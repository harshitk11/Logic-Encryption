module s38417(clk, g51, g563, g1249, g1943, g2637, g3212, g3213, g3214, g3215, g3216, g3217, g3218, g3219, g3220, g3221, g3222, g3223, g3224, g3225, g3226, g3227, g3228, g3229, g3230, g3231, g3232, g3233, g3234, g3993, g4088, g4090, g4200, g4321, g4323, g4450, g4590, g5388, g5437, g5472, g5511, g5549, g5555, g5595, g5612, g5629, g5637, g5648, g5657, g5686, g5695, g5738, g5747, g5796, g6225, g6231, g6313, g6368, g6442, g6447, g6485, g6518, g6573, g6642, g6677, g6712, g6750, g6782, g6837, g6895, g6911, g6944, g6979, g7014, g7052, g7084, g7161, g7194, g7229, g7264, g7302, g7334, g7357, g7390, g7425, g7487, g7519, g7909, g7956, g7961, g8007, g8012, g8021, g8023, g8030, g8082, g8087, g8096, g8106, g8167, g8175, g8249, g8251, g8258, g8259, g8260, g8261, g8262, g8263, g8264, g8265, g8266, g8267, g8268, g8269, g8270, g8271, g8272, g8273, g8274, g8275, g16297, g16355, g16399, g16437, g16496, g24734, g25420, g25435, g25442, g25489, g26104, g26135, g26149, g27380);
input clk, g51, g563, g1249, g1943, g2637, g3212, g3213, g3214, g3215, g3216, g3217, g3218, g3219, g3220, g3221, g3222, g3223, g3224, g3225, g3226, g3227, g3228, g3229, g3230, g3231, g3232, g3233, g3234;
output g3993, g4088, g4090, g4200, g4321, g4323, g4450, g4590, g5388, g5437, g5472, g5511, g5549, g5555, g5595, g5612, g5629, g5637, g5648, g5657, g5686, g5695, g5738, g5747, g5796, g6225, g6231, g6313, g6368, g6442, g6447, g6485, g6518, g6573, g6642, g6677, g6712, g6750, g6782, g6837, g6895, g6911, g6944, g6979, g7014, g7052, g7084, g7161, g7194, g7229, g7264, g7302, g7334, g7357, g7390, g7425, g7487, g7519, g7909, g7956, g7961, g8007, g8012, g8021, g8023, g8030, g8082, g8087, g8096, g8106, g8167, g8175, g8249, g8251, g8258, g8259, g8260, g8261, g8262, g8263, g8264, g8265, g8266, g8267, g8268, g8269, g8270, g8271, g8272, g8273, g8274, g8275, g16297, g16355, g16399, g16437, g16496, g24734, g25420, g25435, g25442, g25489, g26104, g26135, g26149, g27380;
wire clk, g51, g563, g1249, g1943, g2637, g3212, g3213, g3214, g3215, g3216, g3217, g3218, g3219, g3220, g3221, g3222, g3223, g3224, g3225, g3226, g3227, g3228, g3229, g3230, g3231, g3232, g3233, g3234;
wire g2814, g2817, g2933, g2950, g2883, g2888, g2896, g2892, g2903, g2900, g2908;
wire g2912, g2917, g2924, g2920, g2984, g2985, g2930, g2929, g2879, g2934, g2935;
wire g2938, g2941, g2944, g2947, g2953, g2956, g2959, g2962, g2963, g2966, g2969;
wire g2972, g2975, g2978, g2981, g2874, g1506, g1501, g1496, g1491, g1486, g1481;
wire g1476, g1471, g2877, g2861, g813, g2864, g809, g2867, g805, g2870, g801;
wire g2818, g797, g2821, g793, g2824, g789, g2827, g785, g2830, g2873, g2833;
wire g125, g2836, g121, g2839, g117, g2842, g113, g2845, g109, g2848, g105;
wire g2851, g101, g2854, g97, g2858, g2857, g2200, g2195, g2190, g2185, g2180;
wire g2175, g2170, g2165, g2878, g3129, g3117, g3109, g3210, g3211, g3084, g3085;
wire g3086, g3087, g3091, g3092, g3093, g3094, g3095, g3096, g3097, g3098, g3099;
wire g3100, g3101, g3102, g3103, g3104, g3105, g3106, g3107, g3108, g3155, g3158;
wire g3161, g3164, g3167, g3170, g3173, g3176, g3179, g3182, g3185, g3088, g3191;
wire g3194, g3197, g3198, g3201, g3204, g3207, g3188, g3133, g3132, g3128, g3127;
wire g3126, g3125, g3124, g3123, g3120, g3114, g3113, g3112, g3110, g3111, g3139;
wire g3136, g3134, g3135, g3151, g3142, g3147, g185, g138, g135, g165, g130;
wire g131, g129, g133, g134, g132, g142, g143, g141, g145, g146, g144;
wire g148, g149, g147, g151, g152, g150, g154, g155, g153, g157, g158;
wire g156, g160, g161, g159, g163, g164, g162, g169, g170, g168, g172;
wire g173, g171, g175, g176, g174, g178, g179, g177, g186, g189, g192;
wire g231, g234, g237, g195, g198, g201, g240, g243, g246, g204, g207;
wire g210, g249, g252, g255, g213, g216, g219, g258, g261, g264, g222;
wire g225, g228, g267, g270, g273, g92, g88, g83, g79, g74, g70;
wire g65, g61, g56, g52, g180, g182, g181, g276, g405, g401, g309;
wire g354, g343, g346, g369, g358, g361, g384, g373, g376, g398, g388;
wire g391, g408, g411, g414, g417, g420, g423, g427, g428, g426, g429;
wire g432, g435, g438, g441, g444, g448, g449, g447, g312, g313, g314;
wire g315, g316, g317, g318, g319, g320, g322, g323, g321, g403, g404;
wire g402, g450, g451, g452, g453, g454, g279, g280, g281, g282, g283;
wire g284, g285, g286, g287, g288, g289, g290, g291, g299, g305, g308;
wire g297, g296, g295, g294, g304, g303, g302, g301, g300, g298, g342;
wire g349, g350, g351, g352, g353, g357, g364, g365, g366, g367, g368;
wire g372, g379, g380, g381, g382, g383, g387, g394, g395, g396, g397;
wire g324, g325, g331, g337, g545, g551, g550, g554, g557, g510, g513;
wire g523, g524, g564, g569, g570, g571, g572, g573, g574, g565, g566;
wire g567, g568, g489, g474, g481, g485, g486, g487, g488, g455, g458;
wire g461, g477, g478, g479, g480, g484, g464, g465, g468, g471, g528;
wire g535, g542, g543, g544, g548, g549, g499, g558, g559, g576, g577;
wire g575, g579, g580, g578, g582, g583, g581, g585, g586, g584, g587;
wire g590, g593, g596, g599, g602, g614, g617, g620, g605, g608, g611;
wire g490, g493, g496, g506, g507, g508, g509, g514, g515, g516, g517;
wire g518, g519, g520, g525, g529, g530, g531, g532, g533, g534, g536;
wire g537, g538, g541, g623, g626, g629, g630, g659, g640, g633, g653;
wire g646, g660, g672, g666, g679, g686, g692, g699, g700, g698, g702;
wire g703, g701, g705, g706, g704, g708, g709, g707, g711, g712, g710;
wire g714, g715, g713, g717, g718, g716, g720, g721, g719, g723, g724;
wire g722, g726, g727, g725, g729, g730, g728, g732, g733, g731, g735;
wire g736, g734, g738, g739, g737, g826, g823, g853, g818, g819, g817;
wire g821, g822, g820, g830, g831, g829, g833, g834, g832, g836, g837;
wire g835, g839, g840, g838, g842, g843, g841, g845, g846, g844, g848;
wire g849, g847, g851, g852, g850, g857, g858, g856, g860, g861, g859;
wire g863, g864, g862, g866, g867, g865, g873, g876, g879, g918, g921;
wire g924, g882, g885, g888, g927, g930, g933, g891, g894, g897, g936;
wire g939, g942, g900, g903, g906, g945, g948, g951, g909, g912, g915;
wire g954, g957, g960, g780, g776, g771, g767, g762, g758, g753, g749;
wire g744, g740, g868, g870, g869, g963, g1092, g1088, g996, g1041, g1030;
wire g1033, g1056, g1045, g1048, g1071, g1060, g1063, g1085, g1075, g1078, g1095;
wire g1098, g1101, g1104, g1107, g1110, g1114, g1115, g1113, g1116, g1119, g1122;
wire g1125, g1128, g1131, g1135, g1136, g1134, g999, g1000, g1001, g1002, g1003;
wire g1004, g1005, g1006, g1007, g1009, g1010, g1008, g1090, g1091, g1089, g1137;
wire g1138, g1139, g1140, g1141, g966, g967, g968, g969, g970, g971, g972;
wire g973, g974, g975, g976, g977, g978, g986, g992, g995, g984, g983;
wire g982, g981, g991, g990, g989, g988, g987, g985, g1029, g1036, g1037;
wire g1038, g1039, g1040, g1044, g1051, g1052, g1053, g1054, g1055, g1059, g1066;
wire g1067, g1068, g1069, g1070, g1074, g1081, g1082, g1083, g1084, g1011, g1012;
wire g1018, g1024, g1231, g1237, g1236, g1240, g1243, g1196, g1199, g1209, g1210;
wire g1250, g1255, g1256, g1257, g1258, g1259, g1260, g1251, g1252, g1253, g1254;
wire g1176, g1161, g1168, g1172, g1173, g1174, g1175, g1142, g1145, g1148, g1164;
wire g1165, g1166, g1167, g1171, g1151, g1152, g1155, g1158, g1214, g1221, g1228;
wire g1229, g1230, g1234, g1235, g1186, g1244, g1245, g1262, g1263, g1261, g1265;
wire g1266, g1264, g1268, g1269, g1267, g1271, g1272, g1270, g1273, g1276, g1279;
wire g1282, g1285, g1288, g1300, g1303, g1306, g1291, g1294, g1297, g1177, g1180;
wire g1183, g1192, g1193, g1194, g1195, g1200, g1201, g1202, g1203, g1204, g1205;
wire g1206, g1211, g1215, g1216, g1217, g1218, g1219, g1220, g1222, g1223, g1224;
wire g1227, g1309, g1312, g1315, g1316, g1345, g1326, g1319, g1339, g1332, g1346;
wire g1358, g1352, g1365, g1372, g1378, g1385, g1386, g1384, g1388, g1389, g1387;
wire g1391, g1392, g1390, g1394, g1395, g1393, g1397, g1398, g1396, g1400, g1401;
wire g1399, g1403, g1404, g1402, g1406, g1407, g1405, g1409, g1410, g1408, g1412;
wire g1413, g1411, g1415, g1416, g1414, g1418, g1419, g1417, g1421, g1422, g1420;
wire g1424, g1425, g1423, g1520, g1517, g1547, g1512, g1513, g1511, g1515, g1516;
wire g1514, g1524, g1525, g1523, g1527, g1528, g1526, g1530, g1531, g1529, g1533;
wire g1534, g1532, g1536, g1537, g1535, g1539, g1540, g1538, g1542, g1543, g1541;
wire g1545, g1546, g1544, g1551, g1552, g1550, g1554, g1555, g1553, g1557, g1558;
wire g1556, g1560, g1561, g1559, g1567, g1570, g1573, g1612, g1615, g1618, g1576;
wire g1579, g1582, g1621, g1624, g1627, g1585, g1588, g1591, g1630, g1633, g1636;
wire g1594, g1597, g1600, g1639, g1642, g1645, g1603, g1606, g1609, g1648, g1651;
wire g1654, g1466, g1462, g1457, g1453, g1448, g1444, g1439, g1435, g1430, g1426;
wire g1562, g1564, g1563, g1657, g1786, g1782, g1690, g1735, g1724, g1727, g1750;
wire g1739, g1742, g1765, g1754, g1757, g1779, g1769, g1772, g1789, g1792, g1795;
wire g1798, g1801, g1804, g1808, g1809, g1807, g1810, g1813, g1816, g1819, g1822;
wire g1825, g1829, g1830, g1828, g1693, g1694, g1695, g1696, g1697, g1698, g1699;
wire g1700, g1701, g1703, g1704, g1702, g1784, g1785, g1783, g1831, g1832, g1833;
wire g1834, g1835, g1660, g1661, g1662, g1663, g1664, g1665, g1666, g1667, g1668;
wire g1669, g1670, g1671, g1672, g1680, g1686, g1689, g1678, g1677, g1676, g1675;
wire g1685, g1684, g1683, g1682, g1681, g1679, g1723, g1730, g1731, g1732, g1733;
wire g1734, g1738, g1745, g1746, g1747, g1748, g1749, g1753, g1760, g1761, g1762;
wire g1763, g1764, g1768, g1775, g1776, g1777, g1778, g1705, g1706, g1712, g1718;
wire g1925, g1931, g1930, g1934, g1937, g1890, g1893, g1903, g1904, g1944, g1949;
wire g1950, g1951, g1952, g1953, g1954, g1945, g1946, g1947, g1948, g1870, g1855;
wire g1862, g1866, g1867, g1868, g1869, g1836, g1839, g1842, g1858, g1859, g1860;
wire g1861, g1865, g1845, g1846, g1849, g1852, g1908, g1915, g1922, g1923, g1924;
wire g1928, g1929, g1880, g1938, g1939, g1956, g1957, g1955, g1959, g1960, g1958;
wire g1962, g1963, g1961, g1965, g1966, g1964, g1967, g1970, g1973, g1976, g1979;
wire g1982, g1994, g1997, g2000, g1985, g1988, g1991, g1871, g1874, g1877, g1886;
wire g1887, g1888, g1889, g1894, g1895, g1896, g1897, g1898, g1899, g1900, g1905;
wire g1909, g1910, g1911, g1912, g1913, g1914, g1916, g1917, g1918, g1921, g2003;
wire g2006, g2009, g2010, g2039, g2020, g2013, g2033, g2026, g2040, g2052, g2046;
wire g2059, g2066, g2072, g2079, g2080, g2078, g2082, g2083, g2081, g2085, g2086;
wire g2084, g2088, g2089, g2087, g2091, g2092, g2090, g2094, g2095, g2093, g2097;
wire g2098, g2096, g2100, g2101, g2099, g2103, g2104, g2102, g2106, g2107, g2105;
wire g2109, g2110, g2108, g2112, g2113, g2111, g2115, g2116, g2114, g2118, g2119;
wire g2117, g2214, g2211, g2241, g2206, g2207, g2205, g2209, g2210, g2208, g2218;
wire g2219, g2217, g2221, g2222, g2220, g2224, g2225, g2223, g2227, g2228, g2226;
wire g2230, g2231, g2229, g2233, g2234, g2232, g2236, g2237, g2235, g2239, g2240;
wire g2238, g2245, g2246, g2244, g2248, g2249, g2247, g2251, g2252, g2250, g2254;
wire g2255, g2253, g2261, g2264, g2267, g2306, g2309, g2312, g2270, g2273, g2276;
wire g2315, g2318, g2321, g2279, g2282, g2285, g2324, g2327, g2330, g2288, g2291;
wire g2294, g2333, g2336, g2339, g2297, g2300, g2303, g2342, g2345, g2348, g2160;
wire g2156, g2151, g2147, g2142, g2138, g2133, g2129, g2124, g2120, g2256, g2258;
wire g2257, g2351, g2480, g2476, g2384, g2429, g2418, g2421, g2444, g2433, g2436;
wire g2459, g2448, g2451, g2473, g2463, g2466, g2483, g2486, g2489, g2492, g2495;
wire g2498, g2502, g2503, g2501, g2504, g2507, g2510, g2513, g2516, g2519, g2523;
wire g2524, g2522, g2387, g2388, g2389, g2390, g2391, g2392, g2393, g2394, g2395;
wire g2397, g2398, g2396, g2478, g2479, g2477, g2525, g2526, g2527, g2528, g2529;
wire g2354, g2355, g2356, g2357, g2358, g2359, g2360, g2361, g2362, g2363, g2364;
wire g2365, g2366, g2374, g2380, g2383, g2372, g2371, g2370, g2369, g2379, g2378;
wire g2377, g2376, g2375, g2373, g2417, g2424, g2425, g2426, g2427, g2428, g2432;
wire g2439, g2440, g2441, g2442, g2443, g2447, g2454, g2455, g2456, g2457, g2458;
wire g2462, g2469, g2470, g2471, g2472, g2399, g2400, g2406, g2412, g2619, g2625;
wire g2624, g2628, g2631, g2584, g2587, g2597, g2598, g2638, g2643, g2644, g2645;
wire g2646, g2647, g2648, g2639, g2640, g2641, g2642, g2564, g2549, g2556, g2560;
wire g2561, g2562, g2563, g2530, g2533, g2536, g2552, g2553, g2554, g2555, g2559;
wire g2539, g2540, g2543, g2546, g2602, g2609, g2616, g2617, g2618, g2622, g2623;
wire g2574, g2632, g2633, g2650, g2651, g2649, g2653, g2654, g2652, g2656, g2657;
wire g2655, g2659, g2660, g2658, g2661, g2664, g2667, g2670, g2673, g2676, g2688;
wire g2691, g2694, g2679, g2682, g2685, g2565, g2568, g2571, g2580, g2581, g2582;
wire g2583, g2588, g2589, g2590, g2591, g2592, g2593, g2594, g2599, g2603, g2604;
wire g2605, g2606, g2607, g2608, g2610, g2611, g2612, g2615, g2697, g2700, g2703;
wire g2704, g2733, g2714, g2707, g2727, g2720, g2734, g2746, g2740, g2753, g2760;
wire g2766, g2773, g2774, g2772, g2776, g2777, g2775, g2779, g2780, g2778, g2782;
wire g2783, g2781, g2785, g2786, g2784, g2788, g2789, g2787, g2791, g2792, g2790;
wire g2794, g2795, g2793, g2797, g2798, g2796, g2800, g2801, g2799, g2803, g2804;
wire g2802, g2806, g2807, g2805, g2809, g2810, g2808, g2812, g2813, g2811, g3054;
wire g3079, g3080, g3043, g3044, g3045, g3046, g3047, g3048, g3049, g3050, g3051;
wire g3052, g3053, g3055, g3056, g3057, g3058, g3059, g3060, g3061, g3062, g3063;
wire g3064, g3065, g3066, g3067, g3068, g3069, g3070, g3071, g3072, g3073, g3074;
wire g3075, g3076, g3077, g3078, g2997, g2993, g2998, g3006, g3002, g3013, g3010;
wire g3024, g3018, g3028, g3036, g3032, g3040, g2986, g2987, g48, g45, g42;
wire g39, g27, g30, g33, g36, g3083, g26, g2992, g23, g20, g17;
wire g11, g14, g5, g8, g2, g2990, g2991, g1, I13089, g562, I13092;
wire g1248, I13095, g1942, I13098, g2636, I13101, g3235, I13104, g3236, I13107, g3237;
wire I13110, g3238, I13113, g3239, I13116, g3240, I13119, g3241, I13122, g3242, I13125;
wire g3243, I13128, g3244, I13131, g3245, I13134, g3246, I13137, g3247, I13140, g3248;
wire I13143, g3249, I13146, g3250, I13149, g3251, I13152, g3252, I13155, g3253, I13158;
wire g3254, I13161, g3304, g3305, I13165, g3306, g3337, I13169, g3338, g3365, I13173;
wire g3366, I13176, g3398, I13179, g3410, I13182, g3460, g3461, I13186, g3462, g3493;
wire I13190, g3494, g3521, I13194, g3522, I13197, g3554, I13200, g3566, I13203, g3616;
wire g3617, I13207, g3618, g3649, I13211, g3650, g3677, I13215, g3678, I13218, g3710;
wire I13221, g3722, I13224, g3772, g3773, I13228, g3774, g3805, I13232, g3806, g3833;
wire I13236, g3834, I13239, g3866, I13242, g3878, g3897, I13246, g3900, g3919, g3922;
wire g3925, g3928, g3931, g3934, g3937, g3940, g3941, g3942, g3945, g3948, g3951;
wire g3954, g3957, g3960, g3963, g3966, g3969, g3972, g3975, g3978, g3981, g3984;
wire g3987, g3990, I13275, g3993, g3994, g3995, g3996, g3997, g3998, g3999, g4000;
wire g4003, g4006, g4009, g4012, g4015, g4016, g4017, g4020, g4023, g4026, g4029;
wire g4032, g4035, g4038, g4041, g4044, g4047, g4048, g4049, g4052, g4055, g4058;
wire g4061, g4064, g4067, g4070, g4073, g4076, g4079, g4082, g4085, I13316, g4088;
wire g4089, I13320, g4090, g4091, g4092, g4093, g4094, g4095, g4098, g4101, g4104;
wire g4107, g4110, g4111, g4112, g4115, g4118, g4121, g4124, g4127, g4130, g4133;
wire g4136, g4139, g4142, g4143, g4144, g4147, g4150, g4153, g4156, g4159, g4162;
wire g4165, g4168, g4171, g4174, g4175, g4176, g4179, g4182, g4185, g4188, g4191;
wire g4194, g4197, I13366, g4200, g4201, g4202, g4203, g4204, g4205, g4208, g4211;
wire g4214, g4217, g4220, g4221, g4224, g4225, g4228, g4231, g4234, g4237, g4240;
wire g4243, g4246, g4249, g4250, g4251, g4254, g4257, g4260, g4263, g4266, g4269;
wire g4272, g4275, g4278, g4281, g4282, g4283, g4286, g4289, g4292, g4295, g4298;
wire g4301, g4304, g4307, g4310, g4313, g4314, g4315, g4318, I13417, g4321, g4322;
wire I13421, g4323, g4324, g4325, g4326, g4329, g4332, g4335, I13430, g4338, I13433;
wire g4339, g4340, g4343, g4346, g4347, g4348, g4351, g4354, g4357, g4360, g4363;
wire g4366, g4369, g4372, g4375, g4376, g4379, g4380, g4383, g4386, g4389, g4392;
wire g4395, g4398, g4401, g4404, g4405, g4406, g4409, g4412, g4415, g4418, g4421;
wire g4424, g4427, g4430, g4433, g4436, g4437, g4438, g4441, g4444, g4447, I13478;
wire g4450, g4451, g4452, g4453, g4456, g4465, g4468, g4471, g4474, g4475, g4476;
wire g4479, g4480, g4483, g4486, g4489, g4492, g4495, g4498, g4501, g4504, I13501;
wire g4507, I13504, g4508, g4509, g4512, g4515, g4516, g4517, g4520, g4523, g4526;
wire g4529, g4532, g4535, g4538, g4541, g4544, g4545, g4548, g4549, g4552, g4555;
wire g4558, g4561, g4564, g4567, g4570, g4573, g4574, g4575, g4578, g4581, g4584;
wire g4587, I13538, g4590, g4591, g4592, g4595, g4598, g4601, g4602, g4603, g4606;
wire g4609, g4610, g4611, g4614, g4617, g4620, g4623, g4626, g4629, g4632, g4641;
wire g4644, g4647, g4650, g4651, g4652, g4655, g4656, g4659, g4662, g4665, g4668;
wire g4671, g4674, g4677, g4680, I13575, g4683, I13578, g4684, g4685, g4688, g4691;
wire g4692, g4693, g4696, g4699, g4702, g4705, g4708, g4711, g4714, g4717, g4720;
wire g4721, g4724, g4725, g4728, g4731, g4734, I13601, g4735, I13604, g4736, g4737;
wire g4740, g4743, g4746, g4749, g4752, g4753, g4754, g4757, g4760, g4763, g4766;
wire g4769, g4772, g4775, g4778, g4779, g4780, g4783, g4786, g4787, g4788, g4791;
wire g4794, g4797, g4800, g4803, g4806, g4809, g4818, g4821, g4824, g4827, g4828;
wire g4829, g4832, g4833, g4836, g4839, g4842, g4845, g4848, g4851, g4854, g4857;
wire I13652, g4860, I13655, g4861, g4862, g4865, g4868, g4869, g4870, g4873, g4876;
wire g4879, g4882, g4885, g4888, g4891, g4894, g4897, g4898, g4899, g4902, g4905;
wire g4908, I13677, g4911, I13680, g4912, g4913, g4916, g4919, g4922, g4925, g4928;
wire g4929, g4930, g4933, g4936, g4939, g4942, g4945, g4948, g4951, g4954, g4955;
wire g4956, g4959, g4962, g4963, g4964, g4967, g4970, g4973, g4976, g4979, g4982;
wire g4985, g4994, g4997, g5000, g5003, g5004, g5005, g5008, g5009, g5012, g5015;
wire g5018, g5021, g5024, g5027, g5030, g5033, g5034, g5035, g5038, g5041, g5044;
wire g5047, g5050, g5053, g5056, g5057, g5058, g5061, g5064, g5067, I13742, g5070;
wire I13745, g5071, g5072, g5075, g5078, g5081, g5084, g5087, g5088, g5089, g5092;
wire g5095, g5098, g5101, g5104, g5107, g5110, g5113, g5114, g5115, g5118, g5121;
wire g5122, g5123, g5126, g5129, g5132, g5135, g5138, I13775, g5141, g5142, g5145;
wire g5148, g5149, g5150, g5153, g5156, g5159, g5162, g5163, g5164, g5167, g5170;
wire g5173, g5176, g5179, g5182, g5185, g5186, g5187, g5190, g5193, g5196, I13801;
wire g5199, I13804, g5200, g5201, g5204, g5207, g5210, g5213, g5216, g5217, g5218;
wire g5221, g5224, g5227, g5230, g5233, I13820, g5234, g5235, g5238, g5241, g5242;
wire g5243, g5246, g5249, g5252, g5255, g5256, g5257, g5260, g5263, g5266, g5269;
wire g5272, g5275, g5278, g5279, g5280, g5283, g5286, g5289, g5292, g5293, g5296;
wire I13849, g5297, g5298, g5301, g5304, g5305, g5306, g5309, g5312, g5315, g5318;
wire g5319, g5320, g5323, g5326, g5327, g5330, g5333, I13868, g5334, g5335, g5338;
wire g5341, g5342, g5343, g5346, g5349, g5352, g5355, g5358, g5361, g5362, g5363;
wire g5366, g5369, g5372, g5375, g5378, g5379, g5382, g5385, I13892, g5388, g5389;
wire I13896, g5390, g5391, g5394, I13901, g5395, I13904, g5396, I13907, g5397, I13910;
wire g5398, I13913, g5399, I13916, g5400, I13919, g5401, I13922, g5402, I13925, g5403;
wire I13928, g5404, I13931, g5405, I13934, g5406, I13937, g5407, I13940, g5408, I13943;
wire g5409, g5410, I13947, g5411, I13950, g5412, I13953, g5413, I13956, g5414, I13959;
wire g5415, I13962, g5416, I13965, g5417, I13968, g5418, I13971, g5419, I13974, g5420;
wire I13977, g5421, I13980, g5422, g5423, I13984, g5424, I13987, g5425, I13990, g5426;
wire I13993, g5427, g5428, g5431, g5434, I13999, g5437, I14002, g5438, g5469, I14006;
wire g5472, I14009, g5473, g5504, g5507, I14014, g5508, I14017, g5511, I14020, g5512;
wire g5543, g5546, g5547, g5548, I14027, g5549, I14030, g5550, g5551, I14034, g5552;
wire I14037, g5555, I14040, g5556, g5587, g5590, g5591, g5592, g5593, g5594, I14049;
wire g5595, I14052, g5596, g5597, I14056, g5598, g5601, g5604, g5605, g5606, g5609;
wire g5610, g5611, I14066, g5612, I14069, g5613, g5614, I14073, g5615, g5618, g5621;
wire g5622, g5623, g5626, g5627, g5628, I14083, g5629, g5631, g5634, g5635, g5636;
wire I14091, g5637, I14094, g5638, g5639, g5640, g5641, g5642, g5645, g5646, g5647;
wire I14104, g5648, g5651, g5654, g5655, g5656, I14113, g5657, g5659, g5662, g5663;
wire g5664, g5665, g5666, g5667, g5668, g5675, g5679, g5680, g5683, g5684, g5685;
wire I14134, g5686, g5689, g5692, g5693, g5694, I14143, g5695, g5697, g5700, I14149;
wire g5701, g5702, g5703, g5704, g5705, g5706, g5707, g5708, g5712, I14163, g5713;
wire g5714, g5715, g5716, g5717, g5718, g5719, g5720, g5727, g5731, g5732, g5735;
wire g5736, g5737, I14182, g5738, g5741, g5744, g5745, g5746, I14191, g5747, I14195;
wire g5749, g5750, g5751, g5752, g5753, g5754, g5755, g5756, g5759, g5760, g5761;
wire g5762, g5763, g5764, g5765, g5766, g5770, I14219, g5771, g5772, g5773, g5774;
wire g5775, g5776, g5777, g5778, g5785, g5789, g5790, g5793, g5794, g5795, I14238;
wire g5796, I14243, g5799, I14246, g5800, I14249, g5801, g5802, g5803, g5804, g5805;
wire g5806, g5808, g5809, g5810, g5811, g5812, g5813, g5814, g5815, g5818, g5819;
wire g5820, g5821, g5822, g5823, g5824, g5825, g5829, I14280, g5830, g5831, g5832;
wire g5833, g5834, g5835, g5836, g5837, g5844, g5848, I14295, g5849, I14298, g5850;
wire g5851, g5852, g5853, g5854, g5855, I14306, g5856, g5857, g5858, g5859, g5860;
wire g5861, g5862, g5864, g5865, g5866, g5867, g5868, g5869, g5870, g5871, g5874;
wire g5875, g5876, g5877, g5878, g5879, g5880, g5881, g5885, I14338, g5886, g5887;
wire g5888, I14343, g5889, g5890, g5893, g5894, g5895, g5896, g5897, g5898, g5899;
wire g5900, g5901, g5902, I14357, g5903, g5904, g5905, g5906, g5907, g5908, g5909;
wire g5911, g5912, g5913, g5914, g5915, g5916, g5917, g5918, g5921, I14378, g5922;
wire I14381, g5923, I14384, g5924, g5925, g5926, g5927, g5928, g5929, g5932, g5933;
wire g5934, g5935, g5936, g5937, g5938, g5939, g5940, g5941, I14402, g5942, g5943;
wire g5944, g5945, g5946, g5947, g5948, g5950, I14413, g5951, I14416, g5952, g5953;
wire g5954, g5955, g5956, g5957, I14424, g5958, g5959, g5960, g5961, g5962, g5963;
wire g5966, g5967, g5968, g5969, g5970, g5971, g5972, g5973, g5974, g5975, I14442;
wire g5976, g5977, I14446, g5978, I14449, g5979, g5980, g5981, g5982, g5983, g5984;
wire g5985, g5986, I14459, g5987, g5988, g5989, g5990, g5991, g5992, g5995, g5996;
wire g5997, g5998, g5999, I14472, g6000, I14475, g6014, I14478, g6015, g6016, g6017;
wire g6018, g6019, g6020, g6021, g6022, g6023, I14489, g6024, g6025, g6026, g6027;
wire g6028, I14496, g6029, I14499, g6030, I14502, g6031, g6032, g6033, g6034, g6035;
wire g6036, g6037, g6038, g6039, I14513, g6040, I14516, g6041, I14519, g6042, g6043;
wire g6044, g6045, I14525, g6046, g6047, I14529, g6048, I14532, g6051, I14535, g6052;
wire I14538, g6053, I14541, g6054, I14544, g6055, I14547, g6056, I14550, g6057, I14553;
wire g6058, I14556, g6059, I14559, g6060, I14562, g6061, I14565, g6062, I14568, g6063;
wire I14571, g6064, I14574, g6065, I14577, g6066, I14580, g6067, g6068, I14584, g6079;
wire I14587, g6080, I14590, g6081, I14593, g6082, I14596, g6083, I14599, g6084, I14602;
wire g6085, I14605, g6086, g6087, I14609, g6098, I14612, g6099, I14615, g6100, I14618;
wire g6101, I14621, g6102, I14624, g6103, g6104, I14628, g6115, I14631, g6116, I14634;
wire g6117, I14637, g6118, g6119, I14641, g6130, I14644, g6131, I14647, g6134, I14650;
wire g6135, g6136, I14654, g6139, g6140, g6141, g6142, I14660, g6145, g6146, g6149;
wire I14665, g6153, I14668, g6156, g6157, g6161, g6162, g6163, I14675, g6166, g6167;
wire g6170, g6173, g6177, g6180, g6183, g6184, g6188, g6189, g6190, I14688, g6193;
wire g6194, g6197, g6200, g6201, g6204, g6205, g6209, g6212, g6215, g6216, g6220;
wire g6221, g6222, I14704, g6225, g6226, g6227, I14709, g6230, I14712, g6231, I14715;
wire g6232, g6281, g6284, g6288, g6289, g6290, g6293, g6294, g6298, g6301, g6304;
wire g6305, g6309, g6310, I14731, g6313, I14734, g6314, g6363, g6367, I14739, g6368;
wire I14742, g6369, g6418, g6421, g6425, g6426, g6427, g6430, g6431, g6435, g6438;
wire g6441, I14755, g6442, g6443, g6444, I14760, g6447, I14763, g6448, I14766, g6485;
wire I14769, g6486, g6512, g6513, g6517, I14775, g6518, I14778, g6519, g6568, g6572;
wire I14783, g6573, I14786, g6574, g6623, g6626, g6630, g6631, g6632, g6635, g6636;
wire g6637, g6638, g6641, I14799, g6642, I14802, g6643, g6672, g6675, g6676, I14808;
wire g6677, I14811, g6678, g6707, g6711, I14816, g6712, I14819, g6713, I14822, g6750;
wire I14825, g6751, g6776, g6777, g6781, I14831, g6782, I14834, g6783, g6832, g6836;
wire I14839, g6837, I14842, g6838, g6887, g6890, g6894, I14848, g6895, g6896, g6897;
wire g6898, g6901, g6905, g6908, I14857, g6911, I14860, g6912, g6942, g6943, I14865;
wire g6944, I14868, g6945, g6974, g6977, g6978, I14874, g6979, I14877, g6980, g7009;
wire g7013, I14882, g7014, I14885, g7015, I14888, g7052, I14891, g7053, g7078, g7079;
wire g7083, I14897, g7084, I14900, g7085, g7134, g7138, g7139, g7140, g7141, g7142;
wire g7143, g7146, g7149, g7152, g7153, g7156, g7157, g7158, I14917, g7161, I14920;
wire g7162, g7192, g7193, I14925, g7194, I14928, g7195, g7224, g7227, g7228, I14934;
wire g7229, I14937, g7230, g7259, g7263, I14942, g7264, I14945, g7265, I14948, g7302;
wire I14951, g7303, g7328, g7329, g7333, I14957, g7334, g7335, g7336, g7337, g7338;
wire g7342, g7345, g7346, g7347, g7348, g7349, g7352, g7353, g7354, I14973, g7357;
wire I14976, g7358, g7388, g7389, I14981, g7390, I14984, g7391, g7420, g7423, g7424;
wire I14990, g7425, I14993, g7426, g7455, g7459, g7460, g7461, g7462, g7465, g7466;
wire g7471, g7475, g7476, g7477, g7478, g7479, g7482, g7483, g7484, I15012, g7487;
wire I15015, g7488, g7518, I15019, g7519, g7520, g7521, g7522, g7527, g7529, g7530;
wire g7531, g7532, g7533, g7534, g7535, g7538, g7539, g7540, g7541, g7542, g7545;
wire g7548, g7549, g7553, g7554, g7555, g7556, g7557, g7558, g7559, g7560, g7561;
wire g7562, g7566, g7570, g7573, g7574, g7576, g7577, g7578, g7579, g7580, g7581;
wire g7582, g7583, g7587, g7590, g7591, g7592, g7593, g7594, g7595, g7600, g7603;
wire g7604, g7605, g7606, g7607, g7610, g7613, g7614, g7615, g7616, g7619, g7622;
wire g7623, g7626, g7629, g7632, g7635, g7638, g7639, g7642, g7643, g7646, g7649;
wire g7652, g7655, g7658, g7661, g7664, g7667, g7670, g7673, g7676, g7679, g7682;
wire g7685, g7688, g7691, g7694, g7697, g7700, g7703, g7706, g7709, g7712, g7715;
wire g7718, g7721, g7724, g7727, g7730, g7733, g7736, g7739, g7742, g7745, g7748;
wire g7751, g7754, g7757, g7760, g7763, g7766, g7769, g7772, g7776, g7779, g7782;
wire g7785, g7788, g7792, g7796, g7799, g7802, g7806, g7809, g7812, g7815, g7819;
wire g7822, g7823, g7826, g7827, g7830, g7833, g7834, g7837, g7838, g7841, g7842;
wire g7845, g7848, g7849, g7852, g7856, g7857, g7858, g7861, g7862, g7865, g7868;
wire g7869, g7872, g7877, g7878, g7879, g7880, g7888, g7891, g7892, g7897, g7898;
wire g7899, g7900, I15222, g7901, g7906, I15226, g7909, g7910, I15230, g7911, g7912;
wire g7915, g7916, g7919, g7924, g7925, g7926, g7927, g7928, I15256, g7936, g7949;
wire g7950, g7953, I15262, g7956, g7957, g7958, I15267, g7961, g7962, I15271, g7963;
wire g7964, g7967, g7971, g7972, g7973, g7974, g7975, I15288, g7976, g7989, g7990;
wire g7993, g7996, g7999, g8000, g8001, g8004, I15299, g8007, g8008, g8009, I15304;
wire g8012, g8013, I15308, g8014, g8015, g8018, I15313, g8021, g8022, I15317, g8023;
wire g8024, g8025, g8026, g8027, g8028, g8029, I15326, g8030, I15329, g8031, g8044;
wire g8045, g8053, g8056, g8059, g8062, g8065, g8068, g8071, g8074, g8075, g8076;
wire g8079, I15345, g8082, g8083, g8084, I15350, g8087, g8088, I15354, g8089, g8090;
wire g8093, I15359, g8096, g8097, g8098, g8099, g8100, g8101, g8102, g8103, I15369;
wire g8106, I15372, g8107, g8120, g8123, g8126, g8129, g8132, g8135, g8138, g8141;
wire g8144, g8147, g8150, g8153, g8156, g8159, g8160, g8161, g8164, I15392, g8167;
wire g8168, g8169, g8172, I15398, g8175, g8176, g8177, g8178, g8179, g8180, g8181;
wire g8182, g8183, g8191, g8194, g8197, g8200, g8203, g8206, g8209, g8212, g8215;
wire g8218, g8221, g8224, g8227, g8230, g8233, g8236, g8239, g8242, g8245, g8246;
wire I15429, g8249, g8250, I15433, g8251, g8252, g8253, g8254, g8255, g8256, g8257;
wire I15442, g8258, I15445, g8259, I15448, g8260, I15451, g8261, I15454, g8262, I15457;
wire g8263, I15460, g8264, I15463, g8265, I15466, g8266, I15469, g8267, I15472, g8268;
wire I15475, g8269, I15478, g8270, I15481, g8271, I15484, g8272, I15487, g8273, I15490;
wire g8274, I15493, g8275, g8276, g8277, g8278, I15499, g8284, g8285, g8286, g8287;
wire I15505, g8293, g8294, g8295, g8296, I15511, g8302, g8303, g8304, g8305, I15517;
wire g8311, g8312, g8313, g8317, I15523, g8321, I15526, g8324, I15532, g8330, I15535;
wire g8333, I15538, g8336, I15543, g8341, I15546, g8344, I15549, g8347, I15553, g8351;
wire I15556, g8354, I15559, g8357, I15562, g8360, I15565, g8363, I15568, g8366, I15571;
wire g8369, I15574, g8372, I15577, g8375, I15580, g8378, I15584, g8382, I15590, g8388;
wire I15593, g8391, I15599, g8397, I15602, g8400, I15605, g8403, I15610, g8408, I15613;
wire g8411, I15616, g8414, I15620, g8418, I15623, g8421, I15626, g8424, I15629, g8427;
wire I15636, g8434, I15642, g8440, I15645, g8443, I15651, g8449, I15654, g8452, I15657;
wire g8455, I15662, g8460, I15671, g8469, I15677, g8475, I15680, g8478, I15696, g8494;
wire g8514, g8530, g8568, I15771, g8569, I15779, g8575, I15784, g8578, I15787, g8579;
wire g8580, g8587, g8594, I15794, g8602, g8605, I15800, g8614, I15803, g8617, I15806;
wire g8620, I15810, g8622, I15815, g8627, I15818, g8630, I15822, g8632, I15827, g8637;
wire I15830, g8640, I15833, g8643, I15836, g8646, I15839, g8649, I15843, g8651, I15847;
wire g8655, I15850, g8658, I15853, g8659, I15856, g8662, I15859, g8665, I15863, g8667;
wire I15866, g8670, I15869, g8673, I15873, g8677, I15876, g8678, I15879, g8681, I15882;
wire g8684, I15887, g8689, I15890, g8690, I15893, g8693, I15896, g8696, I15899, g8699;
wire I15902, g8700, I15909, g8707, I15912, g8708, I15915, g8711, I15918, g8714, I15922;
wire g8718, I15925, g8719, I15932, g8726, I15935, g8745, I15938, g8748, I15942, g8752;
wire I15946, g8756, I15949, g8757, I15955, g8763, I15958, g8766, I15961, g8769, I15964;
wire g8770, I15967, g8771, I15971, g8775, I15975, g8779, I15978, g8780, I15983, g8785;
wire I15986, g8788, I15989, g8791, I15992, g8792, I15995, g8793, I15998, g8794, I16002;
wire g8798, I16006, g8802, I16009, g8805, I16012, g8808, I16015, g8809, I16018, g8810;
wire I16021, g8811, I16024, g8812, I16027, g8813, I16031, g8817, I16034, g8820, I16037;
wire g8821, g8822, I16041, g8823, I16044, g8824, I16047, g8825, I16050, g8826, I16053;
wire g8827, I16056, g8828, I16059, g8829, I16062, g8832, I16065, g8835, I16068, g8836;
wire I16071, g8839, I16074, g8840, I16079, g8843, I16082, g8844, I16085, g8845, g8846;
wire I16089, g8847, I16092, g8850, I16095, g8851, I16098, g8852, I16101, g8853, I16104;
wire g8856, I16107, g8859, I16110, g8860, I16114, g8862, I16117, g8863, I16120, g8866;
wire I16123, g8867, I16128, g8870, I16131, g8871, I16134, g8872, g8873, I16138, g8874;
wire I16141, g8877, I16144, g8878, I16147, g8879, I16150, g8882, I16153, g8885, I16156;
wire g8888, I16159, g8891, I16163, g8893, I16166, g8894, I16169, g8897, I16172, g8898;
wire I16176, g8900, I16179, g8901, I16182, g8904, I16185, g8905, I16190, g8908, I16193;
wire g8909, I16196, g8910, g8911, I16200, g8912, I16203, g8915, I16206, g8918, I16209;
wire g8921, I16212, g8924, I16215, g8925, I16218, g8928, I16221, g8931, I16225, g8933;
wire I16228, g8934, I16231, g8937, I16234, g8938, I16238, g8940, I16241, g8941, I16244;
wire g8944, I16247, g8945, I16252, g8948, I16255, g8949, I16258, g8952, I16261, g8955;
wire I16264, g8958, I16267, g8961, I16270, g8964, I16273, g8965, I16276, g8968, I16279;
wire g8971, I16283, g8973, I16286, g8974, I16289, g8977, I16292, g8978, I16296, g8980;
wire g8983, I16300, g8984, I16303, g8987, I16306, g8990, I16309, g8993, I16312, g8996;
wire I16315, g8997, I16318, g9000, I16321, g9003, I16325, g9005, I16328, g9006, I16332;
wire g9010, I16335, g9013, I16338, g9016, I16341, g9019, I16344, g9022, I16347, g9025;
wire g9027, I16354, g9035, I16357, g9038, I16360, g9041, I16363, g9044, g9050, I16372;
wire g9058, g9067, g9084, I16432, g9128, I16438, g9134, I16444, g9140, I16450, g9146;
wire I16453, g9149, g9150, I16457, g9159, g9160, g9161, I16462, g9170, I16465, g9173;
wire g9174, I16469, g9183, I16472, g9184, g9187, I16476, g9196, I16479, g9199, I16482;
wire g9202, g9203, I16486, g9212, I16489, g9215, g9216, I16493, g9225, g9226, g9227;
wire g9228, I16499, g9229, g9232, I16504, g9242, I16507, g9245, g9248, I16511, g9257;
wire I16514, g9260, I16517, g9263, g9264, I16521, g9273, I16524, g9276, g9277, g9286;
wire g9287, g9288, g9289, I16532, g9290, g9293, I16538, g9303, I16541, g9306, I16544;
wire g9309, g9310, I16549, g9320, I16552, g9323, g9326, I16556, g9335, I16559, g9338;
wire I16562, g9341, g9342, I16566, g9351, I16569, g9354, g9355, g9356, I16578, g9368;
wire I16581, g9371, g9374, I16587, g9384, I16590, g9387, I16593, g9390, g9391, I16598;
wire g9401, I16601, g9404, g9407, I16605, g9416, I16608, g9419, I16611, g9422, g9423;
wire g9424, g9425, g9426, g9427, I16624, g9443, I16627, g9446, I16630, g9449, I16633;
wire g9450, g9453, I16641, g9465, I16644, g9468, g9471, I16650, g9481, I16653, g9484;
wire I16656, g9487, g9488, I16661, g9498, I16664, g9501, g9504, g9505, g9506, g9507;
wire I16677, g9524, g9527, I16681, g9528, I16684, g9531, g9569, I16694, g9585, I16697;
wire g9588, I16700, g9591, I16703, g9592, g9595, I16711, g9607, I16714, g9610, g9613;
wire I16720, g9623, I16723, g9626, I16726, g9629, I16741, g9640, I16744, g9641, I16747;
wire g9644, g9649, I16759, g9666, g9669, I16763, g9670, I16766, g9673, g9711, I16776;
wire g9727, I16779, g9730, I16782, g9733, I16785, g9734, g9737, I16793, g9749, I16796;
wire g9752, g9755, g9756, g9757, g9758, I16811, g9767, I16814, g9770, I16832, g9786;
wire I16835, g9787, I16838, g9790, g9795, I16850, g9812, g9815, I16854, g9816, I16857;
wire g9819, g9857, I16867, g9873, I16870, g9876, I16873, g9879, I16876, g9880, g9884;
wire g9885, g9886, I16897, g9895, I16900, g9898, I16915, g9913, I16918, g9916, I16936;
wire g9932, I16939, g9933, I16942, g9936, g9941, I16954, g9958, g9961, I16958, g9962;
wire I16961, g9965, I16972, g10004, g10015, I16984, g10016, I16987, g10017, I16990, g10018;
wire I16993, g10021, I17009, g10049, I17012, g10052, I17027, g10067, I17030, g10070, I17048;
wire g10086, I17051, g10087, I17054, g10090, I17066, g10096, g10099, I17070, g10100, I17081;
wire g10109, g10124, I17097, g10125, I17100, g10126, I17103, g10127, I17106, g10130, I17122;
wire g10158, I17125, g10161, I17140, g10176, I17143, g10179, I17159, g10189, I17184, g10214;
wire g10229, I17200, g10230, I17203, g10231, I17206, g10232, I17209, g10235, I17225, g10263;
wire I17228, g10266, I17235, g10273, I17238, g10276, I17278, g10316, g10331, I17294, g10332;
wire I17297, g10333, I17300, g10334, I17303, g10337, I17311, g10357, I17363, g10409, I17370;
wire g10416, I17373, g10419, g10424, g10481, I17433, g10482, g10486, g10500, I17483, g10542;
wire I17486, g10545, g10549, g10560, g10574, I17527, g10601, g10606, g10617, g10631, I17557;
wire g10646, g10653, g10664, g10683, g10694, g10714, g10730, g10735, g10749, g10754, g10765;
wire g10766, g10767, g10772, g10773, I17627, g10779, g10783, I17632, g10787, g10788, I17637;
wire g10792, I17641, g10796, I17645, g10800, I17649, g10804, I17653, g10808, g10809, I17658;
wire g10813, I17662, g10817, I17666, g10821, I17670, g10825, I17673, g10826, g10829, I17677;
wire g10830, I17681, g10834, I17685, g10838, I17689, g10842, I17692, g10843, g10846, g10847;
wire g10848, I17698, g10849, I17701, g10850, I17705, g10854, I17709, g10858, I17712, g10859;
wire I17715, g10862, g10865, g10866, g10867, I17721, g10868, I17724, g10869, I17727, g10870;
wire I17730, g10871, I17734, g10875, I17737, g10876, I17740, g10877, I17743, g10880, I17746;
wire g10883, g10886, I17750, g10887, I17753, g10888, I17756, g10889, I17759, g10890, I17762;
wire g10891, I17765, g10892, I17768, g10895, I17771, g10898, I17774, g10901, g10904, g10905;
wire g10906, I17780, g10907, I17783, g10908, I17786, g10909, I17789, g10910, I17792, g10911;
wire I17795, g10912, I17798, g10915, I17801, g10918, I17804, g10921, I17807, g10924, g10927;
wire g10928, g10929, I17813, g10930, I17816, g10931, I17819, g10932, I17822, g10933, I17825;
wire g10934, I17828, g10935, I17831, g10936, I17834, g10937, I17837, g10940, I17840, g10943;
wire I17843, g10946, I17846, g10949, I17849, g10952, g10961, g10962, I17854, g10963, I17857;
wire g10966, I17860, g10967, I17863, g10968, I17866, g10969, I17869, g10972, I17872, g10973;
wire I17875, g10974, I17878, g10977, I17881, g10980, I17884, g10983, g10986, g10987, I17889;
wire g10988, I17892, g10991, I17895, g10994, I17898, g10995, I17901, g10996, I17904, g10999;
wire I17907, g11002, I17910, g11003, I17913, g11004, I17916, g11007, I17919, g11008, I17922;
wire g11011, I17925, g11014, I17928, g11017, g11020, g11021, I17933, g11022, I17936, g11025;
wire I17939, g11028, I17942, g11031, I17945, g11032, I17948, g11035, I17951, g11036, I17954;
wire g11039, I17957, g11042, I17960, g11045, I17963, g11048, I17966, g11051, I17969, g11054;
wire I17972, g11055, I17975, g11056, I17978, g11059, I17981, g11063, I17984, g11066, g11069;
wire g11078, I17989, g11079, I17992, g11082, I17995, g11085, I17998, g11088, I18001, g11091;
wire I18004, g11092, I18007, g11095, I18010, g11098, I18013, g11101, I18016, g11102, I18019;
wire g11105, I18022, g11108, I18025, g11111, I18028, g11114, I18031, g11117, I18034, g11120;
wire I18037, g11123, I18040, g11126, I18043, g11129, I18046, g11132, I18049, g11135, I18052;
wire g11138, I18055, g11141, I18058, g11144, I18061, g11145, I18064, g11148, I18067, g11151;
wire I18070, g11154, I18073, g11157, I18076, g11160, I18079, g11163, I18082, g11166, I18085;
wire g11169, I18088, g11170, I18091, g11173, I18094, g11176, I18097, g11179, I18100, g11182;
wire I18103, g11185, g11190, I18121, g11199, I18124, g11202, I18127, g11205, I18130, g11208;
wire I18133, g11209, I18136, g11210, I18139, g11213, I18142, g11216, I18145, g11219, I18148;
wire g11222, I18151, g11225, I18154, g11228, I18157, g11231, I18160, g11234, I18163, g11237;
wire I18166, g11240, I18169, g11243, I18172, g11246, I18175, g11249, I18178, g11252, I18181;
wire g11255, I18184, g11256, I18187, g11259, I18211, g11265, I18214, g11268, I18217, g11271;
wire I18220, g11274, I18223, g11277, I18226, g11278, I18229, g11281, I18232, g11284, I18235;
wire g11287, I18238, g11290, I18241, g11291, I18244, g11294, I18247, g11297, I18250, g11300;
wire I18253, g11303, I18256, g11306, I18259, g11309, I18262, g11312, I18265, g11315, I18268;
wire g11318, I18271, g11321, I18274, g11324, I18277, g11327, g11332, I18295, g11341, I18298;
wire g11344, I18302, g11348, I18305, g11351, I18308, g11354, I18311, g11355, I18314, g11358;
wire I18317, g11361, I18320, g11364, I18323, g11367, I18326, g11370, I18329, g11373, I18332;
wire g11376, I18335, g11379, I18338, g11382, I18341, g11385, I18344, g11386, I18347, g11389;
wire I18350, g11392, I18353, g11395, I18356, g11398, I18359, g11401, I18362, g11404, I18365;
wire g11407, I18375, g11411, I18378, g11414, I18381, g11417, I18386, g11422, I18389, g11425;
wire I18392, g11428, I18396, g11432, I18399, g11435, I18402, g11438, I18405, g11441, I18408;
wire g11444, I18411, g11447, I18414, g11450, I18417, g11453, I18420, g11456, I18423, g11459;
wire I18426, g11462, I18429, g11465, I18432, g11468, I18435, g11471, I18438, g11472, I18441;
wire g11475, I18444, g11478, g11481, g11490, I18449, g11491, I18452, g11492, I18455, g11493;
wire I18458, g11494, I18461, g11495, I18464, g11496, I18467, g11497, I18470, g11498, I18473;
wire g11499, I18476, g11500, I18479, g11501, I18482, g11502, I18485, g11503, I18488, g11504;
wire I18491, g11505, I18494, g11506, I18497, g11507, I18500, g11508, I18503, g11509, I18506;
wire g11510, I18509, g11511, I18512, g11512, I18515, g11513, I18518, g11514, I18521, g11515;
wire I18524, g11516, I18527, g11517, I18530, g11518, I18533, g11519, I18536, g11520, I18539;
wire g11521, I18542, g11522, I18545, g11523, I18548, g11524, I18551, g11525, I18554, g11526;
wire I18557, g11527, I18560, g11528, I18563, g11529, I18566, g11530, I18569, g11531, I18572;
wire g11532, I18575, g11533, I18578, g11534, I18581, g11535, I18584, g11536, I18587, g11537;
wire I18590, g11538, I18593, g11539, I18596, g11540, I18599, g11541, I18602, g11542, I18605;
wire g11543, I18608, g11544, I18611, g11545, I18614, g11546, I18617, g11547, I18620, g11548;
wire I18623, g11549, I18626, g11550, I18629, g11551, I18632, g11552, I18635, g11553, I18638;
wire g11554, I18641, g11555, I18644, g11556, I18647, g11557, I18650, g11558, I18653, g11559;
wire I18656, g11560, I18659, g11561, I18662, g11562, I18665, g11563, I18668, g11564, I18671;
wire g11565, I18674, g11566, I18677, g11567, I18680, g11568, I18683, g11569, I18686, g11570;
wire I18689, g11571, I18692, g11572, I18695, g11573, I18698, g11574, I18701, g11575, I18704;
wire g11576, I18707, g11577, I18710, g11578, I18713, g11579, I18716, g11580, I18719, g11581;
wire I18722, g11582, I18725, g11583, I18728, g11584, I18731, g11585, I18734, g11586, I18737;
wire g11587, I18740, g11588, I18743, g11589, I18746, g11590, I18749, g11591, I18752, g11592;
wire I18755, g11593, I18758, g11594, I18761, g11595, I18764, g11596, I18767, g11597, I18770;
wire g11598, I18773, g11599, I18777, g11603, I18780, g11606, I18784, g11608, I18787, g11611;
wire I18791, g11613, I18794, g11616, g11620, g11623, I18810, g11628, I18813, g11629, I18817;
wire g11633, I18820, g11636, I18824, g11638, I18827, g11641, g11642, I18835, g11651, I18838;
wire g11652, I18842, g11656, I18845, g11659, I18854, g11670, I18857, g11671, I18866, g11682;
wire g11706, g11732, g11734, g11735, g11736, g11737, g11740, g11741, g11742, g11743, g11745;
wire g11746, g11747, g11748, I18929, g11749, g11758, g11761, g11762, g11763, g11764, g11765;
wire g11766, I18943, g11769, g11770, g11774, g11775, g11776, g11777, g11778, g11779, g11782;
wire g11783, I18962, g11786, g11787, I18969, g11791, g11794, g11795, g11796, g11797, g11798;
wire g11801, g11802, g11803, g11804, g11808, g11809, I18990, g11812, g11813, g11817, g11818;
wire g11819, g11820, g11821, g11824, g11825, g11826, g11827, g11829, g11834, g11835, g11836;
wire g11837, g11841, g11842, I19025, g11845, g11846, I19030, g11848, g11852, g11853, g11854;
wire g11856, g11857, g11858, g11859, g11862, g11866, g11867, g11868, g11869, g11871, g11876;
wire g11877, g11878, g11879, g11883, g11884, g11886, g11887, g11888, g11891, g11892, g11893;
wire g11894, g11895, g11898, g11899, g11900, g11901, g11904, g11908, g11909, g11910, g11911;
wire g11913, g11918, g11919, g11920, g11921, I19105, g11923, g11927, g11929, g11930, g11931;
wire g11932, g11933, g11936, I19119, g11937, g11941, g11942, g11943, g11944, g11945, g11948;
wire g11949, g11950, g11951, g11954, g11958, g11959, g11960, g11961, g11963, g11968, g11969;
wire g11970, g11971, g11972, g11973, I19160, g11976, g11982, g11983, g11984, g11985, g11986;
wire g11989, I19174, g11990, g11994, g11995, g11996, g11997, g11998, g12001, g12002, g12003;
wire g12004, g12007, I19195, g12009, g12013, g12017, g12020, g12021, g12022, g12023, g12024;
wire g12025, I19208, g12027, I19211, g12030, g12037, g12038, g12039, g12040, g12041, g12042;
wire I19226, g12045, g12051, g12052, g12053, g12054, g12055, g12058, I19240, g12059, g12063;
wire g12064, g12065, g12066, g12067, g12071, g12075, g12076, g12077, g12078, g12084, g12085;
wire g12086, g12087, g12088, g12089, I19271, g12091, I19274, g12094, g12101, g12102, g12103;
wire g12104, g12105, g12106, I19289, g12109, g12115, g12116, g12117, g12118, g12119, g12122;
wire I19303, g12123, I19307, g12125, g12130, g12134, g12135, I19315, g12136, I19318, g12139;
wire I19321, g12142, g12147, g12148, g12149, g12150, g12156, g12157, g12158, g12159, g12160;
wire g12161, I19342, g12163, I19345, g12166, g12173, g12174, g12175, g12176, g12177, g12178;
wire I19360, g12181, g12187, g12191, g12196, g12197, I19374, g12198, I19377, g12201, I19380;
wire g12204, g12209, g12210, g12211, g12212, g12218, g12219, g12220, g12221, g12222, g12223;
wire I19401, g12225, I19404, g12228, g12235, I19412, g12239, I19415, g12242, g12246, g12251;
wire g12252, I19426, g12253, I19429, g12256, I19432, g12259, g12264, g12265, g12266, g12267;
wire g12275, I19449, g12279, I19452, g12282, I19455, g12285, g12289, g12294, g12295, I19466;
wire g12296, I19469, g12299, I19472, g12302, g12308, I19479, g12312, I19482, g12315, I19485;
wire g12318, I19488, g12321, g12325, g12332, I19500, g12333, I19503, g12336, I19507, g12340;
wire I19510, g12343, I19513, g12346, I19516, g12349, g12354, g12362, I19523, g12363, I19526;
wire g12366, I19530, g12370, I19533, g12373, g12378, I19539, g12379, I19542, g12382, I19545;
wire g12385, I19549, g12389, I19552, g12392, g12408, I19557, g12409, I19560, g12412, I19563;
wire g12415, g12420, I19569, g12421, g12424, I19573, g12425, I19576, g12426, g12430, I19582;
wire g12432, g12434, I19587, g12435, I19591, g12437, g12438, I19595, g12439, I19598, g12440;
wire I19602, g12442, I19605, g12443, I19608, g12444, I19611, g12445, I19615, g12447, I19618;
wire g12448, I19621, g12449, I19624, g12450, I19628, g12452, I19631, g12453, I19634, g12454;
wire I19637, g12455, g12456, I19642, g12460, I19645, g12461, I19648, g12462, g12463, g12466;
wire I19654, g12470, I19657, g12471, g12472, g12473, g12476, g12478, g12481, I19667, g12485;
wire g12490, g12493, g12495, g12498, g12502, g12504, g12505, g12510, g12513, g12515, g12518;
wire I19689, g12519, g12521, g12522, g12527, g12530, g12532, g12533, I19702, g12534, g12536;
wire g12537, g12542, I19711, g12543, g12545, g12546, g12547, I19718, g12548, g12551, I19722;
wire g12552, g12553, g12554, I19727, g12555, g12558, g12559, g12560, I19733, g12561, I19736;
wire g12564, I19739, g12565, g12596, g12597, g12598, g12599, g12600, I19747, g12601, I19750;
wire g12604, I19753, g12607, I19756, g12608, I19759, g12611, g12642, g12643, g12644, g12645;
wire g12646, I19767, g12647, I19771, g12651, I19774, g12654, I19777, g12657, g12688, g12689;
wire g12690, g12691, I19784, g12692, I19787, g12695, I19791, g12699, I19794, g12702, I19797;
wire g12705, I19800, g12708, I19803, g12711, g12742, g12743, I19808, g12744, g12748, I19813;
wire g12749, I19816, g12752, I19820, g12756, I19823, g12759, I19826, g12762, I19829, g12765;
wire g12768, I19833, g12769, I19836, g12772, g12775, g12776, g12782, I19844, g12783, I19847;
wire g12786, g12790, I19852, g12791, I19855, g12794, I19859, g12798, I19862, g12801, I19865;
wire g12804, g12807, I19869, g12808, I19872, g12811, g12815, I19877, g12816, g12821, I19883;
wire g12822, I19886, g12825, g12829, I19891, g12830, I19894, g12833, I19898, g12837, I19901;
wire g12840, g12843, I19905, g12844, g12847, g12848, g12850, g12851, g12853, I19915, g12854;
wire g12859, I19921, g12860, I19924, g12863, g12867, I19929, g12868, I19932, g12871, g12874;
wire g12875, g12881, g12882, g12891, g12892, g12894, I19952, g12895, g12900, I19958, g12901;
wire I19961, g12904, g12907, g12909, g12914, g12915, g12921, g12922, g12931, g12932, g12934;
wire I19986, g12935, g12940, g12943, g12944, g12950, g12951, g12960, g12961, I20009, g12962;
wire g12965, g12969, g12972, g12973, g12979, g12980, g12993, g12996, g12997, g12998, g13003;
wire I20062, g13011, g13025, g13033, g13036, g13043, g13046, g13049, g13057, g13060, g13063;
wire g13066, I20117, g13070, g13073, g13076, g13079, g13092, g13095, g13101, g13107, g13117;
wire g13130, g13141, g13148, g13151, g13152, g13153, g13154, g13157, g13158, g13159, g13161;
wire g13162, g13163, g13166, g13167, g13168, g13169, g13170, g13172, g13173, g13174, g13176;
wire g13177, g13178, g13179, g13180, g13181, g13183, g13184, g13185, g13186, g13187, g13188;
wire g13189, g13190, g13191, g13192, g13193, g13195, g13196, g13197, g13198, g13199, g13200;
wire g13201, g13202, g13203, g13204, g13205, g13206, g13207, g13208, g13209, g13210, g13211;
wire g13212, g13213, g13214, I20264, g13215, g13218, g13219, g13220, g13221, g13222, g13223;
wire g13224, g13225, g13226, g13227, I20278, g13229, g13232, g13233, I20283, g13234, g13237;
wire g13238, g13239, g13240, g13241, g13242, g13243, g13244, I20295, g13246, I20299, g13248;
wire g13249, g13250, I20305, g13252, g13255, g13256, I20310, g13257, g13260, g13261, g13262;
wire g13263, g13264, g13265, I20320, g13267, g13268, I20324, g13269, I20328, g13271, g13272;
wire g13273, I20334, g13275, g13278, g13279, I20339, g13280, g13283, g13284, g13285, I20347;
wire g13290, I20351, g13292, g13293, I20355, g13294, I20359, g13296, g13297, g13298, I20365;
wire g13300, g13303, g13304, g13308, g13309, I20376, g13317, I20379, g13318, I20382, g13319;
wire I20386, g13321, I20390, g13323, g13324, I20394, g13325, I20398, g13327, g13328, g13329;
wire g13330, I20407, g13336, I20410, g13339, I20414, g13341, I20417, g13342, I20421, g13344;
wire I20425, g13346, g13347, g13351, g13352, I20441, g13356, I20444, g13359, I20448, g13361;
wire I20451, g13364, I20455, g13366, I20458, g13367, I20462, g13369, g13373, I20476, g13381;
wire I20479, g13384, I20483, g13386, I20486, g13389, I20490, g13391, I20493, g13394, I20497;
wire g13396, I20500, g13397, g13398, g13400, I20514, g13405, I20517, g13406, I20520, g13407;
wire I20523, g13408, I20526, g13409, I20529, g13410, I20532, g13411, I20535, g13412, I20538;
wire g13413, I20541, g13414, I20544, g13415, I20547, g13416, I20550, g13417, I20553, g13418;
wire I20556, g13419, I20559, g13420, I20562, g13421, I20565, g13422, I20568, g13423, I20571;
wire g13424, I20574, g13425, I20577, g13426, I20580, g13427, I20583, g13428, I20586, g13429;
wire I20589, g13430, I20592, g13431, I20595, g13432, I20598, g13433, I20601, g13434, I20604;
wire g13435, I20607, g13436, I20610, g13437, I20613, g13438, I20616, g13439, I20619, g13440;
wire I20622, g13441, I20625, g13442, I20628, g13443, I20631, g13444, I20634, g13445, I20637;
wire g13446, I20640, g13447, I20643, g13448, I20646, g13449, I20649, g13450, I20652, g13451;
wire I20655, g13452, I20658, g13453, I20661, g13454, I20664, g13455, I20667, g13456, I20670;
wire g13457, I20673, g13458, I20676, g13459, I20679, g13460, I20682, g13461, I20685, g13462;
wire I20688, g13463, I20691, g13464, I20694, g13465, I20697, g13466, I20700, g13467, I20703;
wire g13468, I20706, g13469, I20709, g13475, g13519, g13530, g13541, g13552, g13565, g13568;
wire I20791, g13571, I20794, g13572, g13573, g13576, I20799, g13579, I20802, g13580, I20805;
wire g13581, g13582, g13585, I20810, g13588, I20813, g13589, I20816, g13598, I20820, g13600;
wire I20823, g13601, g13602, g13605, I20828, g13608, I20832, g13610, I20836, g13612, I20839;
wire g13613, g13614, I20844, g13620, I20848, g13622, I20852, g13624, g13626, I20858, g13632;
wire I20863, g13635, g13637, g13644, I20873, g13647, g13649, g13657, g13669, g13670, I20886;
wire g13673, g13677, g13687, g13699, g13700, g13706, g13714, g13724, g13736, g13737, I20909;
wire g13741, g13750, g13756, g13764, g13774, g13786, g13791, g13797, g13805, g13817, g13819;
wire g13825, g13836, g13838, g13840, g13848, g13849, g13850, g13852, g13856, g13857, g13858;
wire g13859, g13861, I20959, g13863, g13864, g13866, g13867, g13868, g13869, g13872, g13873;
wire g13879, g13881, g13882, g13883, g13885, g13886, g13894, g13895, g13901, g13903, g13906;
wire g13907, g13918, g13922, g13926, g13927, g13935, g13936, g13942, g13945, g13946, I21012;
wire g13954, g13958, g13962, g13963, g13974, g13978, g13982, g13983, g13991, g13992, g13999;
wire g14000, g14001, I21037, g14008, g14011, g14015, g14016, I21045, g14024, g14028, g14032;
wire g14033, g14044, g14048, g14052, g14053, g14061, g14062, I21064, g14068, g14071, g14079;
wire g14086, g14090, g14091, g14092, I21075, g14099, g14102, g14106, g14107, I21083, g14115;
wire g14119, g14123, g14124, g14135, g14139, I21096, g14144, g14148, g14153, g14158, g14165;
wire g14171, g14175, g14176, g14177, I21108, g14183, g14186, g14194, g14201, g14205, g14206;
wire g14207, I21119, g14214, g14217, g14221, g14222, I21127, g14230, g14234, g14238, g14244;
wire g14249, g14252, g14256, I21137, g14259, g14263, g14268, g14273, g14280, g14286, g14290;
wire g14291, g14292, I21149, g14298, g14301, g14309, g14316, g14320, g14321, g14322, I21160;
wire g14329, g14332, I21165, g14337, g14342, g14347, g14352, g14355, g14359, g14360, g14366;
wire g14371, g14374, g14378, I21178, g14381, g14385, g14390, g14395, g14402, g14408, g14412;
wire g14413, g14414, I21190, g14420, g14423, g14431, g14438, g14442, g14450, g14454, g14459;
wire g14464, g14467, g14471, g14472, g14478, g14483, g14486, g14490, I21208, g14493, g14497;
wire g14502, g14507, g14514, g14520, g14524, g14525, g14529, g14537, g14541, g14546, g14551;
wire g14554, g14558, g14559, g14565, g14570, g14573, g14577, g14580, g14584, g14592, g14596;
wire g14601, g14606, g14609, g14613, g14614, g14618, g14626, I21241, g14630, g14637, g14641;
wire I21246, g14642, I21249, g14650, I21252, g14657, g14668, I21256, g14669, I21259, g14677;
wire I21262, g14684, g14685, I21267, g14691, g14702, I21271, g14703, I21274, g14711, I21277;
wire g14718, g14719, I21282, g14725, g14736, I21286, g14737, I21289, g14745, I21292, g14746;
wire g14747, I21297, g14753, g14764, I21301, g14765, I21304, g14766, g14768, I21310, g14774;
wire I21313, g14775, g14776, g14794, I21318, g14795, I21321, g14796, g14797, g14811, I21326;
wire g14829, I21329, g14830, g14831, g14837, g14849, g14863, g14881, I21337, g14882, I21340;
wire g14883, g14885, g14895, g14904, g14910, g14922, g14936, I21351, g14954, I21354, g14955;
wire g14959, I21361, g14960, I21364, g14963, g14966, g14976, g14985, g14991, g15003, g15017;
wire I21374, g15018, I21377, g15019, I21381, g15021, g15022, g15032, g15033, I21389, g15034;
wire I21392, g15037, I21395, g15040, I21398, g15043, g15048, I21404, g15049, I21407, g15052;
wire g15055, g15065, g15074, g15080, I21415, g15092, I21420, g15095, g15096, I21426, g15106;
wire I21429, g15109, I21432, g15112, I21435, g15115, g15118, g15128, g15129, I21443, g15130;
wire I21446, g15133, I21449, g15136, I21452, g15139, g15144, I21458, g15145, I21461, g15148;
wire g15151, g15161, g15170, g15174, g15175, g15176, g15177, I21476, g15179, I21479, g15182;
wire I21482, g15185, g15188, I21488, g15198, I21491, g15201, I21494, g15204, I21497, g15207;
wire g15210, g15220, g15221, I21505, g15222, I21508, g15225, I21511, g15228, I21514, g15231;
wire g15236, I21520, g15237, I21523, g15240, I21531, g15248, I21534, g15251, I21537, g15254;
wire g15260, g15261, g15262, g15263, I21548, g15265, I21551, g15268, I21554, g15271, g15274;
wire I21560, g15284, I21563, g15287, I21566, g15290, I21569, g15293, g15296, g15306, g15307;
wire I21577, g15308, I21580, g15311, I21583, g15314, I21586, g15317, g15322, g15323, I21595;
wire g15326, I21598, g15329, I21601, g15332, I21609, g15340, I21612, g15343, I21615, g15346;
wire g15352, g15353, g15354, g15355, I21626, g15357, I21629, g15360, I21632, g15363, g15366;
wire I21638, g15376, I21641, g15379, I21644, g15382, I21647, g15385, g15390, I21655, g15393;
wire I21658, g15396, I21661, g15399, I21666, g15404, g15408, g15409, I21674, g15412, I21677;
wire g15415, I21680, g15418, I21688, g15426, I21691, g15429, I21694, g15432, g15438, g15439;
wire g15440, g15441, I21705, g15443, I21708, g15446, I21711, g15449, g15458, I21720, g15461;
wire I21723, g15464, I21726, g15467, I21730, g15471, g15474, I21736, g15477, I21739, g15480;
wire I21742, g15483, I21747, g15488, g15492, g15493, I21755, g15496, I21758, g15499, I21761;
wire g15502, I21769, g15510, I21772, g15513, I21775, g15516, I21780, g15521, g15524, g15525;
wire I21787, g15528, I21790, g15531, I21793, g15534, I21796, g15537, g15544, I21803, g15547;
wire I21806, g15550, I21809, g15553, I21813, g15557, g15560, I21819, g15563, I21822, g15566;
wire I21825, g15569, I21830, g15574, g15578, g15579, I21838, g15582, I21841, g15585, I21844;
wire g15588, I21852, g15596, I21855, g15599, g15602, g15603, I21862, g15606, I21865, g15609;
wire I21868, g15612, I21871, g15615, g15622, I21878, g15625, I21881, g15628, I21884, g15631;
wire I21888, g15635, g15638, I21894, g15641, I21897, g15644, I21900, g15647, I21905, g15652;
wire I21908, g15655, g15659, g15665, I21918, g15667, I21923, g15672, I21926, g15675, g15678;
wire g15679, I21933, g15682, I21936, g15685, I21939, g15688, I21942, g15691, g15698, I21949;
wire g15701, I21952, g15704, I21955, g15707, I21959, g15711, I21962, g15714, g15722, g15724;
wire I21974, g15726, I21979, g15731, I21982, g15734, g15737, g15738, I21989, g15741, I21992;
wire g15744, I21995, g15747, I21998, g15750, g15762, g15764, I22014, g15766, I22019, g15771;
wire I22022, g15774, I22025, g15777, g15790, g15792, I22044, g15794, g15800, g15813, g15859;
wire I22120, g15876, g15880, g15890, g15904, g15913, g15923, g15933, g15942, g15952, g15962;
wire g15971, g15981, I22163, g15989, g15991, g15994, g15997, g16001, g16002, g16005, g16007;
wire g16011, g16012, g16013, g16014, g16023, g16024, g16025, g16026, g16027, g16034, g16035;
wire g16039, g16040, g16041, g16042, g16043, g16044, g16054, g16055, g16056, g16057, g16061;
wire g16062, g16063, g16064, g16065, g16075, g16088, g16090, g16091, g16092, g16093, g16097;
wire g16098, g16099, g16113, g16126, g16128, g16129, g16130, g16131, g16142, g16154, g16164;
wire g16177, g16179, g16180, g16189, g16201, g16213, g16223, g16236, g16243, g16254, g16266;
wire g16278, g16287, g16293, I22382, g16297, g16302, g16313, g16325, g16337, g16351, I22414;
wire g16355, g16360, g16371, g16395, I22444, g16399, g16404, g16433, I22475, g16437, g16466;
wire I22503, g16467, I22506, g16468, I22509, g16469, I22512, g16470, I22515, g16471, I22518;
wire g16472, I22521, g16473, I22524, g16474, I22527, g16475, I22530, g16476, I22533, g16477;
wire I22536, g16478, I22539, g16479, I22542, g16480, I22545, g16481, I22548, g16482, I22551;
wire g16483, I22554, g16484, I22557, g16485, I22560, g16486, I22563, g16487, I22566, g16488;
wire I22569, g16489, I22572, g16490, I22575, g16491, I22578, g16492, I22581, g16493, I22584;
wire g16494, I22587, g16495, I22590, g16496, I22593, g16497, g16501, I22599, g16506, g16507;
wire I22604, g16514, g16515, g16523, I22611, g16528, g16529, I22618, g16540, g16543, g16546;
wire g16554, I22626, g16559, g16560, I22640, g16572, g16575, g16578, g16586, I22651, g16596;
wire g16599, g16602, I22657, g16608, I22663, g16616, g16619, I22667, g16622, I22671, g16626;
wire I22676, g16633, I22679, g16636, I22683, g16640, I22687, g16644, I22690, g16647, I22694;
wire g16651, I22699, g16656, I22702, g16659, g16665, I22715, g16673, I22718, g16676, g16682;
wire g16686, I22726, g16694, g16697, I22730, g16702, g16708, g16712, I22737, g16719, g16722;
wire I22741, g16725, g16728, I22745, g16733, g16739, g16743, g16749, I22752, g16758, I22755;
wire g16761, g16764, I22759, g16767, g16770, I22763, g16775, g16781, I22768, g16785, I22771;
wire g16788, g16791, I22775, g16794, g16797, g16804, g16809, I22783, g16813, I22786, g16814;
wire I22789, g16817, g16820, g16825, I22797, g16830, I22800, g16831, I22803, g16832, g16836;
wire g16840, I22810, g16842, I22813, g16843, g16846, I22820, g16848, I22823, g16849, I22828;
wire g16852, I22836, g16858, I22842, g16862, I22845, g16863, g16867, I22852, g16877, I22855;
wire g16878, I22860, g16881, g16884, g16895, I22866, g16905, I22869, g16906, I22875, g16910;
wire g16913, g16924, I22881, g16934, I22893, g16940, g16943, g16954, I22912, g16971, g16974;
wire g17029, g17057, g17063, g17092, g17098, g17130, g17136, g17157, I23253, g17189, I23274;
wire g17200, g17203, I23287, g17207, g17208, I23292, g17212, g17214, g17217, I23309, g17227;
wire I23314, g17230, I23317, g17233, I23323, g17237, I23326, g17240, I23329, g17243, I23335;
wire g17249, I23338, g17252, I23341, g17255, g17258, I23345, g17259, I23348, g17262, I23351;
wire g17265, I23358, g17272, I23361, g17275, I23364, g17278, g17281, I23368, g17282, I23371;
wire g17285, I23374, g17288, I23377, g17291, I23380, g17294, I23383, g17297, I23386, g17300;
wire I23392, g17304, I23395, g17307, I23398, g17310, g17313, g17314, I23403, g17315, I23406;
wire g17318, I23409, g17321, I23412, g17324, I23415, g17327, I23418, g17330, I23421, g17333;
wire I23424, g17336, I23430, g17342, I23433, g17345, I23436, g17348, g17351, I23442, g17354;
wire I23445, g17357, I23448, g17360, I23451, g17363, I23454, g17366, I23457, g17369, I23460;
wire g17372, I23463, g17375, I23466, g17378, I23472, g17384, I23475, g17387, I23478, g17390;
wire g17394, I23487, g17399, I23490, g17402, I23493, g17405, I23498, g17410, I23501, g17413;
wire I23504, g17416, I23507, g17419, I23510, g17422, I23513, g17425, I23518, g17430, I23521;
wire g17433, I23524, g17436, I23527, g17439, I23530, g17442, g17445, I23539, g17451, I23542;
wire g17454, I23545, g17457, I23553, g17465, I23556, g17468, I23559, g17471, I23564, g17476;
wire I23567, g17479, I23570, g17482, I23575, g17487, I23578, g17490, I23581, g17493, I23584;
wire g17496, g17499, I23588, g17500, I23591, g17503, I23599, g17511, I23602, g17514, I23605;
wire g17517, I23608, g17520, I23611, g17523, I23619, g17531, I23622, g17534, I23625, g17537;
wire I23633, g17545, I23636, g17548, I23639, g17551, I23645, g17557, I23648, g17560, I23651;
wire g17563, g17566, I23655, g17567, I23658, g17570, I23661, g17573, I23667, g17579, I23670;
wire g17582, I23673, g17585, I23676, g17588, I23679, g17591, I23682, g17594, I23689, g17601;
wire I23692, g17604, I23695, g17607, I23698, g17610, I23701, g17613, I23709, g17621, I23712;
wire g17624, I23715, g17627, I23725, g17637, g17640, I23729, g17645, g17648, I23733, g17649;
wire I23739, g17655, I23742, g17658, I23745, g17661, I23748, g17664, I23751, g17667, I23754;
wire g17670, I23760, g17676, I23763, g17679, I23766, g17682, I23769, g17685, I23772, g17688;
wire I23775, g17691, I23782, g17698, I23785, g17701, I23788, g17704, I23791, g17707, I23794;
wire g17710, g17720, g17724, I23817, g17738, g17741, I23821, g17746, I23824, g17749, I23830;
wire g17755, I23833, g17758, I23836, g17761, I23839, g17764, I23842, g17767, I23845, g17770;
wire I23851, g17776, I23854, g17779, I23857, g17782, I23860, g17785, I23863, g17788, I23866;
wire g17791, I23874, g17799, g17802, I23888, g17815, g17825, I23904, g17839, g17842, I23908;
wire g17847, I23911, g17850, I23917, g17856, I23920, g17859, I23923, g17862, I23926, g17865;
wire I23929, g17868, I23932, g17871, g17878, g17882, g17892, g17893, I23954, g17903, g17914;
wire I23976, g17927, g17937, I23992, g17951, g17954, I23996, g17959, I23999, g17962, g17969;
wire g17974, g17984, g17988, g17991, g17993, g18003, g18004, I24049, g18014, g18025, I24071;
wire g18038, g18048, g18063, g18070, g18074, g18084, g18089, g18091, g18101, g18105, g18108;
wire g18110, g18120, g18121, I24144, g18131, g18142, I24166, g18155, I24171, g18166, g18170;
wire g18174, g18179, g18188, g18190, g18200, g18205, g18207, g18217, g18221, g18224, g18226;
wire g18236, g18237, I24247, g18247, I24258, g18258, g18261, g18265, g18275, I24285, g18278;
wire g18281, g18286, g18295, g18297, g18307, g18312, g18314, g18324, g18328, g18331, I24346;
wire g18334, g18337, g18341, g18351, g18353, I24368, g18355, g18358, g18368, I24394, g18371;
wire g18374, g18379, g18388, g18390, g18400, g18405, g18407, g18414, g18415, g18429, I24459;
wire g18432, g18435, g18436, g18446, g18448, I24481, g18450, g18453, g18463, I24507, g18466;
wire g18469, g18474, g18483, g18485, g18486, g18490, g18502, I24560, g18505, g18508, g18509;
wire g18519, g18521, I24582, g18523, g18526, g18536, I24608, g18539, g18543, g18552, g18554;
wire g18566, I24662, g18569, g18572, g18573, g18583, g18585, I24684, g18587, g18593, g18602;
wire g18604, g18616, I24732, g18619, g18622, g18634, g18636, g18643, g18646, g18656, g18670;
wire g18679, g18691, g18692, g18699, g18708, g18720, g18725, g18727, g18728, g18735, g18744;
wire g18756, g18757, g18758, g18764, g18765, g18772, g18783, g18784, g18785, g18786, g18787;
wire g18788, g18789, g18795, g18796, g18805, g18806, g18807, g18808, g18809, g18810, g18811;
wire g18812, g18813, g18814, g18815, g18822, g18823, g18824, g18825, g18826, g18827, g18828;
wire g18829, g18830, g18831, g18832, g18833, g18834, g18838, g18839, g18840, g18841, g18842;
wire g18843, g18844, g18845, g18846, g18847, g18848, g18849, g18850, g18851, g18853, g18854;
wire g18855, g18856, g18857, g18858, g18859, g18860, g18861, g18862, g18863, g18864, g18865;
wire I24894, g18869, g18870, g18871, g18872, g18873, g18874, g18875, g18876, g18877, g18878;
wire g18879, g18880, g18881, g18882, g18884, I24913, g18886, I24916, g18890, g18891, g18892;
wire g18893, g18894, I24923, g18895, g18896, g18897, g18898, g18899, g18900, g18901, g18902;
wire g18903, g18904, g18905, g18908, g18909, g18910, g18911, g18912, I24943, g18913, g18914;
wire g18915, g18916, g18917, I24950, g18918, g18919, g18920, g18921, g18922, g18923, g18924;
wire g18925, g18926, g18927, g18928, g18929, g18930, g18931, I24966, g18932, g18933, g18934;
wire g18935, g18936, I24973, g18937, g18938, g18939, g18940, g18941, g18943, I24982, g18944;
wire g18945, g18946, g18947, g18948, g18949, g18950, g18951, I24992, g18952, g18953, g18954;
wire g18955, g18956, g18958, I25001, g18959, I25004, g18960, g18961, g18962, g18963, g18964;
wire g18965, g18966, g18967, I25015, g18969, I25018, g18970, I25021, g18971, g18972, g18973;
wire g18974, g18976, I25037, g18981, I25041, g18983, I25044, g18984, I25047, g18985, I25050;
wire g18986, g18987, I25054, g18988, I25057, g18989, I25061, g18991, I25064, g18992, I25067;
wire g18993, I25071, g18995, I25074, g18996, I25078, g18998, I25081, g18999, I25084, g19000;
wire g19001, I25089, g19008, I25092, g19009, I25096, g19011, I25099, g19012, I25102, g19013;
wire I25105, g19014, I25108, g19015, I25111, g19016, I25114, g19017, I25117, g19018, I25120;
wire g19019, I25123, g19020, I25126, g19021, I25129, g19022, I25132, g19023, I25135, g19024;
wire I25138, g19025, I25141, g19026, I25144, g19027, I25147, g19028, I25150, g19029, I25153;
wire g19030, I25156, g19031, I25159, g19032, I25162, g19033, I25165, g19034, I25168, g19035;
wire I25171, g19036, I25174, g19037, I25177, g19038, I25180, g19039, I25183, g19040, I25186;
wire g19041, I25189, g19042, I25192, g19043, I25195, g19044, I25198, g19045, I25201, g19046;
wire I25204, g19047, I25207, g19048, I25210, g19049, I25213, g19050, I25216, g19051, I25219;
wire g19052, I25222, g19053, I25225, g19054, I25228, g19055, I25231, g19056, I25234, g19057;
wire I25237, g19058, I25240, g19059, I25243, g19060, I25246, g19061, I25249, g19062, I25253;
wire g19064, g19070, I25258, g19075, g19078, I25264, g19081, I25272, g19091, g19096, I25283;
wire g19098, I25294, g19105, I25303, g19110, I25308, g19113, I25315, g19118, I25320, g19125;
wire I25325, g19132, I25334, g19145, I25338, g19147, I25344, g19151, I25351, g19156, I25355;
wire g19158, I25358, g19159, I25365, g19164, I25371, g19168, I25374, g19169, I25377, g19170;
wire I25383, g19174, I25386, g19175, I25389, g19176, I25395, g19180, I25399, g19182, I25402;
wire g19183, I25406, g19185, I25412, g19189, I25415, g19190, I25423, g19196, I25426, g19197;
wire I25429, g19198, I25432, g19199, I25442, g19207, I25445, g19208, I25456, g19217, I25459;
wire g19218, I25463, g19220, I25474, g19229, I25486, g19237, I25489, g19238, I25492, g19239;
wire I25506, g19247, I25510, g19249, g19251, I25525, g19258, I25528, g19259, g19265, I25557;
wire g19270, I25567, g19272, g19280, g19287, I25612, g19291, g19299, g19301, g19302, g19305;
wire I25660, g19309, g19319, g19322, g19323, g19326, I25717, g19330, I25728, g19335, g19346;
wire g19349, g19350, g19353, I25768, g19358, I25778, g19369, g19380, g19383, g19384, g19387;
wire g19388, I25816, g19390, I25826, g19401, g19412, g19415, g19417, g19418, I25862, g19420;
wire I25872, g19431, g19441, g19444, g19448, g19452, g19454, g19455, I25904, g19457, g19467;
wire g19468, g19471, g19475, g19479, g19481, g19482, g19483, g19484, g19490, g19491, g19494;
wire g19498, g19502, g19504, g19505, g19511, g19512, g19515, g19519, g19523, g19524, g19530;
wire g19533, g19534, I25966, g19543, I25971, g19546, I25977, g19550, I25985, g19556, I25994;
wire g19563, I26006, g19573, g19577, g19578, I26025, g19595, I26028, g19596, g19607, g19608;
wire I26051, g19622, g19640, g19641, I26078, g19652, I26085, g19657, g19680, g19681, I26112;
wire g19689, I26115, g19690, I26123, g19696, I26134, g19705, I26154, g19725, I26171, g19740;
wire I26182, g19749, I26195, g19762, I26198, g19763, I26220, g19783, I26231, g19792, I26237;
wire g19798, I26266, g19825, g19830, I26276, g19838, I26334, g19890, I26337, g19893, I26340;
wire g19894, I26365, g19915, g19918, I26369, g19919, g19933, I26388, g19934, I26401, g19945;
wire g19948, g19950, I26407, g19951, I26413, g19957, I26420, g19972, g19975, g19977, I26426;
wire g19978, I26437, g19987, I26444, g20002, g20005, g20007, I26458, g20016, I26469, g20025;
wire I26476, g20040, g20043, I26481, g20045, I26494, g20058, I26505, g20067, I26512, g20082;
wire g20083, I26535, g20099, I26545, g20105, I26574, g20124, g20127, g20140, g20163, I26612;
wire g20164, g20178, g20193, I26642, g20198, g20212, g20223, I26664, g20228, g20242, g20250;
wire I26679, g20255, g20269, g20273, g20278, g20279, g20281, g20286, g20287, g20288, g20289;
wire g20290, g20292, I26714, g20295, g20296, g20297, g20298, g20302, g20303, g20304, g20305;
wire g20306, g20308, g20311, g20312, g20313, g20315, g20316, g20317, g20321, g20322, g20323;
wire g20324, g20325, g20327, g20328, g20329, g20330, g20331, g20332, g20334, g20335, g20336;
wire g20340, g20341, g20342, g20344, g20345, g20346, g20347, g20348, g20349, g20350, g20351;
wire g20352, g20354, g20355, g20356, I26777, g20360, g20361, g20362, g20363, g20364, g20365;
wire g20366, g20367, g20368, g20369, g20370, g20371, g20372, g20373, g20374, I26796, g20377;
wire g20378, g20379, g20380, g20381, g20382, g20383, g20384, g20385, g20386, g20387, g20388;
wire g20389, g20390, g20391, g20392, g20393, g20394, I26816, g20395, I26819, g20396, g20397;
wire g20398, g20399, g20400, g20401, g20402, g20403, g20404, g20405, g20406, g20407, g20408;
wire g20409, g20410, g20411, g20412, g20413, g20414, g20415, g20416, I26843, g20418, I26846;
wire g20419, g20420, g20421, g20422, g20423, g20424, g20425, g20426, g20427, g20428, g20429;
wire g20430, g20431, g20432, g20433, g20434, g20435, g20436, g20437, g20438, I26868, g20439;
wire I26871, g20440, I26874, g20441, g20442, g20443, g20444, g20445, g20446, g20447, g20448;
wire g20449, g20450, g20451, g20452, g20453, g20454, g20455, g20456, I26892, g20457, I26895;
wire g20458, I26898, g20459, g20461, g20462, g20463, g20464, g20465, g20466, g20467, g20468;
wire I26910, g20469, I26913, g20470, I26916, g20471, g20476, g20477, I26923, g20478, I26926;
wire g20479, I26931, g20484, I26934, g20485, g20490, I26940, g20491, g20496, I26947, g20498;
wire g20500, g20501, g20504, g20505, g20507, I26960, g20513, g20516, g20517, g20518, I26966;
wire g20519, g20526, I26972, g20531, g20534, g20535, g20536, I26980, g20539, g20545, I26985;
wire g20550, g20553, g20554, I26990, g20555, I26993, g20556, I26996, g20557, I26999, g20558;
wire I27002, g20559, I27005, g20560, I27008, g20561, I27011, g20562, I27014, g20563, I27017;
wire g20564, I27020, g20565, I27023, g20566, I27026, g20567, I27029, g20568, I27032, g20569;
wire I27035, g20570, I27038, g20571, I27041, g20572, I27044, g20573, I27047, g20574, I27050;
wire g20575, I27053, g20576, I27056, g20577, I27059, g20578, I27062, g20579, I27065, g20580;
wire I27068, g20581, I27071, g20582, I27074, g20583, I27077, g20584, I27080, g20585, I27083;
wire g20586, I27086, g20587, I27089, g20588, I27092, g20589, I27095, g20590, I27098, g20591;
wire I27101, g20592, I27104, g20593, I27107, g20594, I27110, g20595, I27113, g20596, I27116;
wire g20597, I27119, g20598, I27122, g20599, I27125, g20600, I27128, g20601, I27131, g20602;
wire I27134, g20603, I27137, g20604, I27140, g20605, I27143, g20606, I27146, g20607, I27149;
wire g20608, I27152, g20609, I27155, g20610, I27158, g20611, I27161, g20612, I27164, g20613;
wire I27167, g20614, I27170, g20615, I27173, g20616, I27176, g20617, I27179, g20618, I27182;
wire g20619, I27185, g20620, I27188, g20621, I27191, g20622, I27194, g20623, I27197, g20624;
wire I27200, g20625, I27203, g20626, I27206, g20627, I27209, g20628, I27212, g20629, I27215;
wire g20630, I27218, g20631, I27221, g20632, I27225, g20634, I27228, g20637, I27232, g20641;
wire I27235, g20644, I27240, g20649, I27243, g20652, I27246, g20655, I27250, g20659, I27253;
wire g20662, I27257, g20666, I27260, g20669, I27264, g20673, I27267, g20676, I27270, g20679;
wire I27275, g20684, I27278, g20687, I27281, g20690, I27285, g20694, I27288, g20697, I27293;
wire g20704, I27297, g20708, I27300, g20711, I27303, g20714, I27308, g20719, I27311, g20722;
wire I27314, g20725, I27318, g20729, I27321, g20732, I27324, g20735, I27328, g20739, I27332;
wire g20743, I27335, g20746, I27338, g20749, I27343, g20754, I27346, g20757, I27349, g20760;
wire I27352, g20763, I27355, g20766, I27358, g20769, I27361, g20772, I27365, g20776, I27369;
wire g20780, I27372, g20783, I27375, g20786, I27379, g20790, I27382, g20793, I27385, g20796;
wire I27388, g20799, I27391, g20802, I27395, g20806, I27399, g20810, I27402, g20813, I27405;
wire g20816, I27408, g20819, I27411, g20822, I27416, g20827, I27419, g20830, I27422, g20833;
wire I27426, g20837, g20842, g20850, g20858, g20866, g20885, g20904, g20928, I27488, g20942;
wire I27491, g20943, g20956, I27516, g20971, I27531, g20984, I27534, g20985, I27537, g20986;
wire I27549, g20998, I27565, g21012, I27577, g21024, I27585, g21030, I27593, g21036, g21050;
wire I27614, g21057, I27621, g21064, g21066, g21069, g21076, g21079, I27646, g21087, g21090;
wire g21093, I27658, g21099, g21102, I27667, g21108, I27672, g21113, I27684, g21125, I27689;
wire g21130, I27705, g21144, I27727, g21164, I27749, g21184, g21187, I27766, g21199, g21202;
wire I27779, g21214, g21217, I27785, g21222, g21225, g21241, g21249, g21258, g21266, I27822;
wire g21271, I27827, g21278, I27832, g21285, I27838, g21293, I27868, g21327, I27897, g21358;
wire I27900, g21359, I27917, g21376, I27920, g21377, I27927, g21382, I27942, g21399, g21400;
wire I27949, g21404, I27958, g21415, I27969, g21426, I27972, g21427, I27976, g21429, I27984;
wire g21441, I27992, g21449, I28000, g21457, I28003, g21458, g21461, I28009, g21473, I28013;
wire g21477, I28019, g21483, I28027, g21491, I28031, g21495, I28034, g21496, I28038, g21498;
wire I28043, g21505, g21508, I28047, g21514, I28051, g21518, I28057, g21524, I28061, g21528;
wire g21529, I28065, g21530, I28072, g21537, I28076, g21541, g21544, I28080, g21550, I28084;
wire g21554, I28087, g21557, I28090, g21558, I28093, g21561, g21565, I28100, g21566, I28107;
wire g21573, I28111, g21577, g21580, I28115, g21586, I28119, g21590, I28123, g21594, g21598;
wire I28130, g21599, I28137, g21606, I28143, g21612, I28148, g21619, I28152, g21623, g21627;
wire I28159, g21628, I28169, g21640, I28174, g21647, I28178, g21651, I28184, g21655, g21661;
wire I28201, g21671, I28206, g21678, I28210, g21682, g21690, I28229, g21700, I28235, g21708;
wire g21716, g21726, g21742, g21752, g21766, g21782, I28314, g21795, I28357, g21824, I28360;
wire g21825, g21861, g21867, g21872, g21876, g21883, g21886, g21895, g21902, g21907, I28432;
wire g21914, I28435, g21917, g21921, g21927, I28443, g21928, I28447, g21932, I28450, g21935;
wire g21939, I28455, g21943, I28458, g21944, I28461, g21945, I28464, g21946, I28467, g21947;
wire I28470, g21948, I28473, g21949, I28476, g21950, I28479, g21951, I28482, g21952, I28485;
wire g21953, I28488, g21954, I28491, g21955, I28494, g21956, I28497, g21957, I28500, g21958;
wire I28503, g21959, I28506, g21960, I28509, g21961, I28512, g21962, I28515, g21963, I28518;
wire g21964, I28521, g21965, I28524, g21966, I28527, g21967, I28541, g21982, I28550, g21995;
wire I28557, g22003, I28564, g22014, I28628, g22082, I28649, g22107, I28671, g22133, I28693;
wire g22156, I28712, g22176, g22212, g22213, g22217, I28781, g22219, g22221, g22222, I28789;
wire g22225, I28792, g22226, g22230, I28800, g22232, g22233, g22236, g22237, g22239, g22240;
wire g22241, I28813, g22243, g22246, g22248, g22251, g22252, I28825, g22253, g22256, g22257;
wire g22258, I28833, g22259, g22260, g22261, g22262, g22266, g22268, g22271, g22274, g22275;
wire g22276, g22277, g22278, g22279, g22283, g22286, g22287, g22290, g22293, g22294, g22295;
wire g22296, g22297, g22298, I28876, g22300, g22303, g22304, g22306, g22307, g22310, g22313;
wire g22314, g22315, g22316, g22318, g22319, I28896, g22328, g22331, g22332, g22334, g22335;
wire g22338, g22341, g22343, g22344, I28913, g22353, g22356, g22357, g22359, g22360, g22364;
wire g22366, g22367, I28928, g22376, g22379, g22380, g22384, g22386, g22387, g22401, g22402;
wire g22403, g22404, I28949, g22405, g22408, I28953, g22409, I28956, g22412, I28959, g22415;
wire I28962, g22418, g22421, I28966, g22422, I28969, g22425, I28972, g22428, I28975, g22431;
wire I28978, g22434, I28981, g22437, I28984, g22440, g22443, I28988, g22444, I28991, g22445;
wire I28994, g22448, I28997, g22451, I29001, g22455, I29004, g22458, I29007, g22461, I29010;
wire g22464, I29013, g22467, I29016, g22470, I29019, g22473, g22476, I29023, g22477, I29026;
wire g22480, I29030, g22484, I29033, g22487, I29036, g22490, I29040, g22494, I29043, g22497;
wire I29046, g22500, I29049, g22503, I29052, g22506, I29055, g22509, I29058, g22512, I29064;
wire g22518, I29067, g22519, I29070, g22520, I29073, g22523, I29077, g22527, I29080, g22530;
wire I29083, g22533, I29087, g22537, I29090, g22540, I29093, g22543, g22547, I29098, g22548;
wire I29101, g22549, I29104, g22550, I29107, g22551, I29110, g22552, I29116, g22558, I29119;
wire g22559, I29122, g22560, I29125, g22563, I29129, g22567, I29132, g22570, I29135, g22573;
wire I29142, g22582, I29145, g22583, I29148, g22584, I29151, g22585, I29154, g22586, g22588;
wire I29159, g22589, I29162, g22590, I29165, g22591, I29168, g22592, I29174, g22598, I29177;
wire g22599, I29180, g22600, I29183, g22603, g22609, I29191, g22611, I29194, g22612, I29197;
wire g22613, I29203, g22619, I29206, g22620, I29209, g22621, I29212, g22622, I29215, g22623;
wire g22625, I29220, g22626, I29223, g22627, I29226, g22628, I29229, g22629, I29235, g22635;
wire I29238, g22636, I29243, g22639, I29246, g22640, I29249, g22641, I29252, g22642, g22645;
wire I29259, g22647, I29262, g22648, I29265, g22649, I29271, g22655, I29274, g22656, I29277;
wire g22657, I29280, g22658, I29283, g22659, g22661, I29288, g22662, I29291, g22663, I29294;
wire g22664, I29301, g22669, I29304, g22670, I29307, g22671, I29310, g22672, I29313, g22673;
wire I29317, g22675, I29320, g22676, I29323, g22677, I29326, g22678, g22681, I29333, g22683;
wire I29336, g22684, I29339, g22685, I29345, g22691, I29348, g22692, I29351, g22693, I29354;
wire g22694, I29357, g22695, I29360, g22696, I29366, g22702, I29369, g22703, I29372, g22704;
wire I29375, g22705, I29378, g22706, I29383, g22709, I29386, g22710, I29389, g22711, I29392;
wire g22712, I29395, g22713, I29399, g22715, I29402, g22716, I29405, g22717, I29408, g22718;
wire g22721, I29415, g22723, I29418, g22724, I29421, g22725, I29426, g22728, I29429, g22729;
wire I29432, g22730, I29435, g22731, I29439, g22733, I29442, g22734, I29445, g22735, I29448;
wire g22736, I29451, g22737, I29456, g22740, I29459, g22741, I29462, g22742, I29465, g22743;
wire I29468, g22744, I29472, g22746, I29475, g22747, I29478, g22748, I29481, g22749, I29484;
wire g22750, g22753, I29490, g22756, I29493, g22757, I29496, g22758, I29500, g22760, I29503;
wire g22761, I29506, g22762, I29509, g22763, I29513, g22765, I29516, g22766, I29519, g22767;
wire I29522, g22768, I29525, g22769, I29530, g22772, I29533, g22773, I29536, g22774, I29539;
wire g22775, I29542, g22776, g22777, I29547, g22785, I29550, g22786, g22787, I29556, g22790;
wire I29559, g22791, I29562, g22792, I29566, g22794, I29569, g22795, I29572, g22796, I29575;
wire g22797, I29579, g22799, I29582, g22800, I29585, g22801, I29588, g22802, I29591, g22803;
wire g22805, g22806, I29600, g22812, I29603, g22824, I29606, g22825, I29610, g22827, I29613;
wire g22828, g22829, I29619, g22832, I29622, g22833, I29625, g22834, I29629, g22836, I29632;
wire g22837, I29635, g22838, I29638, g22839, I29641, g22840, g22843, g22847, I29653, g22852;
wire I29656, g22864, I29660, g22866, I29663, g22867, g22868, I29669, g22871, I29672, g22872;
wire I29675, g22873, g22875, g22882, I29687, g22887, I29690, g22899, I29694, g22901, I29697;
wire g22902, I29700, g22903, g22907, g22917, I29712, g22922, I29715, g22934, I29724, g22945;
wire I29727, g22948, g22949, g22954, g22958, g22962, g22966, I29736, g22970, g22971, g22975;
wire I29741, g22979, g22980, g22986, g22988, g22989, g22991, g22995, g22996, g22998, g23001;
wire g23002, g23006, g23007, g23008, g23012, g23015, g23016, g23020, g23021, g23024, g23028;
wire g23031, g23032, g23036, g23037, g23038, g23041, g23045, g23048, g23049, I29797, g23050;
wire I29802, g23055, g23056, g23057, g23060, g23064, I29812, g23065, I29817, g23068, g23069;
wire g23074, g23075, I29827, g23078, g23079, g23082, g23087, g23088, I29841, g23094, g23095;
wire g23098, g23103, I29852, g23105, g23112, g23115, I29863, g23116, I29872, g23125, I29881;
wire g23134, g23140, g23141, g23142, g23143, g23144, g23145, g23146, g23147, I29897, g23148;
wire I29900, g23149, I29903, g23150, I29906, g23151, I29909, g23152, I29912, g23153, I29915;
wire g23154, I29918, g23155, I29921, g23156, I29924, g23157, I29927, g23158, I29930, g23159;
wire I29933, g23160, I29936, g23161, I29939, g23162, I29942, g23163, I29945, g23164, I29948;
wire g23165, I29951, g23166, I29954, g23167, I29957, g23168, I29960, g23169, I29963, g23170;
wire I29966, g23171, I29969, g23172, I29972, g23173, I29975, g23174, I29978, g23175, I29981;
wire g23176, I29984, g23177, I29987, g23178, I29990, g23179, I29993, g23180, I29996, g23181;
wire I29999, g23182, I30002, g23183, I30005, g23184, I30008, g23185, I30011, g23186, I30014;
wire g23187, I30017, g23188, I30020, g23189, I30023, g23190, I30026, g23191, I30029, g23192;
wire I30032, g23193, I30035, g23194, I30038, g23195, I30041, g23196, I30044, g23197, I30047;
wire g23198, I30050, g23199, I30053, g23200, I30056, g23201, I30059, g23202, I30062, g23203;
wire I30065, g23204, I30068, g23205, I30071, g23206, I30074, g23207, I30077, g23208, I30080;
wire g23209, I30083, g23210, I30086, g23211, I30089, g23212, I30092, g23213, I30095, g23214;
wire I30098, g23215, I30101, g23216, I30104, g23217, I30107, g23218, I30110, g23219, I30113;
wire g23220, I30116, g23221, I30119, g23222, I30122, g23223, I30125, g23224, I30128, g23225;
wire I30131, g23226, I30134, g23227, I30137, g23228, I30140, g23229, I30143, g23230, I30146;
wire g23231, I30149, g23232, I30152, g23233, I30155, g23234, I30158, g23235, I30161, g23236;
wire I30164, g23237, I30167, g23238, I30170, g23239, I30173, g23240, I30176, g23241, I30179;
wire g23242, I30182, g23243, I30185, g23244, I30188, g23245, I30191, g23246, I30194, g23247;
wire I30197, g23248, I30200, g23249, I30203, g23250, I30206, g23251, I30209, g23252, I30212;
wire g23253, I30215, g23254, I30218, g23255, I30221, g23256, I30224, g23257, I30227, g23258;
wire I30230, g23259, I30233, g23260, I30236, g23261, I30239, g23262, I30242, g23263, I30245;
wire g23264, I30248, g23265, I30251, g23266, I30254, g23267, I30257, g23268, I30260, g23269;
wire I30263, g23270, I30266, g23271, I30269, g23272, I30272, g23273, I30275, g23274, I30278;
wire g23275, I30281, g23276, I30284, g23277, I30287, g23278, I30290, g23279, I30293, g23280;
wire I30296, g23281, I30299, g23282, I30302, g23283, I30305, g23284, I30308, g23285, I30311;
wire g23286, I30314, g23287, I30317, g23288, I30320, g23289, I30323, g23290, I30326, g23291;
wire I30329, g23292, I30332, g23293, I30335, g23294, I30338, g23295, I30341, g23296, I30344;
wire g23297, I30347, g23298, I30350, g23299, I30353, g23300, I30356, g23301, I30359, g23302;
wire I30362, g23303, I30365, g23304, I30368, g23305, I30371, g23306, I30374, g23307, I30377;
wire g23308, I30380, g23309, I30383, g23310, I30386, g23311, I30389, g23312, I30392, g23313;
wire I30395, g23314, I30398, g23315, I30401, g23316, I30404, g23317, I30407, g23318, g23403;
wire g23410, g23415, g23420, g23424, g23429, g23435, I30467, g23438, I30470, g23439, g23441;
wire g23444, I30476, g23448, I30480, g23452, I30483, g23453, I30486, g23454, I30489, g23455;
wire I30493, g23459, I30496, g23460, I30501, g23463, I30504, g23464, I30508, g23468, I30511;
wire g23469, g23470, I30516, g23472, I30519, g23473, I30525, g23481, g23482, I30531, g23485;
wire I30536, g23492, g23493, I30544, g23500, I30547, g23501, I30552, g23508, g23509, I30560;
wire g23516, I30563, g23517, I30568, g23524, I30575, g23531, I30578, g23532, I30586, g23542;
wire I30589, g23543, I30594, g23546, I30598, g23548, I30601, g23549, I30607, g23553, I30611;
wire g23555, I30614, g23556, I30617, g23557, I30623, g23561, I30626, g23562, I30632, g23566;
wire I30636, g23568, I30639, g23569, I30642, g23570, I30648, g23574, I30651, g23575, I30654;
wire g23576, I30660, g23580, I30663, g23581, I30669, g23585, I30673, g23587, I30676, g23588;
wire I30679, g23589, I30686, g23594, I30689, g23595, I30692, g23596, I30695, g23597, I30701;
wire g23601, I30704, g23602, I30707, g23603, I30713, g23607, I30716, g23608, I30722, g23612;
wire I30725, g23613, I30728, g23614, I30735, g23619, I30738, g23620, I30741, g23621, I30748;
wire g23626, I30751, g23627, I30754, g23628, I30757, g23629, I30763, g23633, I30766, g23634;
wire I30769, g23635, I30776, g23640, I30779, g23641, I30782, g23642, I30786, g23644, I30797;
wire g23661, I30800, g23662, I30803, g23663, I30810, g23668, I30813, g23669, I30816, g23670;
wire I30823, g23675, I30826, g23676, I30829, g23677, I30832, g23678, I30838, g23682, I30841;
wire g23683, I30844, g23684, I30847, g23685, I30854, g23690, I30857, g23691, I30860, g23692;
wire I30864, g23694, I30875, g23711, I30878, g23712, I30881, g23713, I30888, g23718, I30891;
wire g23719, I30894, g23720, I30901, g23725, I30905, g23727, I30908, g23728, I30911, g23729;
wire I30914, g23730, I30917, g23731, I30922, g23736, I30925, g23737, I30928, g23738, I30931;
wire g23739, I30938, g23744, I30941, g23745, I30944, g23746, I30948, g23748, I30959, g23765;
wire I30962, g23766, I30965, g23767, I30973, g23773, I30976, g23774, I30979, g23775, I30985;
wire g23779, I30988, g23782, I30991, g23783, I30994, g23784, I30997, g23785, I31000, g23786;
wire I31005, g23791, I31008, g23792, I31011, g23793, I31014, g23794, I31021, g23799, I31024;
wire g23800, I31027, g23801, I31031, g23803, I31043, g23821, I31050, g23826, I31053, g23827;
wire I31056, g23828, I31062, g23832, I31065, g23835, I31068, g23836, I31071, g23837, I31074;
wire g23838, I31077, g23839, I31082, g23844, I31085, g23845, I31088, g23846, I31091, g23847;
wire g23853, I31102, g23856, I31109, g23861, I31112, g23862, I31115, g23863, I31121, g23867;
wire I31124, g23870, I31127, g23871, I31130, g23872, I31133, g23873, I31136, g23874, I31141;
wire g23879, I31144, g23882, g23885, g23887, I31152, g23890, I31159, g23895, I31162, g23896;
wire I31165, g23897, I31171, g23901, g23905, g23908, I31181, g23911, I31188, g23916, g23918;
wire I31195, g23923, g23940, I31205, g23943, I31213, g23955, I31226, g23984, I31232, g24000;
wire I31235, g24001, I31244, g24014, I31250, g24030, I31253, g24033, I31257, g24035, g24047;
wire I31266, g24051, I31270, g24053, I31274, g24055, g24060, I31282, g24064, I31286, g24066;
wire I31290, g24068, g24073, I31298, g24077, I31302, g24079, g24084, I31310, g24088, g24094;
wire g24095, g24096, g24097, g24098, g24099, g24101, g24102, g24103, g24104, g24105, g24106;
wire g24107, g24108, g24110, g24111, g24112, g24113, g24114, g24115, g24121, g24122, g24123;
wire g24124, g24125, g24127, g24128, g24129, g24130, g24131, g24132, g24133, g24134, g24140;
wire g24141, g24142, g24143, g24144, g24146, g24147, g24148, g24149, g24150, g24151, g24152;
wire g24153, g24159, g24160, g24161, g24162, g24163, g24164, g24165, g24166, g24167, g24168;
wire g24175, g24176, g24177, g24180, I31387, g24183, g24210, g24220, I31417, g24233, I31426;
wire g24240, I31436, g24248, g24251, I31445, g24255, I31451, g24259, I31454, g24260, I31457;
wire g24261, I31460, g24262, I31463, g24263, I31466, g24264, I31469, g24265, I31472, g24266;
wire I31475, g24267, I31478, g24268, I31481, g24269, I31484, g24270, I31487, g24271, I31490;
wire g24272, I31493, g24273, I31496, g24274, I31499, g24275, I31502, g24276, I31505, g24277;
wire I31508, g24278, I31511, g24279, I31514, g24280, I31517, g24281, I31520, g24282, I31523;
wire g24283, I31526, g24284, I31529, g24285, I31532, g24286, I31535, g24287, I31538, g24288;
wire I31541, g24289, I31544, g24290, I31547, g24291, I31550, g24292, I31553, g24293, I31556;
wire g24294, I31559, g24295, I31562, g24296, I31565, g24297, I31568, g24298, I31571, g24299;
wire I31574, g24300, I31577, g24301, I31580, g24302, I31583, g24303, I31586, g24304, I31589;
wire g24305, I31592, g24306, I31595, g24307, I31598, g24308, I31601, g24309, I31604, g24310;
wire I31607, g24311, I31610, g24312, I31613, g24313, I31616, g24314, I31619, g24315, I31622;
wire g24316, I31625, g24317, I31628, g24318, I31631, g24319, I31634, g24320, I31637, g24321;
wire I31640, g24322, I31643, g24323, I31646, g24324, I31649, g24325, I31652, g24326, I31655;
wire g24327, I31658, g24328, I31661, g24329, I31664, g24330, I31667, g24331, I31670, g24332;
wire I31673, g24333, I31676, g24334, I31679, g24335, I31682, g24336, I31685, g24337, I31688;
wire g24338, I31691, g24339, I31694, g24340, I31697, g24341, I31700, g24342, I31703, g24343;
wire I31706, g24344, I31709, g24345, I31712, g24346, I31715, g24347, I31718, g24348, I31721;
wire g24349, I31724, g24350, I31727, g24351, I31730, g24352, I31733, g24353, I31736, g24354;
wire I31739, g24355, I31742, g24356, I31745, g24357, I31748, g24358, I31751, g24359, I31754;
wire g24360, I31757, g24361, I31760, g24362, I31763, g24363, I31766, g24364, I31769, g24365;
wire I31772, g24366, I31775, g24367, I31778, g24368, I31781, g24369, I31784, g24370, I31787;
wire g24371, I31790, g24372, I31793, g24373, I31796, g24374, I31799, g24375, I31802, g24376;
wire I31805, g24377, I31808, g24378, I31811, g24379, I31814, g24380, I31817, g24381, I31820;
wire g24382, I31823, g24383, I31826, g24384, I31829, g24385, I31832, g24386, I31835, g24387;
wire I31838, g24388, I31841, g24389, I31844, g24390, I31847, g24391, I31850, g24392, I31853;
wire g24393, I31856, g24394, I31859, g24395, I31862, g24396, I31865, g24397, I31868, g24398;
wire I31871, g24399, I31874, g24400, I31877, g24401, I31880, g24402, I31883, g24403, I31886;
wire g24404, I31889, g24405, I31892, g24406, I31895, g24407, I31898, g24408, I31901, g24409;
wire I31904, g24410, I31907, g24411, I31910, g24412, I31913, g24413, I31916, g24414, I31919;
wire g24415, I31922, g24416, I31925, g24417, I31928, g24418, I31931, g24419, I31934, g24420;
wire I31937, g24421, I31940, g24422, I31943, g24423, I31946, g24424, I31949, g24425, g24482;
wire I32042, g24518, I32057, g24531, I32067, g24539, I32074, g24544, I32081, g24549, I32085;
wire g24551, I32092, g24556, I32098, g24560, I32102, g24562, I32109, g24567, I32112, g24568;
wire I32116, g24570, I32120, g24572, I32126, g24576, I32129, g24577, I32133, g24579, I32137;
wire g24581, I32140, g24582, I32143, g24583, I32146, g24584, I32150, g24586, I32153, g24587;
wire I32156, g24588, I32159, g24589, I32164, g24592, I32167, g24593, I32170, g24594, I32175;
wire g24597, I32178, g24598, I32181, g24599, I32184, g24600, I32189, g24605, I32193, g24607;
wire I32198, g24612, I32203, g24619, I32210, g24630, g24648, g24668, g24687, g24704, I32248;
wire g24734, I32251, g24735, I32281, g24763, I32320, g24784, I32365, g24805, g24815, I32388;
wire g24816, I32419, g24827, g24834, I32439, g24835, g24850, I32487, g24851, I32506, g24856;
wire g24864, I32535, g24865, I32556, g24872, I32583, g24879, I32604, g24886, g24893, I32642;
wire g24903, g24912, g24916, g24929, g24933, g24939, g24941, g24945, I32704, g24949, g24950;
wire g24952, I32716, g24956, I32719, g24957, g24958, g24962, g24969, g24973, g24982, g24993;
wire g25087, g25094, g25095, I32829, g25103, g25104, g25105, I32835, g25109, g25110, g25111;
wire g25115, g25116, I32844, g25118, I32847, g25119, g25120, I32851, g25121, I32854, g25122;
wire I32857, g25123, I32860, g25124, g25126, I32868, g25130, I32871, g25131, I32874, g25132;
wire I32877, g25133, I32880, g25134, I32883, g25135, I32886, g25136, I32889, g25137, I32892;
wire g25138, I32895, g25139, I32898, g25140, I32901, g25141, I32904, g25142, I32907, g25143;
wire I32910, g25144, I32913, g25145, I32916, g25146, I32919, g25147, I32922, g25148, I32925;
wire g25149, I32928, g25150, I32931, g25151, I32934, g25152, I32937, g25153, I32940, g25154;
wire I32943, g25155, I32946, g25156, I32949, g25157, I32952, g25158, I32955, g25159, I32958;
wire g25160, I32961, g25161, I32964, g25162, I32967, g25163, I32970, g25164, I32973, g25165;
wire I32976, g25166, I32979, g25167, I32982, g25168, I32985, g25169, I32988, g25170, I32991;
wire g25171, I32994, g25172, I32997, g25173, I33000, g25174, I33003, g25175, I33006, g25176;
wire I33009, g25177, I33013, g25179, I33016, g25180, g25274, g25283, g25291, I33128, g25296;
wire g25301, g25305, I33136, g25306, g25313, g25314, I33145, g25315, g25319, g25322, g25323;
wire I33154, g25324, I33157, g25327, g25329, g25330, g25332, g25333, g25335, I33168, g25336;
wire g25338, g25339, g25341, g25347, g25349, I33182, g25350, g25352, g25353, I33188, g25354;
wire g25355, g25361, g25363, I33198, g25364, g25366, g25367, g25368, I33205, g25369, g25370;
wire g25376, g25378, g25379, g25383, g25384, g25385, I33219, g25386, g25387, g25393, g25394;
wire g25395, g25399, g25400, g25401, I33232, g25402, g25403, g25404, g25405, g25409, g25410;
wire g25411, g25412, g25413, g25417, g25419, I33246, g25420, I33249, g25421, g25422, g25430;
wire g25431, I33257, g25435, I33260, g25436, g25437, g25438, I33265, g25442, I33268, g25443;
wire g25444, g25445, g25449, I33278, g25454, I33282, g25458, I33286, g25462, I33289, g25463;
wire I33293, g25467, I33297, g25471, I33300, g25472, I33304, g25476, I33307, g25479, I33312;
wire g25484, I33316, g25488, I33321, g25493, I33324, g25496, I33327, g25499, I33330, g25502;
wire I33335, g25507, I33338, g25510, I33343, g25515, I33347, g25519, I33352, g25524, I33355;
wire g25527, I33358, g25530, I33361, g25533, I33364, g25536, I33368, g25540, I33371, g25543;
wire I33374, g25546, I33377, g25549, I33382, g25554, I33385, g25557, I33390, g25562, I33396;
wire g25573, I33399, g25576, I33402, g25579, I33405, g25582, I33408, g25585, I33411, g25588;
wire I33415, g25590, I33418, g25593, I33421, g25596, I33424, g25599, I33427, g25602, I33431;
wire g25606, I33434, g25609, I33437, g25612, I33440, g25615, I33445, g25620, I33448, g25623;
wire g25630, I33457, g25634, I33460, g25637, I33463, g25640, I33466, g25643, I33469, g25646;
wire I33472, g25647, I33476, g25652, I33479, g25655, I33482, g25658, I33485, g25661, I33488;
wire g25664, I33491, g25667, I33495, g25669, I33498, g25672, I33501, g25675, I33504, g25678;
wire I33507, g25681, I33511, g25685, I33514, g25688, I33517, g25691, I33520, g25694, g25698;
wire I33526, g25700, I33529, g25703, I33532, g25706, I33535, g25707, I33539, g25711, I33542;
wire g25714, I33545, g25717, I33548, g25720, I33551, g25723, I33554, g25724, I33558, g25729;
wire I33561, g25732, I33564, g25735, I33567, g25738, I33570, g25741, I33573, g25744, I33577;
wire g25746, I33580, g25749, I33583, g25752, I33586, g25755, I33589, g25758, I33593, g25762;
wire I33596, g25763, I33600, g25767, I33603, g25770, g25771, I33608, g25773, I33611, g25776;
wire I33614, g25779, I33617, g25780, I33621, g25784, I33624, g25787, I33627, g25790, I33630;
wire g25793, I33633, g25796, I33636, g25797, I33640, g25802, I33643, g25805, I33646, g25808;
wire I33649, g25811, I33652, g25814, I33655, g25817, I33659, g25821, I33662, g25824, g25825;
wire I33667, g25827, I33670, g25830, I33673, g25833, I33676, g25834, I33680, g25838, I33683;
wire g25841, I33686, g25844, I33689, g25847, I33692, g25850, I33695, g25851, I33700, g25856;
wire I33703, g25859, g25860, I33708, g25862, I33711, g25865, I33714, g25868, I33717, g25869;
wire I33723, g25877, I33726, g25880, I33732, g25886, I33737, g25891, g25895, g25899, g25903;
wire g25907, g25911, g25915, g25919, g25923, g25937, g25939, g25942, g25945, g25952, I33790;
wire g25976, I33798, g25982, I33801, g25983, I33804, g25984, I33807, g25985, I33810, g25986;
wire I33813, g25987, I33816, g25988, I33819, g25989, I33822, g25990, I33825, g25991, I33828;
wire g25992, I33831, g25993, I33834, g25994, I33837, g25995, I33840, g25996, I33843, g25997;
wire I33846, g25998, I33849, g25999, I33852, g26000, I33855, g26001, I33858, g26002, I33861;
wire g26003, I33864, g26004, I33867, g26005, I33870, g26006, I33873, g26007, I33876, g26008;
wire I33879, g26009, I33882, g26010, I33885, g26011, I33888, g26012, I33891, g26013, I33894;
wire g26014, I33897, g26015, I33900, g26016, I33903, g26017, I33906, g26018, I33909, g26019;
wire I33912, g26020, I33915, g26021, I33918, g26022, I33954, g26056, I33961, g26063, I33968;
wire g26070, I33974, g26076, I33984, g26086, I33990, g26092, I33995, g26102, I33999, g26104;
wire I34002, g26105, I34009, g26114, I34012, g26118, I34017, g26121, I34020, g26125, I34026;
wire g26131, I34029, g26135, I34032, g26136, I34041, g26149, I34044, g26150, I34051, g26159;
wire I34056, g26164, I34059, g26165, I34063, g26167, I34068, g26172, I34071, g26173, I34074;
wire g26174, I34077, g26175, I34080, g26178, I34083, g26181, I34086, g26182, I34091, g26187;
wire g26189, I34096, g26190, I34099, g26191, I34102, g26192, I34105, g26193, I34108, g26194;
wire I34111, g26195, I34114, g26196, I34118, g26202, I34121, g26205, I34124, g26206, I34128;
wire g26208, g26209, I34132, g26210, I34135, g26211, I34140, g26214, I34143, g26215, I34146;
wire g26216, I34150, g26220, I34153, g26221, I34156, g26222, I34159, g26223, I34162, g26226;
wire I34165, g26229, I34168, g26230, I34172, g26232, g26237, I34180, g26238, I34183, g26239;
wire I34189, g26245, I34192, g26246, I34195, g26247, I34198, g26248, I34201, g26249, I34204;
wire g26250, I34207, g26251, I34210, g26254, I34220, g26264, g26275, I34230, g26276, I34233;
wire g26277, I34238, g26280, I34241, g26281, I34244, g26282, I34254, g26294, I34266, g26308;
wire g26313, I34274, g26314, I34277, g26315, I34296, g26341, I34306, g26349, I34313, g26354;
wire I34316, g26355, I34321, g26358, I34327, g26364, I34343, g26385, I34353, g26393, I34358;
wire g26398, I34363, g26401, I34369, g26407, I34385, g26428, I34388, g26429, I34392, g26433;
wire I34395, g26434, I34400, g26439, I34405, g26442, I34411, g26448, I34421, g26461, I34425;
wire g26465, I34428, g26466, I34433, g26471, I34438, g26474, I34444, g26480, g26481, I34449;
wire g26485, I34453, g26489, I34456, g26490, I34461, g26495, I34464, g26496, g26497, I34469;
wire g26501, I34473, g26505, I34476, g26506, I34479, g26507, g26508, g26512, g26516, g26520;
wire g26521, g26525, g26533, g26538, g26539, g26540, g26542, g26543, g26544, g26546, I34505;
wire g26548, g26549, g26550, g26551, g26552, g26554, g26555, g26556, g26558, g26561, g26562;
wire g26563, g26564, g26565, g26566, g26567, g26568, g26570, g26571, g26572, g26574, I34535;
wire g26576, g26577, g26578, g26579, g26580, g26581, g26582, g26584, g26585, g26586, g26587;
wire g26588, g26589, g26590, g26591, g26593, g26594, g26595, g26597, g26598, g26599, g26600;
wire g26601, g26602, g26603, g26604, g26605, g26606, g26608, g26609, g26610, g26611, g26612;
wire g26613, g26614, g26615, g26617, I34579, g26618, g26619, g26620, g26621, g26622, g26623;
wire g26624, g26625, g26626, g26627, g26628, g26629, g26631, g26632, g26633, g26634, g26635;
wire g26636, g26637, g26638, g26639, g26640, g26641, g26642, g26643, g26644, g26645, g26646;
wire g26647, g26648, g26649, g26650, g26651, g26652, g26653, g26654, g26656, g26657, g26658;
wire g26662, I34641, g26678, I34644, g26679, I34647, g26680, I34650, g26681, I34653, g26682;
wire I34656, g26683, I34659, g26684, I34662, g26685, I34665, g26686, I34668, g26687, I34671;
wire g26688, I34674, g26689, I34677, g26690, I34680, g26691, I34683, g26692, I34686, g26693;
wire I34689, g26694, I34692, g26695, I34695, g26696, I34698, g26697, I34701, g26698, I34704;
wire g26699, I34707, g26700, I34710, g26701, I34713, g26702, I34716, g26703, I34719, g26704;
wire I34722, g26705, I34725, g26706, I34728, g26707, I34731, g26708, I34734, g26709, I34737;
wire g26710, I34740, g26711, I34743, g26712, I34746, g26713, I34749, g26714, I34752, g26715;
wire I34755, g26716, I34758, g26717, I34761, g26718, I34764, g26719, I34767, g26720, I34770;
wire g26721, I34773, g26722, I34776, g26723, I34779, g26724, I34782, g26725, I34785, g26726;
wire I34788, g26727, I34791, g26728, I34794, g26729, I34797, g26730, I34800, g26731, I34803;
wire g26732, I34806, g26733, I34809, g26734, I34812, g26735, I34815, g26736, I34818, g26737;
wire I34821, g26738, I34824, g26739, I34827, g26740, I34830, g26741, I34833, g26742, I34836;
wire g26743, I34839, g26744, I34842, g26745, I34845, g26746, I34848, g26747, I34851, g26748;
wire I34854, g26749, I34857, g26750, I34860, g26751, I34863, g26752, I34866, g26753, I34872;
wire g26757, I34879, g26762, I34901, g26782, I34909, g26788, I34916, g26793, I34921, g26796;
wire I34946, g26819, I34957, g26828, I34961, g26830, I34964, g26831, I34967, g26832, I34971;
wire g26834, I34974, g26835, I34977, g26836, I34980, g26837, I34983, g26840, I34986, g26841;
wire I34990, g26843, I34993, g26844, I34997, g26846, I35000, g26849, I35003, g26850, I35007;
wire g26852, I35011, g26854, I35014, g26855, I35017, g26858, I35028, g26861, I35031, g26864;
wire I35049, g26868, I35053, g26872, I35064, g26875, I35067, g26876, I35072, g26881, I35076;
wire g26883, I35079, g26884, I35083, g26886, I35087, g26890, I35092, g26895, I35095, g26896;
wire I35099, g26900, I35106, g26909, I35109, g26910, I35116, g26921, g26922, g26935, g26944;
wire g26950, I35136, g26953, g26954, I35141, g26956, g26957, I35146, g26959, g26960, I35153;
wire g26964, I35172, g26983, g26987, g27010, g27036, g27064, I35254, g27075, I35283, g27102;
wire I35297, g27114, I35301, g27116, I35313, g27126, I35319, g27132, g27133, g27134, g27135;
wire g27136, g27137, g27138, g27139, g27140, g27141, g27142, g27143, I35334, g27145, g27146;
wire g27148, I35341, g27150, g27151, g27153, I35347, g27154, g27155, I35351, g27156, I35355;
wire g27158, g27159, I35360, g27161, g27162, I35364, g27163, g27164, I35369, g27166, g27167;
wire I35373, g27168, I35376, g27171, g27172, g27173, I35383, g27176, g27177, I35389, g27180;
wire I35394, g27183, I35399, g27186, I35404, g27189, I35407, g27190, I35410, g27191, I35413;
wire g27192, I35416, g27193, I35419, g27194, I35422, g27195, I35425, g27196, I35428, g27197;
wire I35431, g27198, I35434, g27199, I35437, g27200, I35440, g27201, I35443, g27202, I35446;
wire g27203, I35449, g27204, I35452, g27205, I35455, g27206, I35458, g27207, I35461, g27208;
wire I35464, g27209, I35467, g27210, I35470, g27211, I35473, g27212, I35476, g27213, I35479;
wire g27214, I35482, g27215, I35485, g27216, I35488, g27217, I35491, g27218, I35494, g27219;
wire I35497, g27220, I35500, g27221, I35503, g27222, I35506, g27223, I35509, g27224, I35512;
wire g27225, I35515, g27226, I35518, g27227, I35521, g27228, I35524, g27229, I35527, g27230;
wire I35530, g27231, I35533, g27232, I35536, g27233, I35539, g27234, I35542, g27235, I35545;
wire g27236, I35548, g27237, I35551, g27238, I35554, g27239, g27349, I35667, g27353, I35673;
wire g27357, I35678, g27360, I35681, g27361, I35686, g27366, I35689, g27367, I35695, g27373;
wire I35698, g27376, I35708, g27380, I35711, g27381, g27383, g27384, I35723, g27385, g27386;
wire I35727, g27387, I35731, g27391, I35737, g27397, I35741, g27401, I35744, g27404, I35750;
wire g27410, I35756, g27416, I35759, g27419, I35762, g27422, I35768, g27428, I35772, g27432;
wire I35777, g27437, I35780, g27440, I35783, g27443, g27449, I35791, g27451, I35796, g27456;
wire I35799, g27459, I35803, g27463, g27465, I35809, g27467, I35814, g27472, I35817, g27475;
wire I35821, g27479, I35824, g27480, I35829, g27483, g27484, I35834, g27486, I35837, g27489;
wire I35841, g27493, I35844, g27494, I35849, g27497, I35852, g27498, I35856, g27502, I35859;
wire g27503, I35863, g27505, g27506, I35868, g27508, I35872, g27510, I35876, g27514, I35879;
wire g27515, I35883, g27517, I35886, g27518, I35890, g27522, I35893, g27523, I35897, g27525;
wire I35900, g27526, I35915, g27533, I35919, g27535, I35923, g27539, I35926, g27540, I35930;
wire g27542, I35933, g27543, I35937, g27547, I35940, g27548, I35953, g27553, I35957, g27555;
wire I35961, g27559, I35964, g27560, I35968, g27562, I35983, g27569, I36008, g27586, g27589;
wire g27590, g27595, g27599, g27604, g27608, g27613, g27617, g27622, I36032, g27632, I36042;
wire g27662, I36046, g27667, I36052, g27674, I36060, g27683, I36063, g27684, I36066, g27685;
wire I36069, g27686, I36072, g27687, I36075, g27688, I36078, g27689, I36081, g27690, I36084;
wire g27691, I36087, g27692, I36090, g27693, I36093, g27694, I36096, g27695, I36099, g27696;
wire I36102, g27697, I36105, g27698, I36108, g27699, I36111, g27700, I36114, g27701, I36117;
wire g27702, I36120, g27703, I36123, g27704, I36126, g27705, I36129, g27706, I36132, g27707;
wire I36135, g27708, I36138, g27709, I36141, g27710, I36144, g27711, I36147, g27712, I36150;
wire g27713, I36153, g27714, I36156, g27715, I36159, g27716, I36162, g27717, g27748, I36213;
wire g27776, I36217, g27780, I36221, g27784, I36224, g27785, I36227, g27786, I36230, g27787;
wire I36234, g27791, I36237, g27792, I36240, g27793, I36243, g27794, I36246, g27797, I36250;
wire g27799, I36253, g27800, I36264, g27805, I36267, g27806, I36280, g27817, I36283, g27820;
wire I36296, g27831, I36307, g27839, I36311, g27843, I36321, g27847, I36327, g27858, I36330;
wire g27861, I36337, g27872, I36341, g27879, I36347, g27889, I36354, g27903, I36358, g27905;
wire I36362, g27907, I36367, g27910, I36371, g27912, I36379, g27918, I36382, g27919, I36390;
wire g27927, I36393, g27928, I36397, g27932, I36404, g27939, I36407, g27942, I36411, g27946;
wire I36417, g27952, I36420, g27955, I36423, g27956, I36426, g27959, I36432, g27965, g27969;
wire I36438, g27971, I36441, g27972, I36444, g27973, I36447, g27976, I36450, g27977, I36454;
wire g27981, I36459, g27986, I36462, g27987, I36465, g27988, I36468, g27989, g27990, I36473;
wire g27992, I36476, g27993, I36479, g27994, I36483, g27998, I36486, g27999, I36490, g28003;
wire I36493, g28004, I36496, g28005, I36499, g28006, I36502, g28007, I36507, g28010, I36510;
wire g28011, I36513, g28012, I36516, g28013, g28014, I36521, g28016, I36524, g28017, I36527;
wire g28018, I36530, g28021, I36533, g28022, I36536, g28023, I36539, g28024, I36542, g28025;
wire I36545, g28026, I36551, g28030, I36554, g28031, I36557, g28032, I36560, g28033, I36563;
wire g28034, I36568, g28037, I36571, g28038, I36574, g28039, I36577, g28040, g28041, I36582;
wire g28043, I36585, g28044, I36588, g28045, I36598, g28047, I36601, g28048, I36604, g28049;
wire I36609, g28052, I36612, g28053, I36615, g28054, I36618, g28055, I36621, g28056, I36627;
wire g28060, I36630, g28061, I36633, g28062, I36636, g28063, I36639, g28064, I36644, g28067;
wire I36647, g28068, I36650, g28069, I36653, g28070, I36656, g28071, I36659, g28072, I36663;
wire g28074, I36673, g28076, I36676, g28077, I36679, g28078, I36684, g28081, I36687, g28082;
wire I36690, g28083, I36693, g28084, I36696, g28085, I36702, g28089, I36705, g28090, I36708;
wire g28091, I36711, g28092, I36714, g28093, I36718, g28095, I36721, g28096, I36724, g28097;
wire I36728, g28099, I36738, g28101, I36741, g28102, I36744, g28103, I36749, g28106, I36752;
wire g28107, I36755, g28108, I36758, g28109, I36761, g28110, I36766, g28113, I36769, g28114;
wire I36772, g28115, I36776, g28117, I36786, g28119, I36789, g28120, I36792, g28121, I36797;
wire g28124, I36800, g28125, I36803, g28126, g28128, I36808, g28132, g28133, g28137, g28141;
wire g28149, g28150, g28151, g28152, g28153, g28154, g28155, g28156, g28158, g28159, g28160;
wire g28161, g28162, g28163, g28164, g28165, g28166, g28167, g28168, g28169, g28170, g28172;
wire g28173, g28174, g28175, g28177, g28178, I36848, g28179, g28186, g28187, g28190, I36860;
wire g28194, I36864, g28200, I36867, g28206, I36870, g28207, I36873, g28208, I36876, g28209;
wire I36879, g28210, I36882, g28211, I36885, g28212, I36888, g28213, I36891, g28214, I36894;
wire g28215, I36897, g28216, I36900, g28217, I36903, g28218, I36906, g28219, I36909, g28220;
wire I36912, g28221, I36915, g28222, I36918, g28223, I36921, g28224, I36924, g28225, I36927;
wire g28226, I36930, g28227, I36933, g28228, I36936, g28229, I36939, g28230, I36942, g28231;
wire I36945, g28232, I36948, g28233, I36951, g28234, I36954, g28235, I36957, g28236, I36960;
wire g28237, I36963, g28238, I36966, g28239, I36969, g28240, I36972, g28241, I36975, g28242;
wire I36978, g28243, I36981, g28244, I36984, g28245, I36987, g28246, I36990, g28247, I36993;
wire g28248, I36996, g28249, I36999, g28250, I37002, g28251, I37005, g28252, I37008, g28253;
wire I37011, g28254, I37014, g28255, I37017, g28256, I37020, g28257, I37023, g28258, I37026;
wire g28259, I37029, g28260, I37032, g28261, I37035, g28262, I37038, g28263, I37041, g28264;
wire I37044, g28265, I37047, g28266, I37050, g28267, I37053, g28268, I37056, g28269, I37059;
wire g28270, I37062, g28271, I37065, g28272, I37068, g28273, I37071, g28274, I37074, g28275;
wire I37077, g28276, I37080, g28277, I37083, g28278, I37086, g28279, I37089, g28280, I37092;
wire g28281, I37095, g28282, I37098, g28283, I37101, g28284, I37104, g28285, I37107, g28286;
wire I37110, g28287, I37113, g28288, I37116, g28289, I37119, g28290, I37122, g28291, I37125;
wire g28292, I37128, g28293, I37131, g28294, I37134, g28295, I37137, g28296, I37140, g28297;
wire I37143, g28298, I37146, g28299, I37149, g28300, I37152, g28301, I37155, g28302, I37158;
wire g28303, I37161, g28304, I37164, g28305, I37167, g28306, I37170, g28307, I37173, g28308;
wire I37176, g28309, I37179, g28310, I37182, g28311, I37185, g28312, I37188, g28313, I37191;
wire g28314, I37194, g28315, I37197, g28316, I37200, g28317, I37203, g28318, I37228, g28341;
wire I37232, g28343, I37238, g28347, I37252, g28359, I37260, g28365, I37266, g28369, I37269;
wire g28370, I37273, g28372, I37277, g28374, I37280, g28375, I37284, g28377, I37291, g28382;
wire I37319, g28390, I37330, g28393, I37334, g28395, g28419, I37379, g28432, I37386, g28437;
wire I37394, g28443, I37400, g28447, I37410, g28455, I37415, g28458, I37426, g28467, g28483;
wire g28491, g28496, I37459, g28498, g28500, I37467, g28524, I37471, g28526, I37474, g28527;
wire I37481, g28552, I37484, g28553, g28554, I37488, g28555, I37494, g28579, I37497, g28580;
wire g28581, g28582, I37502, g28583, I37508, g28607, g28608, g28609, g28610, I37514, g28611;
wire g28612, g28616, g28617, g28618, g28619, g28623, g28624, g28625, g28629, g28630, g28638;
wire g28639, g28640, g28641, g28642, g28643, g28644, g28645, g28646, g28647, g28648, g28649;
wire g28650, g28651, g28652, g28653, g28655, I37566, g28673, I37569, g28674, I37572, g28675;
wire I37575, g28676, I37578, g28677, I37581, g28678, I37584, g28679, I37587, g28680, I37590;
wire g28681, I37593, g28682, I37596, g28683, I37599, g28684, I37602, g28685, I37605, g28686;
wire I37608, g28687, I37611, g28688, I37614, g28689, I37617, g28690, I37620, g28691, I37623;
wire g28692, I37626, g28693, I37629, g28694, I37632, g28695, I37635, g28696, I37638, g28697;
wire I37641, g28698, I37644, g28699, I37647, g28700, I37650, g28701, I37653, g28702, I37656;
wire g28703, I37659, g28704, I37662, g28705, I37665, g28706, g28720, g28721, g28723, g28725;
wire g28727, g28730, g28734, g28740, I37702, g28741, I37712, g28751, I37716, g28755, I37725;
wire g28764, I37729, g28768, I37736, g28775, I37740, g28779, I37746, g28785, I37752, g28791;
wire I37757, g28796, I37760, g28799, I37765, g28804, I37768, g28807, I37771, g28810, I37775;
wire g28814, I37778, g28817, I37781, g28820, I37784, g28823, I37787, g28826, I37790, g28829;
wire I37793, g28832, I37796, g28833, I37800, g28835, I37804, g28837, I37808, g28839, g28855;
wire g28859, g28863, g28867, I37842, g28871, I37846, g28877, I37851, g28882, I37854, g28883;
wire I37858, g28889, I37863, g28894, I37868, g28899, I37871, g28900, I37875, g28906, I37880;
wire g28911, I37885, g28916, I37891, g28924, I37894, g28925, I37897, g28928, I37901, g28932;
wire I37906, g28937, I37912, g28945, I37917, g28950, I37920, g28951, I37924, g28955, I37928;
wire g28959, I37934, g28967, I37939, g28972, I37942, g28975, I37946, g28979, I37950, g28983;
wire I37956, g28993, I37961, g28998, I37965, g29002, I37968, g29005, I37973, g29010, I37978;
wire g29019, I37982, g29023, I37986, g29027, I37991, g29032, I37994, g29035, I37999, g29042;
wire I38003, g29046, I38007, g29050, I38011, g29054, I38014, g29057, I38018, g29061, I38024;
wire g29065, I38028, g29069, I38032, g29073, I38035, g29074, I38038, g29075, I38042, g29077;
wire I38046, g29081, I38049, g29082, I38053, g29084, I38056, g29085, I38059, g29086, I38064;
wire g29089, I38068, g29091, I38071, g29092, I38074, g29093, I38077, g29094, I38080, g29095;
wire I38085, g29098, I38088, g29099, I38091, g29100, I38094, g29101, I38097, g29102, I38101;
wire g29104, I38104, g29105, I38107, g29106, I38111, g29108, I38119, g29117, I38122, g29118;
wire I38125, g29119, I38128, g29120, I38136, g29131, I38139, g29132, I38142, g29133, I38145;
wire g29134, I38148, g29135, I38151, g29136, I38154, g29137, I38157, g29138, I38160, g29139;
wire I38163, g29140, I38166, g29141, I38169, g29142, I38172, g29143, I38175, g29144, I38178;
wire g29145, I38181, g29146, I38184, g29147, I38187, g29148, I38190, g29149, I38193, g29150;
wire I38196, g29151, I38199, g29152, I38202, g29153, I38205, g29154, I38208, g29155, I38211;
wire g29156, I38214, g29157, I38217, g29158, I38220, g29159, I38223, g29160, I38226, g29161;
wire I38229, g29162, I38232, g29163, I38235, g29164, I38238, g29165, I38241, g29166, I38245;
wire g29168, I38250, g29171, I38258, g29177, I38272, g29189, I38275, g29190, I38278, g29191;
wire g29192, I38282, g29193, I38321, g29230, I38330, g29237, I38339, g29244, I38342, g29245;
wire I38345, g29246, I38348, g29247, I38352, g29249, I38355, g29250, I38360, g29253, I38363;
wire g29254, I38369, g29258, g29266, I38386, g29267, g29268, g29269, I38391, g29270, g29271;
wire g29272, I38396, g29273, g29274, g29275, I38401, g29276, g29277, I38405, g29278, I38408;
wire g29279, g29280, I38412, g29281, g29282, g29283, g29285, g29286, g29287, I38421, g29288;
wire g29290, g29291, g29292, I38428, g29293, g29295, g29296, I38434, g29297, I38437, g29298;
wire I38440, g29299, g29301, I38447, g29304, I38450, g29305, I38453, g29306, I38456, g29307;
wire I38459, g29308, I38462, g29309, I38466, g29311, I38471, g29314, I38474, g29315, I38477;
wire g29316, I38480, g29317, I38483, g29318, I38486, g29319, I38491, g29322, I38496, g29325;
wire I38499, g29326, I38502, g29327, I38505, g29328, I38510, g29331, I38515, g29334, I38518;
wire g29335, I38524, g29339, I38536, g29349, I38539, g29350, g29356, g29358, I38548, g29359;
wire g29360, g29361, g29362, g29363, g29364, g29365, g29366, g29367, g29368, g29369, g29370;
wire g29371, g29372, g29373, g29374, g29375, g29376, g29377, g29378, g29379, g29380, g29381;
wire g29382, g29383, g29384, g29385, g29386, g29387, g29388, g29389, g29390, g29391, g29392;
wire g29393, g29394, g29395, g29396, g29397, g29398, I38591, g29400, I38594, g29401, g29402;
wire I38599, g29404, I38602, g29405, I38606, g29407, I38609, g29408, I38613, g29410, I38617;
wire g29412, I38620, g29413, I38623, g29414, I38626, g29415, I38629, g29416, I38632, g29417;
wire I38635, g29418, I38638, g29419, I38641, g29420, I38644, g29421, I38647, g29422, I38650;
wire g29423, I38653, g29424, I38656, g29425, I38659, g29426, I38662, g29427, I38665, g29428;
wire I38668, g29429, I38671, g29430, I38674, g29431, I38677, g29432, I38680, g29433, I38683;
wire g29434, I38686, g29435, I38689, g29436, I38692, g29437, I38695, g29438, I38698, g29439;
wire I38701, g29440, I38704, g29441, I38707, g29442, I38710, g29443, I38713, g29444, I38716;
wire g29445, I38719, g29446, I38722, g29447, I38725, g29448, I38728, g29449, I38731, g29450;
wire I38734, g29451, I38737, g29452, I38740, g29453, I38743, g29454, I38746, g29455, I38749;
wire g29456, I38752, g29457, I38755, g29458, I38758, g29459, I38761, g29460, I38764, g29461;
wire I38767, g29462, I38770, g29463, g29491, I38801, g29495, I38804, g29496, I38807, g29497;
wire I38817, g29499, I38827, g29501, I38838, g29504, I38848, g29506, I38851, g29507, I38854;
wire g29508, I38857, g29509, I38860, g29510, I38863, g29511, I38866, g29512, I38869, g29513;
wire I38872, g29514, I38875, g29515, I38878, g29516, I38881, g29517, I38885, g29519, I38898;
wire g29530, I38905, g29535, I38909, g29537, I38916, g29542, I38920, g29544, I38924, g29546;
wire I38931, g29551, I38936, g29554, I38940, g29556, I38947, g29561, I38951, g29563, I38958;
wire g29568, I38975, g29583, I38999, g29627, I39002, g29628, I39005, g29629, I39008, g29630;
wire I39011, g29631, I39014, g29632, I39017, g29633, I39020, g29634, I39023, g29635, I39026;
wire g29636, I39029, g29637, I39032, g29638, I39035, g29639, I39038, g29640, I39041, g29641;
wire I39044, g29642, I39047, g29643, I39050, g29644, I39053, g29645, I39056, g29646, I39059;
wire g29647, I39062, g29648, I39065, g29649, I39068, g29650, I39071, g29651, I39074, g29652;
wire I39077, g29653, I39080, g29654, I39083, g29655, I39086, g29656, I39089, g29657, g29658;
wire g29659, g29660, g29661, g29662, g29664, g29666, g29668, g29673, I39121, g29689, I39124;
wire g29690, I39127, g29691, I39130, g29692, I39133, g29693, I39136, g29694, I39139, g29695;
wire I39142, g29696, I39145, g29697, I39148, g29698, I39151, g29699, I39154, g29700, I39157;
wire g29701, I39160, g29702, I39164, g29704, I39168, g29708, g29716, g29724, g29726, g29739;
wire I39234, g29794, I39237, g29795, I39240, g29796, I39243, g29797, I39246, g29798, I39249;
wire g29799, I39252, g29800, I39255, g29801, I39258, g29802, I39261, g29803, I39264, g29804;
wire I39267, g29805, I39270, g29806, I39273, g29807, I39276, g29808, I39279, g29809, g29823;
wire g29829, g29835, g29840, g29844, g29848, g29849, g29853, g29857, g29861, g29865, g29869;
wire g29873, g29877, g29881, g29885, g29889, g29893, g29897, g29901, g29905, I39398, g29932;
wire I39401, g29933, I39404, g29934, I39407, g29935, I39411, g29937, I39414, g29938, I39418;
wire g29940, I39423, g29943, I39454, g29972, I39457, g29973, I39460, g29974, I39463, g29975;
wire I39466, g29976, I39469, g29977, I39472, g29978, I39475, g29979, g30036, g30040, g30044;
wire g30048, I39550, g30052, I39573, g30076, I39577, g30078, I39585, g30084, I39622, g30119;
wire I39625, g30120, I39628, g30121, I39631, g30122, I39635, g30124, I39638, g30125, I39641;
wire g30126, I39647, g30130, g30134, g30139, g30143, g30147, g30151, g30155, g30159, g30163;
wire g30167, g30171, g30175, g30179, g30183, g30187, g30191, g30195, g30199, g30203, g30207;
wire g30211, I39674, g30215, g30229, g30233, g30237, g30241, I39761, g30306, I39764, g30307;
wire I39767, g30308, I39770, g30309, I39773, g30310, I39776, g30311, I39779, g30312, I39782;
wire g30313, I39785, g30314, I39788, g30315, I39791, g30316, I39794, g30317, I39797, g30318;
wire I39800, g30319, I39803, g30320, I39806, g30321, I39809, g30322, I39812, g30323, I39815;
wire g30324, I39818, g30325, I39821, g30326, I39825, g30328, I39828, g30329, I39832, g30331;
wire I39835, g30332, I39840, g30335, I39843, g30336, I39848, g30339, I39853, g30342, I39856;
wire g30343, I39859, g30344, I39863, g30346, I39866, g30347, I39870, g30349, I39873, g30350;
wire I39878, g30353, I39881, g30354, I39886, g30357, I39889, g30358, I39892, g30359, I39895;
wire g30360, I39899, g30362, I39902, g30363, I39906, g30365, I39909, g30366, I39913, g30368;
wire I39916, g30369, I39919, g30370, I39922, g30371, I39926, g30373, I39930, g30375, I39933;
wire g30376, I39936, g30377, I39939, g30378, I39942, g30379, I39945, g30380, I39948, g30381;
wire I39951, g30382, g30383, I39976, g30408, I39982, g30412, I39985, g30435, I39991, g30439;
wire I39997, g30443, I40002, g30446, I40008, g30450, I40016, g30456, I40021, g30459, I40027;
wire g30463, I40032, g30466, I40039, g30471, I40044, g30474, I40051, g30479, I40054, g30480;
wire I40059, g30483, I40066, g30488, I40071, g30491, I40075, g30493, I40078, g30494, I40083;
wire g30497, I40086, g30498, I40091, g30501, I40098, g30506, I40101, g30507, I40104, g30508;
wire I40107, g30509, I40110, g30510, I40113, g30511, I40116, g30512, I40119, g30513, I40122;
wire g30514, I40125, g30515, I40128, g30516, I40131, g30517, I40134, g30518, I40137, g30519;
wire I40140, g30520, I40143, g30521, I40146, g30522, I40149, g30523, I40152, g30524, I40155;
wire g30525, I40158, g30526, I40161, g30527, I40164, g30528, I40167, g30529, I40170, g30530;
wire I40173, g30531, I40176, g30532, I40179, g30533, I40182, g30534, I40185, g30535, I40188;
wire g30536, I40191, g30537, I40194, g30538, I40197, g30539, I40200, g30540, I40203, g30541;
wire I40206, g30542, I40209, g30543, I40212, g30544, I40215, g30545, I40218, g30546, I40221;
wire g30547, I40224, g30548, I40227, g30549, I40230, g30550, I40233, g30551, I40236, g30552;
wire I40239, g30553, I40242, g30554, I40245, g30555, I40248, g30556, I40251, g30557, I40254;
wire g30558, I40257, g30559, I40260, g30560, I40263, g30561, I40266, g30562, I40269, g30563;
wire I40272, g30564, I40275, g30565, g30567, g30568, g30569, g30570, g30571, g30572, g30573;
wire g30574, g30575, I40288, g30578, I40291, g30579, I40294, g30580, I40297, g30581, I40300;
wire g30582, I40303, g30583, I40307, g30585, I40310, g30586, I40313, g30587, I40317, g30591;
wire I40320, g30592, I40326, g30600, I40420, g30710, I40423, g30711, I40426, g30712, I40429;
wire g30713, I40432, g30714, I40435, g30715, I40438, g30716, I40441, g30717, I40444, g30718;
wire I40447, g30719, I40450, g30720, I40453, g30721, I40456, g30722, I40459, g30723, I40462;
wire g30724, I40465, g30725, I40468, g30726, I40471, g30727, I40475, g30729, I40478, g30730;
wire I40481, g30731, I40484, g30732, I40487, g30733, I40490, g30734, I40495, g30737, I40498;
wire g30738, I40501, g30739, I40504, g30740, I40507, g30741, I40510, g30742, I40515, g30745;
wire I40518, g30746, I40521, g30747, I40524, g30748, I40527, g30749, I40531, g30751, I40534;
wire g30752, I40537, g30753, I40542, g30756, g30765, I40555, g30767, I40565, g30769, I40568;
wire g30770, I40578, g30772, I40581, g30773, I40584, g30774, I40594, g30776, I40597, g30777;
wire I40600, g30778, I40611, g30781, I40614, g30782, I40618, g30784, I40634, g30792, I40637;
wire g30793, I40640, g30794, I40643, g30795, I40647, g30797, I40651, g30799, I40654, g30800;
wire I40658, g30802, I40661, g30803, I40664, g30804, I40667, g30805, I40670, g30806, I40673;
wire g30807, I40676, g30808, I40679, g30809, I40682, g30810, I40685, g30811, I40688, g30812;
wire I40691, g30813, I40694, g30814, I40697, g30815, I40700, g30816, I40703, g30817, I40706;
wire g30818, I40709, g30819, I40712, g30820, I40715, g30821, I40718, g30822, I40721, g30823;
wire I40724, g30824, I40727, g30825, I40730, g30826, I40733, g30827, I40736, g30828, I40739;
wire g30829, I40742, g30830, I40745, g30831, I40748, g30832, I40751, g30833, I40754, g30834;
wire I40757, g30835, I40760, g30836, I40763, g30837, I40766, g30838, I40769, g30839, I40772;
wire g30840, I40775, g30841, I40778, g30842, I40781, g30843, I40784, g30844, I40787, g30845;
wire I40790, g30846, I40793, g30847, I40796, g30848, I40799, g30849, I40802, g30850, I40805;
wire g30851, I40808, g30852, I40811, g30853, I40814, g30854, I40817, g30855, I40820, g30856;
wire I40823, g30857, I40826, g30858, I40829, g30859, I40832, g30860, I40835, g30861, I40838;
wire g30862, I40841, g30863, I40844, g30864, I40847, g30865, I40850, g30866, I40853, g30867;
wire I40856, g30868, I40859, g30869, I40862, g30870, I40865, g30871, I40868, g30872, I40871;
wire g30873, I40874, g30874, I40877, g30875, I40880, g30876, I40883, g30877, I40886, g30878;
wire I40889, g30879, I40892, g30880, I40895, g30881, I40898, g30882, I40901, g30883, I40904;
wire g30884, I40907, g30885, I40910, g30886, I40913, g30887, I40916, g30888, I40919, g30889;
wire I40922, g30890, I40925, g30891, I40928, g30892, I40931, g30893, I40934, g30894, I40937;
wire g30895, I40940, g30896, I40943, g30897, I40946, g30898, I40949, g30899, I40952, g30900;
wire I40955, g30901, I40958, g30902, I40961, g30903, I40964, g30904, I40967, g30905, I40970;
wire g30906, I40973, g30907, I40976, g30908, I40979, g30909, I40982, g30910, I40985, g30911;
wire I40988, g30912, I40991, g30913, I40994, g30914, I40997, g30915, I41024, g30928, I41035;
wire g30937, I41038, g30938, I41041, g30939, I41044, g30940, I41047, g30941, I41050, g30942;
wire I41053, g30943, g30962, g30963, g30964, g30965, g30966, g30967, g30968, g30969, g30971;
wire I41090, g30972, I41093, g30973, I41096, g30974, I41099, g30975, I41102, g30976, I41105;
wire g30977, I41108, g30978, I41111, g30979, I41114, g30980, I41117, g30981, I41120, g30982;
wire I41123, g30983, I41126, g30984, I41129, g30985, I41132, g30986, I41135, g30987, I41138;
wire g30988, I41141, g30989, g5630, g5649, g5650, g5658, g5676, g5677, g5678, g5687;
wire g5688, g5696, g5709, g5710, g5711, g5728, g5729, g5730, g5739, g5740, g5748;
wire g5757, g5758, g5767, g5768, g5769, g5786, g5787, g5788, g5797, g5798, g5807;
wire g5816, g5817, g5826, g5827, g5828, g5845, g5846, g5847, g5863, g5872, g5873;
wire g5882, g5883, g5884, g5910, g5919, g5920, g5949, g8327, g8328, g8329, g8339;
wire g8340, g8350, g8385, g8386, g8387, g8394, g8395, g8396, g8406, g8407, g8417;
wire g8431, g8432, g8433, g8437, g8438, g8439, g8446, g8447, g8448, g8458, g8459;
wire g8463, g8464, g8465, g8466, g8467, g8468, g8472, g8473, g8474, g8481, g8482;
wire g8483, g8484, g8485, g8486, g8487, g8488, g8489, g8490, g8491, g8492, g8493;
wire g8497, g8498, g8499, g8500, g8501, g8502, g8503, g8504, g8505, g8506, g8507;
wire g8508, g8509, g8510, g8511, g8512, g8513, g8515, g8516, g8517, g8518, g8519;
wire g8520, g8521, g8522, g8523, g8524, g8525, g8526, g8527, g8528, g8529, g8531;
wire g8532, g8534, g8535, g8536, g8537, g8538, g8539, g8540, g8541, g8542, g8543;
wire g8544, g8545, g8546, g8548, g8549, g8551, g8552, g8553, g8554, g8555, g8556;
wire g8557, g8558, g8559, g8561, g8562, g8564, g8565, g8566, g8567, g8570, g8572;
wire g8573, g8576, g8601, g8612, g8613, g8621, g8625, g8626, g8631, g8635, g8636;
wire g8650, g8654, g8666, g8676, g8687, g8688, g8703, g8704, g8705, g8706, g8717;
wire g8722, g8723, g8724, g8725, g8751, g8755, g8760, g8761, g8762, g8774, g8778;
wire g8783, g8784, g8797, g8801, g8816, g8841, g8842, g8861, g8868, g8869, g8892;
wire g8899, g8906, g8907, g8932, g8939, g8946, g8947, g8972, g8979, g9004, g9009;
wire g9026, g9033, g9034, g9047, g9048, g9049, g9056, g9057, g9061, g9062, g9063;
wire g9064, g9065, g9066, g9073, g9074, g9075, g9076, g9077, g9078, g9079, g9080;
wire g9081, g9082, g9083, g9090, g9091, g9092, g9093, g9094, g9095, g9096, g9097;
wire g9098, g9099, g9100, g9101, g9102, g9103, g9104, g9105, g9106, g9107, g9108;
wire g9109, g9110, g9111, g9112, g9113, g9114, g9115, g9116, g9117, g9118, g9119;
wire g9120, g9121, g9122, g9123, g9124, g9125, g9126, g9127, g9131, g9132, g9133;
wire g9137, g9138, g9139, g9143, g9145, g9241, g9301, g9302, g9319, g9364, g9365;
wire g9366, g9367, g9382, g9383, g9400, g9438, g9439, g9440, g9441, g9442, g9461;
wire g9462, g9463, g9464, g9479, g9480, g9497, g9518, g9519, g9520, g9521, g9522;
wire g9523, g9534, g9580, g9581, g9582, g9583, g9584, g9603, g9604, g9605, g9606;
wire g9621, g9622, g9630, g9631, g9632, g9633, g9634, g9635, I16735, I16736, g9636;
wire g9639, g9647, g9648, g9660, g9661, g9662, g9663, g9664, g9665, g9676, g9722;
wire g9723, g9724, g9725, g9726, g9745, g9746, g9747, g9748, g9759, g9760, g9761;
wire g9762, g9763, g9764, g9765, g9766, g9773, g9774, g9775, g9776, g9777, g9778;
wire g9779, g9780, g9781, I16826, I16827, g9782, g9785, g9793, g9794, g9806, g9807;
wire g9808, g9809, g9810, g9811, g9822, g9868, g9869, g9870, g9871, g9872, g9887;
wire g9888, g9889, g9890, g9891, g9892, g9893, g9894, g9901, g9902, g9903, g9904;
wire g9905, g9906, g9907, g9908, g9909, g9910, g9911, g9912, g9919, g9920, g9921;
wire g9922, g9923, g9924, g9925, g9926, g9927, I16930, I16931, g9928, g9931, g9939;
wire g9940, g9952, g9953, g9954, g9955, g9956, g9957, g9968, g10007, g10008, g10009;
wire g10010, g10011, g10012, g10013, g10014, g10024, g10035, g10036, g10037, g10041, g10042;
wire g10043, g10044, g10045, g10046, g10047, g10048, g10055, g10056, g10057, g10058, g10059;
wire g10060, g10061, g10062, g10063, g10064, g10065, g10066, g10073, g10074, g10075, g10076;
wire g10077, g10078, g10079, g10080, g10081, I17042, I17043, g10082, g10085, g10093, g10094;
wire g10101, g10102, g10103, g10104, g10105, g10106, g10107, g10108, g10112, g10113, g10114;
wire g10115, g10116, g10117, g10118, g10119, g10120, g10121, g10122, g10123, g10133, g10144;
wire g10145, g10146, g10150, g10151, g10152, g10153, g10154, g10155, g10156, g10157, g10164;
wire g10165, g10166, g10167, g10168, g10169, g10170, g10171, g10172, g10173, g10174, g10175;
wire g10182, g10183, g10184, I17156, g10186, g10192, g10193, g10194, g10195, g10196, g10197;
wire g10198, g10199, g10200, g10201, g10202, g10203, g10204, g10205, g10206, g10207, g10208;
wire g10209, g10210, g10211, g10212, g10213, g10217, g10218, g10219, g10220, g10221, g10222;
wire g10223, g10224, g10225, g10226, g10227, g10228, g10238, g10249, g10250, g10251, g10255;
wire g10256, g10257, g10258, g10259, g10260, g10261, g10262, g10269, g10270, g10271, g10272;
wire g10279, g10280, g10281, g10282, g10283, g10284, g10285, g10286, g10287, g10288, g10289;
wire g10290, g10291, g10292, g10293, g10294, g10295, g10296, g10297, g10298, g10299, g10300;
wire g10301, g10302, g10303, g10304, g10305, g10306, g10307, g10308, g10309, g10310, g10311;
wire g10312, g10313, g10314, g10315, g10319, g10320, g10321, g10322, g10323, g10324, g10325;
wire g10326, g10327, g10328, g10329, g10330, g10340, g10351, g10352, g10353, g10360, g10361;
wire g10362, g10363, g10364, g10365, g10366, g10367, g10368, g10369, g10370, g10371, g10372;
wire g10373, g10374, g10375, g10376, g10377, g10378, g10379, g10380, g10381, g10382, g10383;
wire g10384, g10385, g10386, g10387, g10388, g10389, g10390, g10391, g10392, g10393, g10394;
wire g10395, g10396, g10397, g10398, g10399, g10400, g10401, g10402, g10403, g10404, g10405;
wire g10406, g10407, g10408, g10412, g10413, g10414, g10415, g10422, g10423, g10430, g10431;
wire g10432, g10433, g10434, g10435, g10436, g10437, g10438, g10439, g10440, g10441, g10442;
wire g10443, g10444, g10445, g10446, g10447, g10448, g10449, g10450, g10451, g10452, g10453;
wire g10454, g10455, g10456, g10457, g10458, g10459, g10460, g10461, g10462, g10463, g10464;
wire g10465, g10466, g10467, g10468, g10469, g10470, g10471, g10472, g10473, g10474, g10475;
wire g10476, g10477, g10478, g10479, I17429, g10480, g10485, g10492, g10493, g10494, g10495;
wire g10496, g10497, g10498, g10499, g10506, g10507, g10508, g10509, g10510, g10511, g10512;
wire g10513, g10514, g10515, g10516, g10517, g10518, g10519, g10520, g10521, g10522, g10523;
wire g10524, g10525, g10526, g10527, g10528, g10529, g10530, g10531, g10532, g10533, g10534;
wire g10535, g10536, g10537, g10538, g10539, g10540, g10541, g10548, g10555, g10556, g10557;
wire g10558, g10559, g10566, g10567, g10568, g10569, g10570, g10571, g10572, g10573, g10580;
wire g10581, g10582, g10583, g10584, g10585, g10586, g10587, g10588, g10589, g10590, g10591;
wire g10592, g10593, g10594, g10595, g10596, g10597, g10598, g10599, g10600, g10604, g10605;
wire g10612, g10613, g10614, g10615, g10616, g10623, g10624, g10625, g10626, g10627, g10628;
wire g10629, g10630, g10637, g10638, g10639, g10640, g10641, g10642, g10643, g10644, g10645;
wire g10650, g10651, g10652, g10659, g10660, g10661, g10662, g10663, g10670, g10671, g10672;
wire g10673, g10674, g10675, g10678, g10680, g10681, g10682, g10689, g10690, g10691, g10692;
wire g10693, g10704, g10707, g10709, g10710, I17599, g10711, g10724, g10727, g10729, g10745;
wire g10748, g10764, g11347, g11420, g11421, g11431, g11607, g11612, g11637, g11771, g11788;
wire g11805, g11814, g11816, g11838, g11847, g11851, g11880, g11885, g11922, g11926, g11966;
wire g11967, g12012, g12069, g12070, g12128, g12129, g12186, g12273, g12274, g12307, g12330;
wire g12331, g12353, g12376, g12419, g12429, g12477, g12494, g12514, g12531, g12650, I19937;
wire I19938, g12876, g12908, I19971, I19972, g12916, g12938, I19996, I19997, g12945, g12966;
wire I20021, I20022, g12974, g12989, g12990, g13000, g13004, g13009, g13010, g13023, g13031;
wire g13032, g13042, I20100, g13055, g13056, I20131, I20132, g13082, g13110, g13247, g13266;
wire g13270, g13289, g13291, g13295, g13316, g13320, g13322, g13326, g13335, g13340, g13343;
wire g13345, g13355, g13360, g13365, g13368, g13385, g13390, g13395, g13477, g13479, g13480;
wire g13481, g13483, g13484, g13485, g13486, g13487, g13488, g13489, g13490, g13491, g13492;
wire g13493, g13496, g13498, g13499, g13500, g13502, g13503, g13504, g13505, g13506, g13513;
wire g13515, g13516, g13517, g13527, g13609, g13619, g13623, g13625, g13631, g13634, g13636;
wire g13642, g13643, g13645, g13646, g13648, g13654, g13655, g13656, g13671, g13672, g13674;
wire g13675, g13676, g13701, g13702, g13703, g13704, g13705, g13738, g13739, g13740, g13755;
wire g13787, g13788, g13789, g13790, g13796, g13815, g13816, g13818, g13824, g13833, g13834;
wire g13835, g13837, g13839, g13845, g13846, g13847, g13851, g13853, g13854, g13855, g13860;
wire g13862, g13865, g13870, g13871, g13878, g13880, g13884, g13892, g13900, g13902, g13904;
wire g13905, g13913, g13914, g13933, g13941, g13943, g13944, g13952, g13953, g13969, g13970;
wire g13989, g13997, g13998, g14006, g14007, g14022, g14023, g14039, g14040, g14059, g14067;
wire g14097, g14098, g14113, g14114, g14130, g14131, g14143, g14182, g14212, g14213, g14228;
wire g14229, g14297, g14327, g14328, g14336, g14419, g14690, g14724, g14752, g14767, g14773;
wire g14884, g14894, g14956, g14957, g14958, g14975, g15020, g15030, g15031, g15046, g15047;
wire g15064, g15093, g15094, g15104, g15105, g15126, g15127, g15142, g15143, g15160, g15171;
wire g15172, g15173, g15178, g15196, g15197, g15218, g15219, g15234, g15235, g15243, g15244;
wire g15245, g15246, g15247, g15257, g15258, g15259, g15264, g15282, g15283, g15304, g15305;
wire g15320, g15321, g15324, g15325, g15335, g15336, g15337, g15338, g15339, g15349, g15350;
wire g15351, g15356, g15374, g15375, g15388, g15389, g15391, g15392, g15402, g15403, g15407;
wire g15410, g15411, g15421, g15422, g15423, g15424, g15425, g15435, g15436, g15437, g15442;
wire g15452, g15453, g15459, g15460, g15470, g15475, g15476, g15486, g15487, g15491, g15494;
wire g15495, g15505, g15506, g15507, g15508, g15509, g15519, g15520, g15526, g15527, g15545;
wire g15546, g15556, g15561, g15562, g15572, g15573, g15577, g15580, g15581, g15591, g15592;
wire g15593, g15594, g15595, g15604, g15605, g15623, g15624, g15634, g15639, g15640, g15650;
wire g15651, g15658, g15666, g15670, g15671, g15680, g15681, g15699, g15700, g15710, g15717;
wire g15725, g15729, g15730, g15739, g15740, g15753, g15754, g15755, g15765, g15769, g15770;
wire I22028, g15780, g15781, g15793, g15801, g15802, g15817, g15828, g15829, g15840, g15852;
wire I22136, g15902, g15998, g16003, g16004, g16008, g16009, g16010, g16015, g16016, g16017;
wire g16018, g16019, g16028, g16029, g16030, g16031, g16032, g16033, g16045, g16046, g16047;
wire g16048, g16049, g16050, g16051, g16052, g16053, g16066, g16067, g16068, g16069, g16070;
wire g16071, g16072, g16073, g16074, g16081, g16089, g16100, g16101, g16102, g16103, g16104;
wire g16105, g16106, g16107, g16108, g16109, g16110, g16111, g16112, g16119, g16127, g16133;
wire g16134, g16135, g16136, g16137, g16138, g16139, g16140, g16141, g16152, g16153, g16158;
wire g16159, g16160, g16161, g16162, g16163, g16170, g16178, g16182, g16183, g16184, g16185;
wire g16186, g16187, g16188, g16197, g16198, g16199, g16200, g16211, g16212, g16217, g16218;
wire g16219, g16220, g16221, g16222, g16229, g16237, g16238, g16239, g16240, g16241, g16242;
wire g16250, g16251, g16252, g16253, g16262, g16263, g16264, g16265, g16276, g16277, g16282;
wire g16283, g16284, g16285, g16286, g16288, g16289, g16290, g16291, g16292, g16298, g16299;
wire g16300, g16301, g16309, g16310, g16311, g16312, g16321, g16322, g16323, g16324, g16335;
wire g16336, g16342, g16343, g16344, g16345, g16346, g16347, g16348, g16349, g16350, g16356;
wire g16357, g16358, g16359, g16367, g16368, g16369, g16370, g16379, g16380, g16381, g16382;
wire g16383, g16384, g16385, g16386, g16387, g16388, g16389, g16390, g16391, g16392, g16393;
wire g16394, g16400, g16401, g16402, g16403, g16411, g16413, g16414, g16415, g16416, g16417;
wire g16418, g16419, g16420, g16421, g16422, g16423, g16424, g16425, g16426, g16427, g16428;
wire g16429, g16430, g16431, g16432, g16438, g16443, g16444, g16445, g16447, g16448, g16449;
wire g16450, g16451, g16452, g16453, g16454, g16455, g16456, g16457, g16458, g16459, g16460;
wire g16461, g16462, g16505, g16513, g16527, g16535, g16558, g16590, g16607, g16625, g16639;
wire g16650, g16850, g16855, g16856, g16859, g16864, g16865, g16879, g16894, g16907, g16908;
wire g16909, g16923, g16938, g16939, g16953, g16964, g16966, g16967, g16968, g16969, g16970;
wire g16984, g16987, g16988, g16989, g16990, g16991, g16993, g16994, g16997, g16998, g16999;
wire g17001, g17015, g17017, g17018, g17021, g17022, g17023, g17028, g17031, g17045, g17047;
wire g17048, g17055, g17056, g17062, g17065, g17079, g17081, g17082, g17084, g17090, g17091;
wire g17097, g17100, g17114, g17116, g17117, g17122, g17128, g17129, g17135, g17138, g17143;
wire g17144, g17149, g17155, g17156, g17161, g17166, g17167, g17172, g17176, g17181, g17182;
wire g17193, g17268, g17301, g17339, g17352, g17353, g17381, g17382, g17393, g17395, g17396;
wire g17397, g17398, g17408, g17409, g17428, g17446, g17447, g17448, g17449, g17450, g17460;
wire g17461, g17462, g17463, g17464, g17474, g17475, g17485, g17486, g17506, g17508, g17509;
wire g17510, g17526, g17527, g17528, g17529, g17530, g17540, g17541, g17542, g17543, g17544;
wire g17554, g17555, g17556, g17576, g17577, g17578, g17597, g17598, g17599, g17600, g17616;
wire g17617, g17618, g17619, g17620, g17630, g17631, g17632, g17633, g17634, g17635, g17636;
wire g17652, g17653, g17654, g17673, g17674, g17675, g17694, g17695, g17696, g17697, g17713;
wire g17714, g17715, g17716, g17717, g17718, g17719, g17734, g17735, g17736, g17737, g17752;
wire g17753, g17754, g17773, g17774, g17775, g17794, g17795, g17796, g17797, g17798, g17812;
wire g17813, g17814, g17824, g17835, g17836, g17837, g17838, g17853, g17854, g17855, g17874;
wire g17875, g17876, g17877, g17900, g17901, g17902, g17912, g17924, g17925, g17926, g17936;
wire g17947, g17948, g17949, g17950, g17965, g17966, g17967, g17989, g17990, g18011, g18012;
wire g18013, g18023, g18035, g18036, g18037, g18047, g18058, g18059, g18060, g18061, g18062;
wire g18088, g18106, g18107, g18128, g18129, g18130, g18140, g18152, g18153, g18154, g18164;
wire g18165, g18169, g18204, g18222, g18223, g18244, g18245, g18246, g18256, g18311, g18329;
wire g18330, g18333, g18404, I24619, g18547, I24689, g18597, I24738, g18629, I24758, g18638;
wire g18645, g18647, g18648, g18649, g18650, g18651, g18652, g18653, g18654, g18655, g18665;
wire g18666, g18667, g18668, g18688, g18689, g18690, g18717, g18718, g18753, g18982, g18990;
wire g18994, g18997, g19007, g19010, g19063, g19079, g19080, g19087, g19088, g19089, g19090;
wire g19092, g19093, g19094, g19095, I25280, g19097, g19099, g19100, g19101, g19102, I25291;
wire g19104, g19106, g19107, g19108, I25300, g19109, g19111, g19112, I25311, g19116, g19117;
wire g19124, g19131, g19142, g19143, g19146, g19148, g19150, g19155, g19161, g19166, g19228;
wire g19236, g19241, g19248, g19252, g19254, g19260, g19267, g19282, g19284, g19285, g19289;
wire g19303, g19307, g19316, g19317, g19320, g19324, g19328, g19347, g19351, g19355, g19356;
wire g19381, g19385, g19413, g19449, g19476, g19499, g19520, g19531, g19540, g19541, g19544;
wire g19545, g19547, g19548, g19549, g19551, g19552, g19553, g19554, g19555, g19557, g19558;
wire g19559, g19560, g19561, g19562, g19564, g19565, g19566, g19567, g19568, g19569, g19570;
wire g19571, g19572, g19574, g19575, g19576, g19584, g19585, g19586, g19587, g19588, g19589;
wire g19590, g19591, g19592, g19593, g19594, g19597, g19598, g19599, g19600, g19601, g19602;
wire g19603, g19604, g19605, g19606, g19614, g19615, g19616, g19617, g19618, g19619, g19620;
wire g19621, g19623, g19624, g19625, g19626, g19627, g19628, g19629, g19630, g19631, g19632;
wire g19633, g19634, g19635, g19636, g19637, g19638, g19639, g19647, g19648, g19649, g19650;
wire g19651, g19653, g19654, g19655, g19656, g19660, g19661, g19662, g19663, g19664, g19665;
wire g19666, g19667, g19668, g19669, g19670, g19671, g19672, g19673, g19674, g19675, g19676;
wire g19677, g19678, g19679, g19687, g19688, g19691, g19692, g19693, g19694, g19695, g19697;
wire g19698, g19699, g19700, g19701, g19702, g19703, g19704, g19708, g19709, g19710, g19711;
wire g19712, g19713, g19714, g19715, g19716, g19717, g19718, g19719, g19720, g19721, g19722;
wire g19723, g19724, g19726, g19727, g19728, g19729, g19730, g19731, g19732, g19733, g19734;
wire g19735, g19736, g19737, g19738, g19739, g19741, g19742, g19743, g19744, g19745, g19746;
wire g19747, g19748, g19752, g19753, g19754, g19755, g19756, g19757, g19758, g19759, g19760;
wire g19761, g19764, g19765, g19766, g19767, g19768, g19769, g19770, g19771, g19772, g19773;
wire g19774, g19775, g19776, g19777, g19778, g19779, g19780, g19781, g19782, g19784, g19785;
wire g19786, g19787, g19788, g19789, g19790, g19791, g19795, g19796, g19797, I26240, g19799;
wire g19802, g19803, g19804, g19805, g19806, g19807, g19808, g19809, g19810, g19811, g19812;
wire g19813, g19814, g19815, g19816, g19817, g19818, g19819, g19820, g19821, g19822, g19823;
wire g19824, g19826, g19827, g19828, g19829, g19836, g19837, g19839, g19840, g19841, I26282;
wire g19842, I26285, g19843, g19846, g19847, g19848, g19849, g19850, g19851, g19852, g19853;
wire g19854, g19855, g19856, g19857, g19858, g19859, g19860, g19861, g19862, g19863, g19864;
wire g19868, g19869, g19870, I26311, g19871, g19872, g19873, g19874, I26317, g19875, I26320;
wire g19876, g19879, g19880, g19881, g19882, g19883, g19884, g19885, g19886, g19887, g19888;
wire g19889, g19895, g19899, g19900, g19901, I26348, g19902, g19903, g19904, g19905, I26354;
wire g19906, I26357, g19907, g19910, g19911, g19912, g19913, g19914, g19920, g19924, g19925;
wire g19926, I26377, g19927, g19928, g19929, g19930, I26383, g19931, g19932, g19935, g19939;
wire g19940, g19941, I26396, g19942, g19943, g19944, g19949, g19952, g19953, I26416, g19970;
wire g19971, g19976, I26432, g19982, g19983, I26440, g20000, g20001, g20006, g20011, g20012;
wire g20013, g20014, I26464, g20020, g20021, I26472, g20038, g20039, g20044, g20048, g20049;
wire g20050, g20051, g20052, g20053, I26500, g20062, g20063, I26508, g20080, g20081, g20084;
wire g20085, g20086, g20087, g20088, g20089, g20090, g20091, g20092, I26525, g20093, I26528;
wire g20094, I26541, g20103, g20104, g20106, g20107, g20108, g20109, g20110, g20111, g20112;
wire g20113, g20114, g20115, I26558, g20116, I26561, g20117, I26564, g20118, I26567, g20119;
wire g20131, g20132, g20133, g20134, g20135, g20136, g20137, g20138, g20139, g20144, g20145;
wire I26590, g20146, I26593, g20147, I26596, g20148, I26599, g20149, g20156, g20157, g20158;
wire g20159, g20160, g20161, g20162, I26615, g20177, g20182, g20183, I26621, g20184, I26624;
wire g20185, I26627, g20186, I26630, g20187, g20188, g20189, g20190, g20191, g20192, I26639;
wire g20197, I26645, g20211, g20216, g20217, I26651, g20218, I26654, g20219, g20220, g20221;
wire g20222, I26661, g20227, I26667, g20241, g20246, g20247, g20248, g20249, I26676, g20254;
wire I26682, g20268, g20270, g20271, g20272, I26690, g20277, I26695, g20280, g20282, g20283;
wire g20284, g20285, I26708, g20291, g20293, g20294, I26726, g20307, g20309, I26745, g20326;
wire g20460, g20472, g20480, g20486, g20492, g20499, g20502, g20503, g20506, g20512, g20525;
wire g20538, g20640, g20647, g20665, g20809, g20826, g20836, g20840, g21049, g21067, g21068;
wire g21077, g21078, g21085, g21086, g21091, g21092, g21097, g21098, g21103, g21107, g21111;
wire g21112, g21121, g21122, g21123, g21124, g21128, g21129, I27695, g21136, g21137, g21138;
wire g21140, g21141, g21142, g21143, I27711, g21152, g21153, g21154, g21155, I27717, g21156;
wire g21157, g21158, g21160, g21161, g21162, g21163, I27733, g21172, g21173, g21174, g21175;
wire I27739, g21176, g21177, g21178, g21180, g21181, g21182, g21188, I27755, g21192, g21193;
wire g21194, g21195, I27761, g21196, g21197, g21198, g21203, I27772, g21207, g21208, g21209;
wire g21210, g21218, g21226, g21229, g21234, g21243, g21245, g21251, g21252, g21254, g21259;
wire g21260, g21262, g21267, g21268, g21270, g21276, g21277, g21283, g21284, g21290, g21291;
wire g21292, g21298, g21299, g21300, g21301, g21302, g21303, g21304, g21305, g21306, g21307;
wire g21308, g21309, g21310, g21311, g21312, g21313, g21314, g21315, g21319, g21320, g21321;
wire g21322, g21323, g21324, g21325, g21326, g21328, g21329, g21330, g21334, g21335, g21336;
wire g21337, g21338, g21339, g21340, g21341, g21342, g21343, g21344, g21345, g21349, g21350;
wire g21351, g21352, g21353, g21354, g21355, g21356, g21357, g21360, g21361, g21362, g21363;
wire g21367, g21368, g21369, g21370, g21371, g21372, g21373, g21374, g21375, g21378, g21379;
wire g21380, g21381, g21388, g21389, g21390, g21391, g21392, g21393, g21394, g21395, g21396;
wire g21397, g21398, g21401, g21402, g21403, g21410, g21411, g21412, g21413, g21414, g21418;
wire g21419, g21420, g21421, g21422, g21423, g21424, g21425, g21428, g21438, g21439, g21440;
wire g21444, g21445, g21446, g21447, g21448, g21452, g21453, g21454, g21455, g21456, g21476;
wire g21480, g21481, g21482, g21486, g21487, g21488, g21489, g21490, g21494, g21497, g21517;
wire g21521, g21522, g21523, g21527, I28068, g21533, g21553, I28096, g21564, I28103, g21569;
wire g21589, g21593, I28126, g21597, I28133, g21602, g21610, g21611, g21622, I28155, g21626;
wire I28162, g21631, g21635, g21639, g21650, I28181, g21654, g21658, g21666, g21670, g21681;
wire g21687, g21695, g21699, g21707, g21723, g21731, g21735, g21749, g21757, g21758, g21773;
wire g21805, g21812, g21818, g21822, g21891, g21892, g21899, g21900, g21906, g21911, g21912;
wire g21913, g21920, g21925, g21926, g21931, g21938, g21990, g22004, g22015, g22020, I28582;
wire g22036, I28594, g22046, I28609, g22062, g22187, g22196, g22201, g22202, g22206, g22207;
wire g22208, g22211, g22214, g22215, g22220, g22223, g22224, g22228, g22229, g22235, g22238;
wire g22244, g22245, g22250, g22254, g22255, g22264, g22265, g22270, g22272, g22273, g22281;
wire g22282, g22285, g22289, g22291, g22292, g22305, g22309, g22311, g22312, g22333, g22337;
wire g22340, g22358, g22363, g22383, g22398, g22483, g22515, g22516, g22517, g22526, g22546;
wire g22555, g22556, g22557, g22566, g22577, g22581, g22587, g22595, g22596, g22597, g22606;
wire g22607, g22610, g22614, g22618, g22624, g22632, g22633, g22634, g22637, g22638, g22643;
wire g22646, g22650, g22654, g22660, g22665, g22666, g22667, g22674, g22679, g22682, g22686;
wire g22690, g22699, g22700, g22701, g22707, g22714, g22719, g22722, g22726, g22727, g22732;
wire g22738, g22745, g22754, g22759, g22764, g22770, g22788, g22793, g22798, g22804, g22830;
wire g22835, g22841, g22842, g22869, g22874, g22906, g22984, g23104, g23106, g23118, g23119;
wire g23127, g23128, g23138, g23139, g23409, g23414, g23419, g23423, g23428, g23432, g23434;
wire g23440, g23451, g23458, g23462, g23467, g23471, g23476, g23483, g23484, g23494, g23496;
wire g23510, g23512, g23525, g23527, g23536, g23538, g23544, g23547, g23550, g23551, g23552;
wire g23554, g23558, g23559, g23560, g23563, g23564, g23565, g23567, g23571, g23572, g23573;
wire g23577, g23578, g23579, g23582, g23583, g23584, g23586, g23590, g23591, g23592, g23593;
wire g23598, g23599, g23600, g23604, g23605, g23606, g23609, g23610, g23611, g23615, g23616;
wire g23617, g23618, g23622, g23623, g23624, g23625, g23630, g23631, g23632, g23636, g23637;
wire g23638, g23639, g23643, g23659, g23664, g23665, g23666, g23667, g23671, g23672, g23673;
wire g23674, g23679, g23680, g23681, g23686, g23687, g23689, g23693, g23709, g23714, g23715;
wire g23716, g23717, g23721, g23722, g23723, g23724, g23726, g23734, g23735, g23740, g23741;
wire g23743, g23747, g23763, g23768, g23769, g23770, g23771, g23772, g23776, g23777, g23778;
wire g23789, g23790, g23795, g23796, g23798, g23802, g23818, g23820, g23822, g23824, g23825;
wire g23829, g23830, g23831, g23842, g23843, g23848, g23849, g23851, g23852, g23854, g23855;
wire g23857, g23859, g23860, g23864, g23865, g23866, g23877, g23878, g23886, g23888, g23889;
wire g23891, g23893, g23894, g23898, g23899, g23900, g23904, g23907, g23909, g23910, g23912;
wire g23914, g23915, g23917, g23939, g23941, g23942, g23944, g23971, g23972, g24029, g24211;
wire g24217, g24221, g24224, g24229, g24236, g24241, g24246, g24247, g24253, g24256, g24427;
wire g24429, g24431, g24432, g24433, g24435, g24436, g24437, g24439, g24440, g24441, g24478;
wire g24529, g24540, g24541, g24542, g24550, g24552, g24553, g24554, g24559, g24561, g24563;
wire g24564, g24565, g24569, g24571, g24573, g24574, g24578, g24580, g24585, g24590, g24591;
wire g24595, g24596, g24603, g24604, g24610, g24611, g24644, g24664, g24676, g24683, g24695;
wire g24700, g24712, g24723, g24745, g24746, g24747, g24748, g24749, g24750, g24751, g24752;
wire g24754, g24755, g24757, g24758, g24759, g24760, g24761, g24762, g24767, g24768, g24769;
wire g24772, g24773, g24774, g24775, g24776, g24777, g24779, g24780, g24781, g24788, g24789;
wire g24790, g24792, g24793, g24794, g24795, g24796, g24798, g24799, g24802, g24803, g24804;
wire g24809, g24810, g24811, g24813, g24818, g24821, g24822, g24824, g24825, g24826, g24831;
wire g24838, g24840, g24841, g24843, g24846, g24853, g24855, g24858, g24861, g24867, g24869;
wire g24870, g24874, g24876, g24878, g24881, g24882, g24884, g24885, g24888, g24898, g24899;
wire g24901, g24902, g24905, g24906, g24907, g24908, g24921, g24922, g24924, g24938, g24964;
wire g24974, g25086, g25102, g25117, g25128, g25178, g25181, g25182, g25184, g25187, g25188;
wire g25192, g25193, g25196, g25198, g25269, g25277, g25278, g25281, g25282, g25286, g25287;
wire g25289, g25290, g25294, g25295, g25299, g25300, g25304, g25309, g25310, g25318, g25321;
wire g25328, g25334, g25337, g25342, g25346, g25348, g25351, g25356, g25360, g25362, g25365;
wire g25371, g25375, g25377, g25388, g25392, g25453, g25457, g25461, g25466, g25470, g25475;
wire g25482, g25483, g25487, g25505, g25506, g25513, g25514, g25518, g25552, g25553, g25560;
wire g25561, g25565, g25618, g25619, g25626, g25627, g25628, g25629, g25697, g25881, g25951;
wire g25953, g25957, g25961, g25963, g25968, g25972, g25973, g25975, g25977, g25978, g25980;
wire g25981, g26023, g26024, g26026, g26027, g26028, g26029, g26030, g26032, g26033, g26034;
wire g26035, g26036, g26038, g26039, g26040, g26051, g26052, g26053, g26054, g26060, g26061;
wire g26062, g26067, g26068, g26069, g26074, g26075, g26080, g26082, g26085, g26091, g26157;
wire g26158, g26163, g26166, g26171, g26186, g26188, g26207, g26212, g26213, g26231, g26233;
wire g26234, g26235, g26236, g26243, g26244, g26257, g26258, g26259, g26260, g26261, g26262;
wire g26263, g26268, g26269, g26270, g26271, g26278, g26279, g26288, g26289, g26290, g26291;
wire g26292, g26293, g26298, g26299, g26300, g26301, g26302, g26303, g26307, g26309, g26310;
wire g26311, g26312, g26316, g26317, g26318, g26319, g26324, g26325, g26326, g26332, g26333;
wire g26334, g26335, g26339, g26340, g26342, g26343, g26344, g26345, g26346, g26347, g26348;
wire g26350, g26351, g26352, g26353, g26357, g26361, g26362, g26363, g26365, g26366, g26371;
wire g26372, g26373, g26379, g26380, g26381, g26382, g26383, g26384, g26386, g26387, g26388;
wire g26389, g26390, g26391, g26392, g26396, g26397, g26400, g26404, g26405, g26406, g26408;
wire g26409, g26414, g26415, g26416, g26422, g26423, g26424, g26425, g26426, g26427, g26432;
wire g26437, g26438, g26441, g26445, g26446, g26447, g26449, g26450, g26455, g26456, g26457;
wire g26464, g26469, g26470, g26473, g26477, g26478, g26479, g26488, g26493, g26494, g26504;
wire g26663, g26668, g26673, g26674, g26754, g26755, g26756, g26758, g26759, g26760, g26761;
wire g26763, g26764, g26765, g26766, g26767, g26768, g26769, g26770, g26771, g26773, g26774;
wire g26775, g26777, g26778, g26780, g26783, g26784, g26787, g26790, g26791, g26794, g26797;
wire g26829, g26833, g26842, g26845, g26851, g26853, g26860, g26866, g26955, g26958, g26961;
wire g26962, g26963, g26965, g26966, g26967, g26968, g26969, g26970, g26971, g26972, g26973;
wire g26977, g26978, g26979, g26980, g26981, g26982, g26984, g26985, g26986, g26993, g26994;
wire g26995, g26996, g26997, g26998, g26999, g27000, g27001, g27002, g27003, g27004, g27005;
wire g27006, g27007, g27008, g27009, g27016, g27017, g27018, g27019, g27020, g27021, g27022;
wire g27023, g27024, g27025, g27026, g27027, g27028, g27029, g27030, g27031, g27032, g27033;
wire g27034, g27035, g27042, g27043, g27044, g27045, g27046, g27047, g27048, g27049, g27050;
wire g27052, g27053, g27054, g27055, g27056, g27057, g27058, g27059, g27060, g27061, g27062;
wire g27063, g27070, g27071, g27072, g27073, g27074, g27076, g27077, g27079, g27080, g27081;
wire g27082, g27083, g27084, g27085, g27086, g27087, g27088, g27089, g27090, g27091, g27092;
wire g27093, g27095, g27096, g27097, g27098, g27099, g27100, g27101, g27103, g27104, g27105;
wire g27107, g27108, g27109, g27110, g27111, g27112, g27115, g27178, g27181, g27182, g27185;
wire g27187, g27240, g27241, g27242, g27244, g27245, g27246, g27247, g27248, g27249, g27355;
wire g27356, g27358, g27359, g27364, g27365, g27370, g27371, g27372, g27394, g27396, g27407;
wire g27409, g27425, g27427, g27446, g27448, g27495, g27509, g27516, g27530, g27534, g27541;
wire g27552, g27554, g27561, g27568, g27570, g27578, g27656, g27657, g27659, g27660, g27661;
wire g27666, g27671, g27673, g27679, g27680, g27681, g27719, g27720, g27721, g27723, g27725;
wire g27726, g27727, g27728, g27729, g27730, g27731, g27732, g27733, g27734, g27737, g27770;
wire g27772, g27773, g27774, g27775, g27779, g27783, g27790, g27904, g27908, g27909, g27913;
wire g27914, g27915, g27922, g27923, g27924, g27926, g27931, g27935, g27936, g27938, g27945;
wire g27949, g27951, g27963, g27968, g27970, g27984, g27985, g27991, g28008, g28009, g28015;
wire g28027, g28028, g28035, g28036, g28042, g28050, g28051, g28057, g28058, g28065, g28066;
wire g28073, g28079, g28080, g28086, g28087, g28094, g28098, g28104, g28105, g28111, g28112;
wire g28116, g28122, g28123, g28127, g28171, g28176, g28188, g28193, g28319, g28320, g28322;
wire g28323, g28324, g28326, g28327, g28329, g28330, g28331, g28332, g28333, g28334, g28335;
wire g28336, g28337, g28338, g28339, g28340, g28373, g28376, g28378, g28379, g28380, g28381;
wire g28383, g28385, g28387, g28389, g28396, g28398, g28399, g28401, g28402, g28404, g28405;
wire g28407, g28408, g28411, g28412, g28416, g28422, g28423, g28424, g28426, g28427, g28428;
wire g28429, g28430, g28431, g28433, g28434, g28435, g28436, g28438, g28439, g28440, g28441;
wire g28442, g28444, g28445, g28446, g28448, g28450, g28451, g28452, g28453, g28454, g28456;
wire g28457, g28459, g28460, g28462, g28463, g28464, g28465, g28466, g28468, g28469, g28471;
wire g28472, g28474, g28475, g28476, g28477, g28478, g28479, g28480, g28481, g28484, g28485;
wire g28486, g28487, g28492, g28493, g28494, g28497, g28657, g28659, g28660, g28662, g28663;
wire g28664, g28665, g28666, g28667, g28669, g28670, g28671, g28672, g28707, g28708, g28709;
wire g28710, g28711, g28712, g28713, g28714, g28715, g28716, g28717, g28718, g28719, g28722;
wire g28724, g28726, g28729, g28834, g28836, g28838, g28840, g28841, g28843, g28844, g28846;
wire g28847, g28848, g28849, g28850, g28851, g28852, g28853, g28854, g28880, g28881, g28892;
wire g28893, g28897, g28898, g28909, g28910, g28914, g28915, g28919, g28923, g28931, g28935;
wire g28936, g28940, g28944, g28948, g28949, g28958, g28962, g28966, g28970, g28971, g28986;
wire g28996, g28997, g29022, g29130, g29174, g29175, g29176, g29180, g29183, g29186, g29188;
wire g29196, g29200, g29203, g29208, g29211, g29217, g29220, g29225, g29229, g29232, g29233;
wire g29234, g29235, g29236, g29238, g29239, g29240, g29241, g29242, g29243, g29248, g29251;
wire g29252, g29255, g29256, g29257, g29259, g29260, g29261, g29262, g29263, g29264, g29284;
wire g29289, g29294, g29300, g29302, g29310, g29312, g29320, g29321, g29323, g29329, g29330;
wire g29332, g29336, g29337, g29338, g29341, g29342, g29344, g29346, g29411, g29464, g29465;
wire g29466, g29467, g29468, g29469, g29470, g29471, g29472, g29473, g29474, g29475, g29476;
wire g29477, g29478, g29479, g29480, g29481, g29482, g29483, g29484, g29485, g29486, g29487;
wire g29488, g29489, g29490, g29502, g29518, g29520, g29521, g29522, g29523, g29524, g29525;
wire g29526, g29527, g29528, g29529, g29531, g29532, g29533, g29534, g29536, g29538, g29539;
wire g29540, g29541, g29543, g29545, g29547, g29548, g29549, g29550, g29553, g29555, g29557;
wire g29558, g29559, g29560, g29562, g29564, g29565, g29566, g29567, g29572, g29573, g29575;
wire g29607, g29610, g29614, g29615, g29619, g29622, g29624, g29625, g29626, g29790, g29792;
wire g29793, g29810, g29811, g29812, g29813, g29814, g29815, g29816, g29817, g29818, g29819;
wire g29820, g29821, g29822, g29827, g29828, g29833, g29834, g29839, g29909, g29910, g29942;
wire g29944, g29945, g29946, g29947, g29948, g29949, g29950, g29951, g29952, g29953, g29954;
wire g29955, g29956, g29957, g29958, g29959, g29960, g29961, g29962, g29963, g29964, g29965;
wire g29966, g29967, g29968, g29969, g29970, g29971, g29980, g29981, g29982, g29983, g29984;
wire g29985, g29986, g29987, g29988, g29989, g29990, g29991, g29992, g29993, g29994, g29995;
wire g29996, g29997, g29998, g29999, g30000, g30001, g30002, g30003, g30004, g30005, g30006;
wire g30007, g30008, g30009, g30077, g30079, g30080, g30081, g30082, g30083, g30085, g30086;
wire g30087, g30088, g30089, g30090, g30091, g30092, g30093, g30094, g30095, g30096, g30097;
wire g30098, g30099, g30100, g30101, g30102, g30103, g30104, g30105, g30106, g30107, g30108;
wire g30109, g30110, g30111, g30112, g30113, g30114, g30115, g30116, g30117, g30118, g30123;
wire g30127, g30128, g30129, g30131, g30132, g30133, g30138, g30216, g30217, g30218, g30219;
wire g30220, g30221, g30222, g30223, g30224, g30225, g30226, g30227, g30327, g30330, g30333;
wire g30334, g30337, g30340, g30345, g30348, g30351, g30352, g30355, g30361, g30364, g30367;
wire g30372, g30374, g30387, g30388, g30389, g30390, g30391, g30392, g30393, g30394, g30395;
wire g30396, g30397, g30398, g30407, g30409, g30410, g30411, g30436, g30437, g30438, g30440;
wire g30441, g30442, g30444, g30445, g30447, g30448, g30449, g30451, g30452, g30453, g30454;
wire g30457, g30458, g30460, g30461, g30462, g30464, g30465, g30467, g30469, g30472, g30473;
wire g30475, g30476, g30477, g30478, g30481, g30484, g30486, g30489, g30490, g30492, g30495;
wire g30496, g30499, g30502, g30504, g30696, g30697, g30698, g30728, g30735, g30736, g30743;
wire g30744, g30750, g30754, g30755, g30757, g30758, g30759, g30760, g30761, g30762, g30763;
wire g30764, g30766, g30916, g30917, g30918, g30919, g30920, g30921, g30922, g30923, g30924;
wire g30925, g30944, g30945, g30946, g30947, g30948, g30949, g30950, g30951, g30953, g9144;
wire g10778, g12377, g12407, g12886, g12926, g12955, g12984, g16539, g16571, g16595, g16615;
wire g17973, g19181, g19186, g19187, g19188, g19191, g19192, g19193, g19194, g19195, g19200;
wire g19201, g19202, g19203, g19204, g19205, g19206, g19209, g19210, g19211, g19212, g19213;
wire g19214, g19215, g19216, g19221, g19222, g19223, g19224, g19225, g19226, g19227, I25477;
wire g19230, g19231, g19232, g19233, g19234, g19235, I25495, g19240, g19242, I25500, g19243;
wire g19244, g19245, g19246, g19250, I25516, g19253, g19255, I25521, g19256, g19257, g19263;
wire g19264, I25549, g19266, g19268, I25554, g19269, g19275, g19278, g19279, I25588, g19281;
wire g19283, g19294, g19297, g19298, g19312, g19315, g19333, g19450, g19477, g19500, g19503;
wire g19521, g19522, g19532, g19542, I26429, g19981, I26455, g20015, I26461, g20019, I26491;
wire g20057, I26497, g20061, I26532, g20098, I26538, g20102, I26571, g20123, g21120, g21139;
wire g21159, g21179, g21244, g21253, g21261, g21269, g21501, g21536, g21540, g21572, g21576;
wire g21605, g21609, g21634, g21774, g21787, I28305, g21788, g21789, I28318, g21799, g21800;
wire g21801, I28323, g21802, g21803, g21806, I28330, g21807, g21808, g21809, I28335, g21810;
wire g21811, g21813, I28341, g21814, g21815, g21816, I28346, g21817, g21819, I28351, g21820;
wire g21821, g21823, I28365, g21844, I28369, g21846, I28374, g21849, I28380, g21856, g22175;
wire g22190, g22199, g22205, g22811, g23052, g23071, g23084, g23089, g23100, g23107, g23120;
wire g23129, g23319, g23688, g23742, g23797, g23850, g23919, g24239, g24244, g24245, g24252;
wire g24254, g24257, g24258, g24633, g24653, g24672, g24691, g24890, g24909, g24925, g24965;
wire g24978, g24989, g25000, g25183, g25186, g25190, g25195, g25489, g25490, g25520, g25566;
wire g26320, g26367, g26410, g26451, g26974, g27113, g28501, g28512, g28529, g28540, g28556;
wire g28567, g28584, g28595, g29348, g30305, I15167, I15168, I15169, g7855, I15183, I15184;
wire I15185, g7875, I15190, I15191, I15192, g7876, I15204, I15205, I15206, g7895, I15211;
wire I15212, I15213, g7896, I15237, I15238, I15239, g7922, I15244, I15245, I15246, g7923;
wire I15276, I15277, I15278, g7970, g8381, g8533, g8547, g8550, g8560, g8563, g8571;
wire g8574, g8577, I16879, I16880, I16881, g9883, I16965, I16966, I16967, g10003, g10038;
wire I17059, I17060, I17061, g10095, g10147, I17149, I17150, I17151, g10185, g10252, g10354;
wire g10649, g10676, g10677, g10679, g10703, g10705, g10706, g10708, g10723, g10725, g10726;
wire g10728, g10744, g10746, g10747, g10763, I18106, I18107, I18108, g11188, I18113, I18114;
wire I18115, g11189, I18190, I18191, I18192, g11262, I18197, I18198, I18199, g11263, I18204;
wire I18205, I18206, g11264, I18280, I18281, I18282, g11330, I18287, I18288, I18289, g11331;
wire I18368, I18369, I18370, g11410, g11617, I18799, I18800, I18801, g11621, g11661, g11662;
wire g11672, g11673, g11674, g11683, g11684, g11685, g11686, g11691, g11692, g11693, g11694;
wire g11695, g11696, g11698, g11699, g11700, g11701, g11702, g11704, g11705, g11707, g11708;
wire g11709, g11710, g11712, g11713, g11716, g11717, g11718, g11719, g11720, g11721, g11722;
wire g11723, g11724, g11725, g11726, g11727, g11728, g11729, g11730, g11731, g11733, g12433;
wire g12486, g12503, g12506, g12520, g12523, g12535, g12538, g12544, I20031, I20032, I20033;
wire g12988, I20048, I20049, I20050, g12999, g13020, g13021, g13026, g13027, g13028, g13029;
wire g13030, g13034, g13035, g13037, g13038, g13039, g13040, g13041, g13044, g13045, g13047;
wire g13048, g13050, g13051, g13052, g13053, g13054, g13058, g13059, g13061, g13062, g13064;
wire g13065, g13067, g13068, g13069, g13071, g13072, g13074, g13075, g13077, g13078, g13080;
wire g13081, g13087, g13088, g13089, g13090, g13091, g13093, g13094, g13096, g13097, g13098;
wire g13099, g13100, g13102, g13103, g13104, g13105, g13106, g13108, g13109, g13112, g13113;
wire g13114, g13115, g13116, g13118, g13119, g13120, g13121, g13122, g13123, g13125, g13126;
wire g13127, g13128, g13129, g13131, g13132, g13133, g13134, g13136, g13137, g13138, g13139;
wire g13140, g13142, g13144, g13145, g13146, g13147, g13150, g13156, g13165, g13245, g13305;
wire I20429, I20430, I20431, g13348, I20465, I20466, I20467, g13370, I20504, I20505, I20506;
wire g13399, g13476, g13478, g13482, g13494, g13495, g13497, g13501, I20743, I20744, I20745;
wire g13507, g13510, g13511, g13512, g13514, g13518, g13524, g13525, g13526, g13528, g13529;
wire g13535, g13536, g13537, g13538, g13539, g13540, g13546, g13547, g13548, g13549, g13550;
wire g13551, g13557, g13558, g13559, g13560, g13561, g13562, g13563, g13564, g13599, g13611;
wire g13621, g13633, g13893, g13915, g13934, g13957, g13971, g13990, g14027, g14041, g14060;
wire g14118, g14132, g14233, g15454, g15540, g15618, g15660, g15664, g15694, g15718, g15719;
wire g15720, g15721, g15723, g15756, g15757, g15758, g15759, g15760, g15761, g15763, g15782;
wire g15783, g15784, g15785, g15786, g15787, g15788, g15789, g15791, g15803, g15804, g15805;
wire g15806, g15807, g15808, g15809, g15810, g15811, g15812, I22062, I22063, I22064, g15814;
wire g15818, g15819, g15820, g15821, g15822, g15823, g15824, g15825, g15826, g15827, g15830;
wire g15831, g15832, g15833, g15834, g15835, g15836, g15837, g15838, g15839, g15841, g15842;
wire g15843, g15844, g15845, g15846, g15847, g15848, g15849, g15850, g15851, g15853, g15854;
wire g15855, g15856, g15857, g15858, g15866, g15867, g15868, g15869, g15870, g15871, g15872;
wire g15877, g15878, g15879, g15887, g15888, g15889, g15897, g15898, g15899, g15900, g15901;
wire g15903, g15912, g15920, g15921, g15922, g15930, g15931, g15932, g15941, g15949, g15950;
wire g15951, g15970, g15990, g15992, g15993, g15995, g15996, g15999, g16000, g16006, g16085;
wire g16123, I22282, I22283, I22284, g16132, g16174, I22316, I22317, I22318, g16181, g16233;
wire g16341, g16412, g16439, g16442, g16446, g16463, g16536, I22630, I22631, I22632, g16566;
wire I22705, I22706, I22707, g16662, I22884, I22885, I22886, g16935, I22900, I22901, I22902;
wire g16965, I22917, I22918, I22919, g16985, I22924, I22925, I22926, g16986, I22936, I22937;
wire I22938, g16992, I22945, I22946, I22947, g16995, I22952, I22953, I22954, g16996, I22962;
wire I22963, I22964, g17000, I22972, I22973, I22974, g17016, I22981, I22982, I22983, g17019;
wire I22988, I22989, I22990, g17020, I22998, I22999, I23000, g17024, I23008, I23009, I23010;
wire g17030, I23018, I23019, I23020, g17046, I23027, I23028, I23029, g17049, I23034, I23035;
wire I23036, g17050, I23045, I23046, I23047, g17058, I23055, I23056, I23057, g17064, I23065;
wire I23066, I23067, g17080, I23074, I23075, I23076, g17083, I23082, I23083, I23084, g17085;
wire I23093, I23094, I23095, g17093, I23103, I23104, I23105, g17099, I23113, I23114, I23115;
wire g17115, g17118, I23123, I23124, I23125, g17121, I23131, I23132, I23133, g17123, I23142;
wire I23143, I23144, g17131, I23152, I23153, I23154, g17137, g17139, I23161, I23162, I23163;
wire g17142, g17145, I23171, I23172, I23173, g17148, I23179, I23180, I23181, g17150, I23190;
wire I23191, I23192, g17158, g17159, I23198, I23199, I23200, g17160, g17162, I23207, I23208;
wire I23209, g17165, g17168, I23217, I23218, I23219, g17171, I23225, I23226, I23227, g17173;
wire g17174, I23233, I23234, I23235, g17175, g17177, I23242, I23243, I23244, g17180, g17183;
wire I23256, I23257, I23258, g17190, g17191, I23264, I23265, I23266, g17192, g17194, I23277;
wire I23278, I23279, g17201, g17202, I23806, I23807, I23808, g17729, I23878, I23879, I23880;
wire g17807, I23893, I23894, I23895, g17830, I23941, I23942, I23943, g17887, I23958, I23959;
wire I23960, g17913, I23966, I23967, I23968, g17919, I23981, I23982, I23983, g17942, I24005;
wire I24006, I24007, g17968, I24015, I24016, I24017, g17979, g17985, I24028, I24029, I24030;
wire g17992, I24036, I24037, I24038, g17998, I24053, I24054, I24055, g18024, I24061, I24062;
wire I24063, g18030, I24076, I24077, I24078, g18053, I24091, I24092, I24093, g18079, I24102;
wire I24103, I24104, g18090, I24110, I24111, I24112, g18096, g18102, I24123, I24124, I24125;
wire g18109, I24131, I24132, I24133, g18115, I24148, I24149, I24150, g18141, I24156, I24157;
wire I24158, g18147, I24178, I24179, I24180, g18183, I24186, I24187, I24188, g18189, I24194;
wire I24195, I24196, g18195, I24205, I24206, I24207, g18206, I24213, I24214, I24215, g18212;
wire g18218, I24226, I24227, I24228, g18225, I24234, I24235, I24236, g18231, I24251, I24252;
wire I24253, g18257, I24263, I24264, I24265, g18270, I24271, I24272, I24273, g18276, I24278;
wire I24279, I24280, g18277, I24290, I24291, I24292, g18290, I24298, I24299, I24300, g18296;
wire I24306, I24307, I24308, g18302, I24317, I24318, I24319, g18313, I24325, I24326, I24327;
wire g18319, g18325, I24338, I24339, I24340, g18332, I24351, I24352, I24353, g18346, I24361;
wire I24362, I24363, g18354, I24372, I24373, I24374, g18363, I24380, I24381, I24382, g18369;
wire I24387, I24388, I24389, g18370, I24399, I24400, I24401, g18383, I24407, I24408, I24409;
wire g18389, I24415, I24416, I24417, g18395, I24426, I24427, I24428, g18406, I24436, I24437;
wire I24438, g18419, I24443, I24444, I24445, g18424, I24452, I24453, I24454, g18431, I24464;
wire I24465, I24466, g18441, I24474, I24475, I24476, g18449, I24485, I24486, I24487, g18458;
wire I24493, I24494, I24495, g18464, I24500, I24501, I24502, g18465, I24512, I24513, I24514;
wire g18478, I24520, I24521, I24522, g18484, I24530, I24531, I24532, g18491, I24537, I24538;
wire I24539, g18492, I24544, I24545, I24546, g18497, I24553, I24554, I24555, g18504, I24565;
wire I24566, I24567, g18514, I24575, I24576, I24577, g18522, I24586, I24587, I24588, g18531;
wire I24594, I24595, I24596, g18537, I24601, I24602, I24603, g18538, I24611, I24612, I24613;
wire g18542, I24624, I24625, I24626, g18553, I24632, I24633, I24634, g18555, I24639, I24640;
wire I24641, g18556, I24646, I24647, I24648, g18561, I24655, I24656, I24657, g18568, I24667;
wire I24668, I24669, g18578, I24677, I24678, I24679, g18586, I24694, I24695, I24696, g18603;
wire I24702, I24703, I24704, g18605, I24709, I24710, I24711, g18606, I24716, I24717, I24718;
wire g18611, I24725, I24726, I24727, g18618, I24743, I24744, I24745, g18635, I24751, I24752;
wire I24753, g18637, I24763, I24764, I24765, g18644, g18977, I25030, I25031, I25032, g18980;
wire g19067, g19084, g19103, g19121, g19128, g19135, g19138, g19141, g19152, I25532, I25533;
wire I25534, g19261, I25539, I25540, I25541, g19262, I25560, I25561, I25562, g19271, I25571;
wire I25572, I25573, g19276, I25578, I25579, I25580, g19277, I25595, I25596, I25597, g19286;
wire g19288, I25605, I25606, I25607, g19290, I25616, I25617, I25618, g19295, I25623, I25624;
wire I25625, g19296, I25633, I25634, I25635, g19300, I25643, I25644, I25645, g19304, g19306;
wire I25653, I25654, I25655, g19308, I25664, I25665, I25666, g19313, I25671, I25672, I25673;
wire g19314, I25681, I25682, I25683, g19318, I25690, I25691, I25692, g19321, I25700, I25701;
wire I25702, g19325, g19327, I25710, I25711, I25712, g19329, I25721, I25722, I25723, g19334;
wire I25731, I25732, I25733, g19345, I25740, I25741, I25742, g19348, I25750, I25751, I25752;
wire g19352, g19354, I25761, I25762, I25763, g19357, I25771, I25772, I25773, g19368, I25781;
wire I25782, I25783, g19379, I25790, I25791, I25792, g19382, I25800, I25801, I25802, g19386;
wire I25809, I25810, I25811, g19389, I25819, I25820, I25821, g19400, I25829, I25830, I25831;
wire g19411, I25838, I25839, I25840, g19414, I25846, I25847, I25848, g19416, I25855, I25856;
wire I25857, g19419, I25865, I25866, I25867, g19430, I25880, I25881, I25882, g19451, I25888;
wire I25889, I25890, g19453, I25897, I25898, I25899, g19456, I25913, I25914, I25915, g19478;
wire I25921, I25922, I25923, g19480, I25938, I25939, I25940, g19501, g19865, g19896, g19921;
wire g19936, g19954, g19984, g20022, g20064, g20473, g20481, g20487, g20493, g20497, g20522;
wire g20537, g20542, g20633, g20648, g20658, g20672, g20683, g20693, g20700, g20703, g20707;
wire g20718, g20728, g20738, g20742, g20753, g20775, g20779, g20805, g20825, g21659, I28189;
wire I28190, I28191, g21660, g21685, g21686, g21688, I28217, I28218, I28219, g21689, g21714;
wire g21715, g21720, g21721, g21722, g21724, I28247, I28248, I28249, g21725, g21736, g21737;
wire g21740, g21741, g21746, g21747, g21748, g21750, I28271, I28272, I28273, g21751, g21759;
wire g21760, g21761, g21764, g21765, g21770, g21771, g21772, g21775, g21776, g21777, g21780;
wire g21781, g21786, g21790, g21791, g21792, g21804, g21848, g21850, g21855, g21857, g21858;
wire g21859, g21860, g21862, g21863, g21864, g21865, g21866, g21868, g21869, g21870, g21871;
wire g21873, g21874, g21875, g21877, g21879, g21881, g21885, g21888, g21903, g21976, g21983;
wire g21989, g21991, g21996, g22002, g22005, g22009, g22016, g22021, g22050, g22069, g22083;
wire g22093, g22108, g22118, g22134, g22157, I28726, I28727, I28728, g22188, I28741, I28742;
wire I28743, g22197, I28753, I28754, I28755, g22203, I28765, I28766, I28767, g22209, g22317;
wire g22339, g22342, g22362, g22365, g22381, g22382, g22385, g22396, g22397, g22399, g22400;
wire g22608, g22644, g22668, g22680, g22708, g22720, g22739, g22771, g22809, g22844, g22845;
wire g22846, g22850, g22876, g22879, g22880, g22881, g22885, g22911, g22914, g22915, g22916;
wire g22920, g22936, g22939, g22940, g22941, g22942, g22992, g23003, g23017, g23033, g23320;
wire g23325, g23331, g23335, g23340, g23344, g23349, g23353, g23360, g23364, g23368, g23372;
wire g23376, g23377, g23381, g23387, g23388, g23394, g23395, g23402, g23478, g23486, g23489;
wire g23495, g23502, g23505, g23511, g23518, g23521, g23526, g23533, g23537, I30790, I30791;
wire I30792, g23660, I30868, I30869, I30870, g23710, I30952, I30953, I30954, g23764, I31035;
wire I31036, I31037, g23819, g23906, g23936, g23937, g23938, g23953, g23968, g23969, g23970;
wire g23973, g23982, g23997, g23998, g23999, g24002, g24003, g24012, g24027, g24028, g24034;
wire g24036, g24037, g24046, g24052, g24054, g24056, g24057, g24058, g24065, g24067, g24069;
wire g24070, g24071, g24078, g24080, g24081, g24082, g24089, g24090, g24091, g24093, g24100;
wire g24109, g24126, g24145, g24442, g24443, g24444, g24447, g24448, g24449, g24450, g24451;
wire g24452, g24453, g24454, g24455, g24456, g24457, g24458, g24459, g24460, g24461, g24462;
wire g24463, g24464, g24465, g24466, g24467, g24468, g24469, g24470, g24471, g24472, g24474;
wire g24475, g24477, g24616, g24627, g24641, g24660, I32265, I32266, I32267, g24753, I32284;
wire I32285, I32286, g24766, I32295, I32296, I32297, g24771, I32308, I32309, I32310, g24778;
wire I32323, I32324, I32325, g24787, I32333, I32334, I32335, g24791, I32345, I32346, I32347;
wire g24797, I32355, I32356, I32357, g24801, I32368, I32369, I32370, g24808, I32378, I32379;
wire I32380, g24812, g24814, I32391, I32392, I32393, g24817, I32400, I32401, I32402, g24820;
wire I32409, I32410, I32411, g24823, I32422, I32423, I32424, g24830, I32430, I32431, I32432;
wire g24832, g24833, I32443, I32444, I32445, g24837, I32451, I32452, I32453, g24839, I32460;
wire I32461, I32462, g24842, I32468, I32469, I32470, g24844, I32478, I32479, I32480, g24848;
wire g24849, I32490, I32491, I32492, g24852, I32498, I32499, I32500, g24854, I32509, I32510;
wire I32511, g24857, I32518, I32519, I32520, g24860, I32526, I32527, I32528, g24862, g24863;
wire I32538, I32539, I32540, g24866, I32546, I32547, I32548, g24868, I32559, I32560, I32561;
wire g24873, I32567, I32568, I32569, g24875, I32575, I32576, I32577, g24877, I32586, I32587;
wire I32588, g24880, I32595, I32596, I32597, g24883, I32607, I32608, I32609, g24887, I32615;
wire I32616, I32617, g24889, I32624, I32625, I32626, g24897, I32633, I32634, I32635, g24900;
wire I32645, I32646, I32647, g24904, I32659, I32660, I32661, g24920, I32668, I32669, I32670;
wire g24923, I32677, I32678, I32679, g24928, I32686, I32687, I32688, g24937, I32695, I32696;
wire I32697, g24940, I32708, I32709, I32710, g24951, I32724, I32725, I32726, g24963, g24975;
wire g24986, g24997, g25004, g25005, g25008, g25009, g25010, g25011, g25012, g25013, g25014;
wire g25015, g25016, g25017, g25018, g25019, g25020, g25021, g25022, g25023, g25024, g25025;
wire g25026, g25028, g25029, g25030, g25031, g25032, g25033, g25034, g25035, g25036, g25037;
wire g25038, g25039, g25040, g25041, g25043, g25044, g25045, g25046, g25047, g25048, g25049;
wire g25050, g25051, g25052, g25053, g25054, g25055, g25057, g25058, g25059, g25060, g25061;
wire g25062, g25063, g25064, g25065, g25066, g25068, g25069, g25070, g25071, g25072, g25073;
wire g25074, g25088, g25096, g25106, g25112, g25200, g25203, g25205, g25210, g25312, g25320;
wire g25331, g25340, g25927, g25928, g25929, g25930, g25931, g25933, g25934, g25936, g25954;
wire g25958, g25964, g25969, g26059, g26066, g26073, g26079, g26106, g26119, g26120, g26129;
wire g26130, g26143, g26144, g26148, g26356, g26399, g26440, g26458, g26472, g26482, g26498;
wire g26513, g26772, g26779, g26785, g26792, I35020, I35021, I35022, g26859, I35034, I35035;
wire I35036, g26865, I35042, I35043, I35044, g26867, I35057, I35058, I35059, g26874, g26892;
wire g26902, g26906, g26911, g26915, g26918, g26925, g26928, g26931, I35123, I35124, I35125;
wire g26934, g26938, g26941, g26947, g27117, g27118, g27119, g27121, g27122, g27124, g27125;
wire g27130, I35701, I35702, I35703, g27379, I35714, I35715, I35716, g27382, g27390, g27395;
wire g27400, g27408, g27413, g27426, g27431, g27447, I35904, I35905, I35906, g27528, I35944;
wire I35945, I35946, g27550, I35974, I35975, I35976, g27566, g27571, I35992, I35993, I35994;
wire g27576, g27580, g27583, g27587, g27626, g27627, g27628, g27630, g27738, g27743, g27751;
wire g27756, I36256, I36257, I36258, g27801, I36270, I36271, I36272, g27809, I36289, I36290;
wire I36291, g27830, I36300, I36301, I36302, g27838, I36314, I36315, I36316, g27846, I36591;
wire I36592, I36593, g28046, I36666, I36667, I36668, g28075, I36731, I36732, I36733, g28100;
wire I36779, I36780, I36781, g28118, I37295, I37296, I37297, g28384, I37303, I37304, I37305;
wire g28386, I37311, I37312, I37313, g28388, I37322, I37323, I37324, g28391, I37356, I37357;
wire I37358, g28415, I37813, I37814, I37815, g28842, I37822, I37823, I37824, g28845, g28978;
wire g29001, g29008, g29026, g29030, g29038, g29045, g29049, g29053, g29060, g29062, g29068;
wire g29072, g29076, g29080, g29087, g29088, g29096, g29103, g29107, I38378, I38379, I38380;
wire g29265, I38810, I38811, I38812, g29498, I38820, I38821, I38822, g29500, I38831, I38832;
wire I38833, g29503, I38841, I38842, I38843, g29505, I39323, I39324, I39325, g29911, I39331;
wire I39332, I39333, g29913, I39339, I39340, I39341, g29915, I39347, I39348, I39349, g29917;
wire I39359, I39360, I39361, g29923, I39367, I39368, I39369, g29925, I39375, I39376, I39377;
wire g29927, I39384, I39385, I39386, g29930, I39391, I39392, I39393, g29931, I39532, I39533;
wire I39534, g30034, I39539, I39540, I39541, g30035, I39689, I39690, I39691, g30228, I40558;
wire I40559, I40560, g30768, I40571, I40572, I40573, g30771, I40587, I40588, I40589, g30775;
wire I40603, I40604, I40605, g30779, I40627, I40628, I40629, g30791, I41010, I41011, I41012;
wire g30926, I41017, I41018, I41019, g30927, I41064, I41065, I41066, g30952, g7528, g7575;
wire g7795, g8430, g10784, g10789, g10793, g10797, g10801, g10805, g10810, g10814, g10818;
wire g10822, g10831, g10835, g10839, g10851, g10855, g10872, g11600, g11622, g11624, g11627;
wire g11630, g11643, g11644, g11647, g11650, g11653, g11660, g11663, g11666, g11669, g11675;
wire g11678, g11681, g11687, g11690, g11697, g11703, g11711, g11744, g11759, g11760, g11767;
wire g11768, g11772, g11773, g11780, g11781, g11784, g11785, g11789, g11790, g11799, g11800;
wire g11806, g11807, g11810, g11811, g11815, g11822, g11823, g11828, g11830, g11831, g11832;
wire g11833, g11839, g11840, g11843, g11844, g11855, g11860, g11861, g11863, g11864, g11865;
wire g11870, g11872, g11873, g11874, g11875, g11881, g11882, g11889, g11890, g11896, g11897;
wire g11902, g11903, g11905, g11906, g11907, g11912, g11914, g11915, g11916, g11917, g11928;
wire g11934, g11935, g11938, g11939, g11940, g11946, g11947, g11952, g11953, g11955, g11956;
wire g11957, g11962, g11964, g11965, g11974, g11975, g11979, g11980, g11981, g11987, g11988;
wire g11991, g11992, g11993, g11999, g12000, g12005, g12006, g12008, g12026, g12033, g12034;
wire g12035, g12036, g12043, g12044, g12048, g12049, g12050, g12056, g12057, g12060, g12061;
wire g12062, g12068, g12079, g12080, g12081, g12082, g12083, g12090, g12097, g12098, g12099;
wire g12100, g12107, g12108, g12112, g12113, g12114, g12120, g12121, g12124, g12145, g12146;
wire g12151, g12152, g12153, g12154, g12155, g12162, g12169, g12170, g12171, g12172, g12179;
wire g12180, g12184, g12185, g12192, g12193, g12194, g12195, g12207, g12208, g12213, g12214;
wire g12215, g12216, g12217, g12224, g12231, g12232, g12233, g12234, g12245, g12247, g12248;
wire g12249, g12250, g12262, g12263, g12268, g12269, g12270, g12271, g12272, g12288, g12290;
wire g12291, g12292, g12293, g12305, g12306, g12324, g12326, g12327, g12328, g12329, g12339;
wire g12352, g12369, g12388, g12418, g12431, g12436, g12441, g12446, g12451, g12457, g12467;
wire g12482, g12487, g12499, g12507, g12524, g12539, g12698, g12747, g12755, g12780, g12781;
wire g12789, g12797, g12814, g12819, g12820, g12828, g12836, g12849, g12852, g12857, g12858;
wire g12866, g12880, g12883, g12890, g12893, g12898, g12899, g12912, g12913, g12920, g12923;
wire g12930, g12933, g12939, g12941, g12942, g12949, g12952, g12959, g12967, g12968, g12970;
wire g12971, g12978, g12981, g12991, g12992, g12994, g12995, g13001, g13002, g13022, g13024;
wire g13111, g13124, g13135, g13143, g13149, g13155, g13160, g13164, g13171, g13175, g13182;
wire g13194, g13228, g13251, g13274, g13286, g13299, g13310, g13313, g13331, g13332, g13353;
wire g13354, g13374, g13375, g13378, g13401, g13404, g15661, g15797, g15873, g15959, g15978;
wire g16020, g16036, g16058, g16082, g16094, g16120, g16171, g16230, g16498, g16520, g16551;
wire g16567, g16570, g16583, g16591, g16594, g16611, g16614, g16629, g16632, g16643, g16654;
wire g16655, g16671, g16672, g16679, g16692, g16693, g16705, g16718, g16736, g16778, g16802;
wire g16803, g16823, g16824, g16829, g16835, g16841, g16844, g16845, g16847, g16851, g16853;
wire g16854, g16857, g16860, g16861, g16866, g16880, g17012, g17025, g17042, g17051, g17059;
wire g17076, g17086, g17094, g17111, g17124, g17132, g17151, g17186, g17197, g17204, g17209;
wire g17213, g17215, g17216, g17218, g17219, g17220, g17221, g17222, g17223, g17224, g17225;
wire g17226, g17228, g17229, g17234, g17235, g17236, g17246, g17247, g17248, g17269, g17270;
wire g17271, g17302, g17303, g17340, g17341, g17383, g17429, g17507, g17896, g18007, g18085;
wire g18124, g18201, g18240, g18308, g18352, g18401, g18430, g18447, g18503, g18520, g18548;
wire g18567, g18584, g18590, g18598, g18617, g18623, g18626, g18630, g18639, g18669, g18678;
wire g18707, g18719, g18726, g18743, g18754, g18755, g18763, g18780, g18781, g18782, g18794;
wire g18803, g18804, g18820, g18821, g18835, g18836, g18837, g18852, g18866, g18867, g18868;
wire g18883, g18885, g18906, g18907, g18942, g18957, g18968, g18975, g19144, g19149, g19153;
wire g19154, g19157, g19160, g19162, g19163, g19165, g19167, g19171, g19172, g19173, g19177;
wire g19178, g19179, g19184, g19219, g20008, g20054, g20095, g20120, g20150, g20153, g20299;
wire g20310, g20314, g20318, g20333, g20337, g20343, g20353, g20357, g20375, g20376, g20417;
wire g20682, g20717, g20752, g20789, g20841, g20874, g20875, g20876, g20877, g20878, g20879;
wire g20880, g20881, g20882, g20883, g20884, g20891, g20892, g20893, g20894, g20895, g20896;
wire g20897, g20898, g20899, g20900, g20901, g20902, g20903, g20910, g20911, g20912, g20913;
wire g20914, g20915, g20916, g20917, g20918, g20919, g20920, g20921, g20922, g20923, g20924;
wire g20925, g20926, g20927, g20934, g20935, g20936, g20937, g20938, g20939, g20940, g20941;
wire g20944, g20945, g20946, g20947, g20948, g20949, g20950, g20951, g20952, g20953, g20954;
wire g20955, g20962, g20963, g20964, g20965, g20966, g20967, g20968, g20969, g20970, g20972;
wire g20973, g20974, g20975, g20976, g20977, g20978, g20979, g20980, g20981, g20982, g20983;
wire g20989, g20990, g20991, g20992, g20993, g20994, g20995, g20996, g20997, g20999, g21000;
wire g21001, g21002, g21003, g21004, g21005, g21006, g21007, g21008, g21009, g21010, g21011;
wire g21015, g21016, g21017, g21018, g21019, g21020, g21021, g21022, g21023, g21025, g21026;
wire g21027, g21028, g21029, g21031, g21032, g21033, g21034, g21035, g21039, g21040, g21041;
wire g21042, g21043, g21044, g21045, g21046, g21047, g21048, g21051, g21052, g21053, g21054;
wire g21055, g21056, g21060, g21061, g21062, g21063, g21065, g21070, g21071, g21072, g21073;
wire g21074, g21075, g21080, g21081, g21082, g21083, g21084, g21094, g21095, g21096, g21104;
wire g21105, g21106, g21116, g21117, g21118, g21119, g21133, g21134, g21135, g21147, g21148;
wire g21149, g21167, g21168, g21169, g21183, g21189, g21204, g21211, g21219, g21227, g21228;
wire g21230, g21233, g21235, g21238, g21242, g21246, g21250, g21255, g21263, g21316, g21331;
wire g21346, g21364, g21385, g21407, g21432, g21435, g21467, g21470, g21502, g21615, g21618;
wire g21636, g21643, g21646, g21665, g21667, g21674, g21677, g21694, g21696, g21703, g21706;
wire g21711, g21730, g21732, g21738, g21739, g21756, g21762, g21763, g21778, g21779, g21793;
wire g21794, g21796, g21842, g21843, g21845, g21847, g21851, g21878, g21880, g21882, g21884;
wire g21887, g21889, g21890, g21893, g21894, g21901, g21968, g21969, g21970, g21971, g21972;
wire g21973, g21974, g21975, g21980, g21981, g21987, g21988, g22000, g22001, g22013, g22025;
wire g22026, g22027, g22028, g22029, g22030, g22031, g22032, g22033, g22034, g22035, g22037;
wire g22038, g22039, g22040, g22041, g22042, g22043, g22044, g22045, g22047, g22048, g22049;
wire g22054, g22055, g22056, g22057, g22058, g22059, g22060, g22061, g22063, g22064, g22065;
wire g22066, g22067, g22068, g22073, g22074, g22075, g22076, g22077, g22078, g22079, g22080;
wire g22081, g22087, g22088, g22089, g22090, g22091, g22092, g22097, g22098, g22099, g22100;
wire g22101, g22102, g22103, g22104, g22105, g22106, g22112, g22113, g22114, g22115, g22116;
wire g22117, g22122, g22123, g22124, g22125, g22126, g22127, g22128, g22129, g22130, g22131;
wire g22132, g22138, g22139, g22140, g22141, g22142, g22143, g22144, g22145, g22146, g22147;
wire g22148, g22149, g22150, g22151, g22152, g22153, g22154, g22155, g22161, g22162, g22163;
wire g22164, g22165, g22166, g22167, g22168, g22169, g22170, g22171, g22172, g22173, g22174;
wire g22177, g22178, g22179, g22180, g22181, g22182, g22183, g22184, g22185, g22186, g22189;
wire g22191, g22192, g22193, g22194, g22195, g22198, g22200, g22204, g22210, g22216, g22218;
wire g22227, g22231, g22234, g22242, g22247, g22249, g22263, g22267, g22269, g22280, g22284;
wire g22288, g22299, g22308, g22336, g22361, g22454, g22493, g22536, g22576, g22578, g22615;
wire g22651, g22687, g22755, g22784, g22789, g22810, g22826, g22831, g22851, g22865, g22870;
wire g22886, g22900, g22921, g22935, g22953, g22985, g22987, g22990, g22997, g22999, g23000;
wire g23009, g23013, g23014, g23022, g23023, g23025, g23029, g23030, g23039, g23040, g23042;
wire g23046, g23047, g23051, g23058, g23059, g23061, g23066, g23067, g23070, g23076, g23077;
wire g23080, g23081, g23083, g23092, g23093, g23096, g23097, g23099, g23110, g23111, g23113;
wire g23114, g23117, g23123, g23124, g23126, g23132, g23133, g23135, g23136, g23137, g23324;
wire g23329, g23330, g23339, g23348, g23357, g23358, g23359, g23385, g23386, g23392, g23393;
wire g23399, g23400, g23401, g23406, g23407, g23408, g23413, g23418, g23427, g23433, g23461;
wire g23477, g23497, g23513, g23528, g23539, g23545, g23823, g23858, g23892, g23913, g23922;
wire g23945, g23950, g23954, g23974, g23979, g23983, g24004, g24009, g24013, g24038, g24043;
wire g24059, g24072, g24083, g24092, g24174, g24178, g24179, g24181, g24182, g24206, g24207;
wire g24208, g24209, g24212, g24213, g24214, g24215, g24216, g24218, g24219, g24222, g24223;
wire g24225, g24226, g24227, g24228, g24230, g24231, g24232, g24234, g24235, g24237, g24238;
wire g24242, g24243, g24249, g24250, g24426, g24428, g24430, g24434, g24438, g24445, g24446;
wire g24473, g24476, g24479, g24480, g24481, g24485, g24486, g24487, g24488, g24489, g24490;
wire g24491, g24492, g24493, g24494, g24495, g24496, g24497, g24498, g24499, g24500, g24501;
wire g24502, g24503, g24504, g24505, g24506, g24507, g24508, g24509, g24510, g24511, g24512;
wire g24513, g24514, g24515, g24516, g24517, g24519, g24520, g24521, g24522, g24523, g24524;
wire g24525, g24526, g24527, g24528, g24530, g24532, g24533, g24534, g24535, g24536, g24537;
wire g24538, g24543, g24545, g24546, g24547, g24548, g24555, g24557, g24558, g24566, g24575;
wire g24606, g24613, g24622, g24623, g24624, g24636, g24637, g24638, g24652, g24656, g24657;
wire g24663, g24675, g24681, g24682, g24694, g24708, g24711, g24717, g24720, g24728, g24731;
wire g24736, g24739, g24742, g24756, g24770, g24782, g24783, g24800, g24819, g24836, g24845;
wire g24847, g24859, g24871, g25027, g25042, g25056, g25067, g25075, g25076, g25077, g25078;
wire g25081, g25082, g25085, g25091, g25099, g25125, g25127, g25129, g25185, g25189, g25191;
wire g25194, g25197, g25199, g25201, g25202, g25204, g25206, g25207, g25208, g25209, g25211;
wire g25212, g25213, g25214, g25215, g25216, g25217, g25218, g25219, g25220, g25221, g25222;
wire g25223, g25224, g25225, g25226, g25227, g25228, g25229, g25230, g25231, g25232, g25233;
wire g25234, g25235, g25236, g25237, g25238, g25239, g25240, g25241, g25242, g25243, g25244;
wire g25245, g25246, g25247, g25248, g25249, g25250, g25251, g25252, g25253, g25254, g25255;
wire g25256, g25257, g25258, g25259, g25260, g25261, g25262, g25263, g25264, g25265, g25266;
wire g25267, g25268, g25270, g25271, g25272, g25273, g25279, g25280, g25288, g25311, g25343;
wire g25357, g25372, g25389, g25418, g25426, g25429, g25450, g25451, g25452, g25523, g25539;
wire g25569, g25589, g25605, g25631, g25648, g25668, g25684, g25699, g25708, g25725, g25745;
wire g25761, g25764, g25772, g25781, g25798, g25818, g25826, g25835, g25852, g25853, g25861;
wire g25870, g25873, g25874, g25882, g25885, g25887, g25890, g25892, g25932, g25935, g25938;
wire g25940, g25941, g25943, g25944, g25946, g25947, g25948, g25949, g25950, g25962, g25967;
wire g25974, g25979, g26025, g26031, g26037, g26041, g26042, g26043, g26044, g26045, g26046;
wire g26047, g26048, g26049, g26050, g26055, g26081, g26083, g26084, g26087, g26090, g26096;
wire g26099, g26103, g26107, g26110, g26113, g26126, g26137, g26140, g26145, g26151, g26154;
wire g26160, g26168, g26183, g26199, g26217, g26240, g26265, g26272, g26283, g26295, g26304;
wire g26327, g26336, g26374, g26417, g26529, g26530, g26531, g26532, g26534, g26541, g26545;
wire g26547, g26553, g26557, g26559, g26560, g26569, g26573, g26575, g26583, g26592, g26596;
wire g26607, g26616, g26630, g26655, g26659, g26660, g26661, g26664, g26665, g26666, g26667;
wire g26669, g26670, g26671, g26672, g26675, g26676, g26677, g26776, g26781, g26786, g26789;
wire g26795, g26798, g26799, g26800, g26801, g26802, g26803, g26804, g26805, g26806, g26807;
wire g26808, g26809, g26810, g26811, g26812, g26813, g26814, g26815, g26816, g26817, g26818;
wire g26820, g26821, g26822, g26823, g26824, g26825, g26826, g26827, g26869, g26873, g26877;
wire g26878, g26882, g26885, g26887, g26891, g26897, g26901, g26905, g26914, g26988, g26989;
wire g27011, g27012, g27037, g27038, g27051, g27065, g27066, g27078, g27094, g27106, g27120;
wire g27123, g27129, g27131, g27144, g27147, g27149, g27152, g27157, g27160, g27165, g27174;
wire g27175, g27179, g27184, g27188, g27243, g27250, g27251, g27252, g27253, g27254, g27255;
wire g27256, g27257, g27258, g27259, g27260, g27261, g27262, g27263, g27264, g27265, g27266;
wire g27267, g27268, g27269, g27270, g27271, g27272, g27273, g27274, g27275, g27276, g27277;
wire g27278, g27279, g27280, g27281, g27282, g27283, g27284, g27285, g27286, g27287, g27288;
wire g27289, g27290, g27291, g27292, g27293, g27294, g27295, g27296, g27297, g27298, g27299;
wire g27300, g27301, g27302, g27303, g27304, g27305, g27306, g27307, g27308, g27309, g27310;
wire g27311, g27312, g27313, g27314, g27315, g27316, g27317, g27318, g27319, g27320, g27321;
wire g27322, g27323, g27324, g27325, g27326, g27327, g27328, g27329, g27330, g27331, g27332;
wire g27333, g27334, g27335, g27336, g27337, g27338, g27339, g27340, g27341, g27342, g27343;
wire g27344, g27345, g27346, g27347, g27348, g27354, g27414, g27415, g27435, g27436, g27450;
wire g27454, g27455, g27462, g27464, g27466, g27470, g27471, g27478, g27481, g27482, g27485;
wire g27492, g27496, g27501, g27504, g27507, g27513, g27521, g27524, g27527, g27529, g27531;
wire g27532, g27538, g27546, g27549, g27551, g27558, g27563, g27564, g27565, g27567, g27572;
wire g27573, g27574, g27575, g27577, g27579, g27581, g27582, g27584, g27585, g27588, g27594;
wire g27603, g27612, g27621, g27629, g27631, g27655, g27658, g27672, g27678, g27682, g27718;
wire g27722, g27724, g27735, g27736, g27741, g27742, g27746, g27747, g27754, g27755, g27759;
wire g27760, g27761, g27762, g27763, g27764, g27765, g27766, g27767, g27768, g27769, g27771;
wire g27798, g27802, g27810, g27811, g27814, g27823, g27824, g27827, g27834, g27842, g27850;
wire g27854, g27855, g27864, g27865, g27868, g27869, g27875, g27882, g27883, g27886, g27892;
wire g27896, g27897, g27900, g27906, g27911, g27916, g27917, g27925, g27937, g27950, g27962;
wire g27964, g27980, g27997, g28002, g28029, g28059, g28088, g28145, g28146, g28147, g28148;
wire g28157, g28185, g28189, g28191, g28192, g28199, g28321, g28325, g28328, g28342, g28344;
wire g28345, g28346, g28348, g28349, g28350, g28351, g28352, g28353, g28354, g28355, g28356;
wire g28357, g28358, g28360, g28361, g28362, g28363, g28364, g28366, g28367, g28368, g28371;
wire g28392, g28394, g28397, g28400, g28403, g28406, g28409, g28410, g28413, g28414, g28417;
wire g28418, g28420, g28421, g28425, g28449, g28461, g28470, g28473, g28482, g28488, g28489;
wire g28490, g28495, g28499, g28523, g28525, g28528, g28551, g28578, g28606, g28634, g28635;
wire g28636, g28637, g28654, g28656, g28658, g28661, g28668, g28728, g28731, g28732, g28733;
wire g28735, g28736, g28737, g28738, g28739, g28744, g28745, g28746, g28747, g28748, g28749;
wire g28750, g28754, g28758, g28759, g28760, g28761, g28762, g28763, g28767, g28771, g28772;
wire g28773, g28774, g28778, g28782, g28783, g28784, g28788, g28789, g28790, g28794, g28795;
wire g28802, g28803, g28813, g28874, g28886, g28903, g28920, g28941, g28954, g28963, g28982;
wire g28987, g28990, g29009, g29013, g29016, g29031, g29039, g29063, g29064, g29083, g29090;
wire g29097, g29109, g29110, g29111, g29112, g29113, g29126, g29127, g29128, g29129, g29167;
wire g29169, g29170, g29172, g29173, g29178, g29179, g29181, g29182, g29184, g29185, g29187;
wire g29194, g29195, g29197, g29198, g29199, g29201, g29202, g29204, g29205, g29206, g29207;
wire g29209, g29210, g29212, g29213, g29214, g29215, g29216, g29218, g29219, g29221, g29222;
wire g29223, g29224, g29226, g29227, g29228, g29231, g29303, g29313, g29324, g29333, g29340;
wire g29343, g29345, g29347, g29353, g29354, g29355, g29357, g29399, g29403, g29406, g29409;
wire g29552, g29569, g29570, g29571, g29574, g29576, g29577, g29578, g29579, g29580, g29581;
wire g29582, g29606, g29608, g29609, g29611, g29612, g29613, g29616, g29617, g29618, g29620;
wire g29621, g29623, g29663, g29665, g29667, g29669, g29670, g29671, g29672, g29676, g29677;
wire g29678, g29679, g29680, g29681, g29682, g29683, g29684, g29685, g29686, g29687, g29688;
wire g29703, g29705, g29709, g29710, g29713, g29717, g29718, g29721, g29725, g29727, g29728;
wire g29731, g29732, g29735, g29736, g29740, g29741, g29744, g29747, g29748, g29751, g29754;
wire g29755, g29756, g29757, g29758, g29759, g29760, g29761, g29762, g29763, g29764, g29765;
wire g29766, g29767, g29768, g29769, g29770, g29771, g29772, g29773, g29774, g29775, g29776;
wire g29777, g29778, g29779, g29780, g29781, g29782, g29783, g29784, g29785, g29786, g29787;
wire g29788, g29789, g29791, g29912, g29914, g29916, g29918, g29919, g29920, g29921, g29922;
wire g29924, g29926, g29928, g29929, g29936, g29939, g29941, g30010, g30011, g30012, g30013;
wire g30014, g30015, g30016, g30017, g30018, g30019, g30020, g30021, g30022, g30023, g30024;
wire g30025, g30026, g30027, g30028, g30029, g30030, g30031, g30032, g30033, g30053, g30054;
wire g30055, g30056, g30057, g30058, g30059, g30060, g30061, g30062, g30063, g30064, g30065;
wire g30066, g30067, g30068, g30069, g30070, g30071, g30072, g30245, g30246, g30247, g30248;
wire g30249, g30250, g30251, g30252, g30253, g30254, g30255, g30256, g30257, g30258, g30259;
wire g30260, g30261, g30262, g30263, g30264, g30265, g30266, g30267, g30268, g30269, g30270;
wire g30271, g30272, g30273, g30274, g30275, g30276, g30277, g30278, g30279, g30280, g30281;
wire g30282, g30283, g30284, g30285, g30286, g30287, g30288, g30289, g30290, g30291, g30292;
wire g30293, g30294, g30295, g30296, g30297, g30298, g30299, g30300, g30301, g30302, g30303;
wire g30304, g30338, g30341, g30356, g30399, g30400, g30401, g30402, g30403, g30404, g30405;
wire g30406, g30455, g30468, g30470, g30482, g30485, g30487, g30500, g30503, g30505, g30566;
wire g30584, g30588, g30593, g30594, g30597, g30601, g30602, g30605, g30608, g30609, g30610;
wire g30613, g30614, g30617, g30618, g30621, g30622, g30625, g30628, g30629, g30632, g30635;
wire g30636, g30637, g30638, g30639, g30640, g30641, g30642, g30643, g30644, g30645, g30646;
wire g30647, g30648, g30649, g30650, g30651, g30652, g30653, g30654, g30655, g30656, g30657;
wire g30658, g30659, g30660, g30661, g30662, g30663, g30664, g30665, g30666, g30667, g30668;
wire g30669, g30670, g30671, g30672, g30673, g30674, g30675, g30676, g30677, g30678, g30679;
wire g30680, g30681, g30682, g30683, g30684, g30685, g30686, g30687, g30688, g30689, g30690;
wire g30691, g30692, g30693, g30694, g30695, g30699, g30700, g30701, g30702, g30703, g30704;
wire g30705, g30706, g30707, g30708, g30709, g30780, g30783, g30785, g30786, g30787, g30788;
wire g30789, g30790, g30796, g30798, g30801, g30929, g30930, g30931, g30932, g30933, g30934;
wire g30935, g30936, g30954, g30955, g30956, g30957, g30958, g30959, g30960, g30961, g30970;
wire line1, line2, line3, line4, line5, line6, line7, line8, line9, line10, line11;
wire line12, line13, line14, line15, line16, line17, line18, line19, line20, line21, line22;
wire line23, line24, line25, line26, line27, line28, line29, line30, line31, line32, line33;
wire line34, line35, line36, line37, line38, line39, line40, line41, line42, line43, line44;
wire line45, line46, line47, line48, line49, line50, line51, line52, line53, line54, line55;
wire line56, line57, line58, line59, line60, line61, line62, line63, line64, line65, line66;
wire line67, line68, line69, line70, line71, line72, line73, line74, line75, line76, line77;
wire line78, line79, line80, line81, line82, line83, line84, line85, line86, line87, line88;
wire line89, line90, line91, line92, line93, line94, line95, line96, line97, line98, line99;
wire line100, line101, line102, line103, line104, line105, line106, line107, line108, line109, line110;
wire line111, line112, line113, line114, line115, line116, line117, line118, line119, line120, line121;
wire line122, line123, line124, line125, line126, line127, line128, line129, line130, line131, line132;
wire line133, line134, line135, line136, line137, line138, line139, line140, line141, line142, line143;
wire line144, line145, line146, line147, line148, line149, line150, line151, line152, line153, line154;
wire line155, line156, line157, line158, line159, line160, line161, line162, line163, line164, line165;
wire line166, line167, line168, line169, line170, line171, line172, line173, line174, line175, line176;
wire line177, line178, line179, line180, line181, line182, line183, line184, line185, line186, line187;
wire line188, line189, line190, line191, line192, line193, line194, line195, line196, line197, line198;
wire line199, line200, line201, line202, line203, line204, line205, line206, line207, line208, line209;
wire line210, line211, line212, line213, line214, line215, line216, line217, line218, line219, line220;
wire line221, line222, line223, line224, line225, line226, line227, line228, line229, line230, line231;
wire line232, line233, line234, line235, line236, line237, line238, line239, line240, line241, line242;
wire line243, line244, line245, line246, line247, line248, line249, line250, line251, line252, line253;
wire line254, line255, line256, line257, line258, line259, line260, line261, line262, line263, line264;
wire line265, line266, line267, line268, line269, line270, line271, line272, line273, line274, line275;
wire line276, line277, line278, line279, line280, line281, line282, line283, line284, line285, line286;
wire line287, line288, line289, line290, line291, line292, line293, line294, line295, line296, line297;
wire line298, line299, line300, line301, line302, line303, line304, line305, line306, line307, line308;
wire line309, line310, line311, line312, line313, line314, line315, line316, line317, line318, line319;
wire line320, line321, line322, line323, line324, line325, line326, line327, line328, line329, line330;
wire line331, line332, line333, line334, line335, line336, line337, line338, line339, line340, line341;
wire line342, line343, line344, line345, line346, line347, line348, line349, line350, line351, line352;
wire line353, line354, line355, line356, line357, line358, line359, line360, line361, line362, line363;
wire line364, line365, line366, line367, line368, line369, line370, line371, line372, line373, line374;
wire line375, line376, line377, line378, line379, line380, line381, line382, line383, line384, line385;
wire line386, line387, line388, line389, line390, line391, line392, line393, line394, line395, line396;
wire line397, line398, line399, line400, line401, line402, line403, line404, line405, line406, line407;
wire line408, line409, line410, line411, line412, line413, line414, line415, line416, line417, line418;
wire line419, line420, line421, line422, line423, line424, line425, line426, line427, line428, line429;
wire line430, line431, line432, line433, line434, line435, line436, line437, line438, line439, line440;
wire line441, line442, line443, line444, line445, line446, line447, line448, line449, line450, line451;
wire line452, line453, line454, line455, line456, line457, line458, line459, line460, line461, line462;
wire line463, line464, line465, line466, line467, line468, line469, line470, line471, line472, line473;
wire line474, line475, line476, line477, line478, line479, line480, line481, line482, line483, line484;
wire line485, line486, line487, line488, line489, line490, line491, line492, line493, line494, line495;
wire line496, line497, line498, line499, line500, line501, line502, line503, line504, line505, line506;
wire line507, line508, line509, line510, line511, line512, line513, line514, line515, line516, line517;
wire line518, line519, line520, line521, line522, line523, line524, line525, line526, line527, line528;
wire line529, line530, line531, line532, line533, line534, line535, line536, line537, line538, line539;
wire line540, line541, line542, line543, line544, line545, line546, line547, line548, line549, line550;
wire line551, line552, line553, line554, line555, line556, line557, line558, line559, line560, line561;
wire line562, line563, line564, line565, line566, line567, line568, line569, line570, line571, line572;
wire line573, line574, line575, line576, line577, line578, line579, line580, line581, line582, line583;
wire line584, line585, line586, line587, line588, line589, line590, line591, line592, line593, line594;
wire line595, line596, line597, line598, line599, line600, line601, line602, line603, line604, line605;
wire line606, line607, line608, line609, line610, line611, line612, line613, line614, line615, line616;
wire line617, line618, line619, line620, line621, line622, line623, line624, line625, line626, line627;
wire line628, line629, line630, line631, line632, line633, line634, line635, line636, line637, line638;
wire line639, line640, line641, line642, line643, line644, line645, line646, line647, line648, line649;
wire line650, line651, line652, line653, line654, line655, line656, line657, line658, line659, line660;
wire line661, line662, line663, line664, line665, line666, line667, line668, line669, line670, line671;
wire line672, line673, line674, line675, line676, line677, line678, line679, line680, line681, line682;
wire line683, line684, line685, line686, line687, line688, line689, line690, line691, line692, line693;
wire line694, line695, line696, line697, line698, line699, line700, line701, line702, line703, line704;
wire line705, line706, line707, line708, line709, line710, line711, line712, line713, line714, line715;
wire line716, line717, line718, line719, line720, line721, line722, line723, line724, line725, line726;
wire line727, line728, line729, line730, line731, line732, line733, line734, line735, line736, line737;
wire line738, line739, line740, line741, line742, line743, line744, line745, line746, line747, line748;
wire line749, line750, line751, line752, line753, line754, line755, line756, line757, line758, line759;
wire line760, line761, line762, line763, line764, line765, line766, line767, line768, line769, line770;
wire line771, line772, line773, line774, line775, line776, line777, line778, line779, line780, line781;
wire line782, line783, line784, line785, line786, line787, line788, line789, line790, line791, line792;
wire line793, line794, line795, line796, line797, line798, line799, line800, line801, line802, line803;
wire line804, line805, line806, line807, line808, line809, line810, line811, line812, line813, line814;
wire line815, line816, line817, line818, line819, line820, line821, line822, line823, line824, line825;
wire line826, line827, line828, line829, line830, line831, line832, line833, line834, line835, line836;
wire line837, line838, line839, line840, line841, line842, line843, line844, line845, line846, line847;
wire line848, line849, line850, line851, line852, line853, line854, line855, line856, line857, line858;
wire line859, line860, line861, line862, line863, line864, line865, line866, line867, line868, line869;
wire line870, line871, line872, line873, line874, line875, line876, line877, line878, line879, line880;
wire line881, line882, line883, line884, line885, line886, line887, line888, line889, line890, line891;
wire line892, line893, line894, line895, line896, line897, line898, line899, line900, line901, line902;
wire line903, line904, line905, line906, line907, line908, line909, line910, line911, line912, line913;
wire line914, line915, line916, line917, line918, line919, line920, line921, line922, line923, line924;
wire line925, line926, line927, line928, line929, line930, line931, line932, line933, line934, line935;
wire line936, line937, line938, line939, line940, line941, line942, line943, line944, line945, line946;
wire line947, line948, line949, line950, line951, line952, line953, line954, line955, line956, line957;
wire line958, line959, line960, line961, line962, line963, line964, line965, line966, line967, line968;
wire line969, line970, line971, line972, line973, line974, line975, line976, line977, line978, line979;
wire line980, line981, line982, line983, line984, line985, line986, line987, line988, line989, line990;
wire line991, line992, line993, line994, line995, line996, line997, line998, line999, line1000, line1001;
wire line1002, line1003, line1004, line1005, line1006, line1007, line1008, line1009, line1010, line1011, line1012;
wire line1013, line1014, line1015, line1016, line1017, line1018, line1019, line1020, line1021, line1022, line1023;
wire line1024, line1025, line1026, line1027, line1028, line1029, line1030, line1031, line1032, line1033, line1034;
wire line1035, line1036, line1037, line1038, line1039, line1040, line1041, line1042, line1043, line1044, line1045;
wire line1046, line1047, line1048, line1049, line1050, line1051, line1052, line1053, line1054, line1055, line1056;
wire line1057, line1058, line1059, line1060, line1061, line1062, line1063, line1064, line1065, line1066, line1067;
wire line1068, line1069, line1070, line1071, line1072, line1073, line1074, line1075, line1076, line1077, line1078;
wire line1079, line1080, line1081, line1082, line1083, line1084, line1085, line1086, line1087, line1088, line1089;
wire line1090, line1091, line1092, line1093, line1094, line1095, line1096, line1097, line1098, line1099, line1100;
wire line1101, line1102, line1103, line1104, line1105, line1106, line1107, line1108, line1109, line1110, line1111;
wire line1112, line1113, line1114, line1115, line1116, line1117, line1118, line1119, line1120, line1121, line1122;
wire line1123, line1124, line1125, line1126, line1127, line1128, line1129, line1130, line1131, line1132, line1133;
wire line1134, line1135, line1136, line1137, line1138, line1139, line1140, line1141, line1142, line1143, line1144;
wire line1145, line1146, line1147, line1148, line1149, line1150, line1151, line1152, line1153, line1154, line1155;
wire line1156, line1157, line1158, line1159, line1160, line1161, line1162, line1163, line1164, line1165, line1166;
wire line1167, line1168, line1169, line1170, line1171, line1172, line1173, line1174, line1175, line1176, line1177;
wire line1178, line1179, line1180, line1181, line1182, line1183, line1184, line1185, line1186, line1187, line1188;
wire line1189, line1190, line1191, line1192, line1193, line1194, line1195, line1196, line1197, line1198, line1199;
wire line1200, line1201, line1202, line1203, line1204, line1205, line1206, line1207, line1208, line1209, line1210;
wire line1211, line1212, line1213, line1214, line1215, line1216, line1217, line1218, line1219, line1220, line1221;
wire line1222, line1223, line1224, line1225, line1226, line1227, line1228, line1229, line1230, line1231, line1232;
wire line1233, line1234, line1235, line1236, line1237, line1238, line1239, line1240, line1241, line1242, line1243;
wire line1244, line1245, line1246, line1247, line1248, line1249, line1250, line1251, line1252, line1253, line1254;
wire line1255, line1256, line1257, line1258, line1259, line1260, line1261, line1262, line1263, line1264, line1265;
wire line1266, line1267, line1268, line1269, line1270, line1271, line1272, line1273, line1274, line1275, line1276;
wire line1277, line1278, line1279, line1280, line1281, line1282, line1283, line1284, line1285, line1286, line1287;
wire line1288, line1289, line1290, line1291, line1292, line1293, line1294, line1295, line1296, line1297, line1298;
wire line1299, line1300, line1301, line1302, line1303, line1304, line1305, line1306, line1307, line1308, line1309;
wire line1310, line1311, line1312, line1313, line1314, line1315, line1316, line1317, line1318, line1319, line1320;
wire line1321, line1322, line1323, line1324, line1325, line1326, line1327, line1328, line1329, line1330, line1331;
wire line1332, line1333, line1334, line1335, line1336, line1337, line1338, line1339, line1340, line1341, line1342;
wire line1343, line1344, line1345, line1346, line1347, line1348, line1349, line1350, line1351, line1352, line1353;
wire line1354, line1355, line1356, line1357, line1358, line1359, line1360, line1361, line1362, line1363, line1364;
wire line1365, line1366, line1367, line1368, line1369, line1370, line1371, line1372, line1373, line1374, line1375;
wire line1376, line1377, line1378, line1379, line1380, line1381, line1382, line1383, line1384, line1385, line1386;
wire line1387, line1388, line1389, line1390, line1391, line1392, line1393, line1394, line1395, line1396, line1397;
wire line1398, line1399, line1400, line1401, line1402, line1403, line1404, line1405, line1406, line1407, line1408;
wire line1409, line1410, line1411, line1412, line1413, line1414, line1415, line1416, line1417, line1418, line1419;
wire line1420, line1421, line1422, line1423, line1424, line1425, line1426, line1427, line1428, line1429, line1430;
wire line1431, line1432, line1433, line1434, line1435, line1436, line1437, line1438, line1439, line1440, line1441;
wire line1442, line1443, line1444, line1445, line1446, line1447, line1448, line1449, line1450, line1451, line1452;
wire line1453, line1454, line1455, line1456, line1457, line1458, line1459, line1460, line1461, line1462, line1463;
wire line1464, line1465, line1466, line1467, line1468, line1469, line1470, line1471, line1472, line1473, line1474;
wire line1475, line1476, line1477, line1478, line1479, line1480, line1481, line1482, line1483, line1484, line1485;
wire line1486, line1487, line1488, line1489, line1490, line1491, line1492, line1493, line1494, line1495, line1496;
wire line1497, line1498, line1499, line1500, line1501, line1502, line1503, line1504, line1505, line1506, line1507;
wire line1508, line1509, line1510, line1511, line1512, line1513, line1514, line1515, line1516, line1517, line1518;
wire line1519, line1520, line1521, line1522, line1523, line1524, line1525, line1526, line1527, line1528, line1529;
wire line1530, line1531, line1532, line1533, line1534, line1535, line1536, line1537, line1538, line1539, line1540;
wire line1541, line1542, line1543, line1544, line1545, line1546, line1547, line1548, line1549, line1550, line1551;
wire line1552, line1553, line1554, line1555, line1556, line1557, line1558, line1559, line1560, line1561, line1562;
wire line1563, line1564, line1565, line1566, line1567, line1568, line1569, line1570, line1571, line1572, line1573;
wire line1574, line1575, line1576, line1577, line1578, line1579, line1580, line1581, line1582, line1583, line1584;
wire line1585, line1586, line1587, line1588, line1589, line1590, line1591, line1592, line1593, line1594, line1595;
wire line1596, line1597, line1598, line1599, line1600, line1601, line1602, line1603, line1604, line1605, line1606;
wire line1607, line1608, line1609, line1610, line1611, line1612, line1613, line1614, line1615, line1616, line1617;
wire line1618, line1619, line1620, line1621, line1622, line1623, line1624, line1625, line1626, line1627, line1628;
wire line1629, line1630, line1631, line1632, line1633, line1634, line1635, line1636;
DFFX1 gate1(.Q (g2814), .QB (line1), .D(g16475), .CK(clk));
DFFX1 gate2(.Q (g2817), .QB (line2), .D(g20571), .CK(clk));
DFFX1 gate3(.Q (g2933), .QB (line3), .D(g20588), .CK(clk));
DFFX1 gate4(.Q (g2950), .QB (line4), .D(g21951), .CK(clk));
DFFX1 gate5(.Q (g2883), .QB (line5), .D(g23315), .CK(clk));
DFFX1 gate6(.Q (g2888), .QB (line6), .D(g24423), .CK(clk));
DFFX1 gate7(.Q (g2896), .QB (line7), .D(g25175), .CK(clk));
DFFX1 gate8(.Q (g2892), .QB (line8), .D(g26019), .CK(clk));
DFFX1 gate9(.Q (g2903), .QB (line9), .D(g26747), .CK(clk));
DFFX1 gate10(.Q (g2900), .QB (line10), .D(g27237), .CK(clk));
DFFX1 gate11(.Q (g2908), .QB (line11), .D(g27715), .CK(clk));
DFFX1 gate12(.Q (g2912), .QB (line12), .D(g24424), .CK(clk));
DFFX1 gate13(.Q (g2917), .QB (line13), .D(g25174), .CK(clk));
DFFX1 gate14(.Q (g2924), .QB (line14), .D(g26020), .CK(clk));
DFFX1 gate15(.Q (g2920), .QB (line15), .D(g26746), .CK(clk));
DFFX1 gate16(.Q (g2984), .QB (line16), .D(g19061), .CK(clk));
DFFX1 gate17(.Q (g2985), .QB (line17), .D(g19060), .CK(clk));
DFFX1 gate18(.Q (g2930), .QB (line18), .D(g19062), .CK(clk));
DFFX1 gate19(.Q (g2929), .QB (line19), .D(g2930), .CK(clk));
DFFX1 gate20(.Q (g2879), .QB (line20), .D(g16494), .CK(clk));
DFFX1 gate21(.Q (g2934), .QB (line21), .D(g16476), .CK(clk));
DFFX1 gate22(.Q (g2935), .QB (line22), .D(g16477), .CK(clk));
DFFX1 gate23(.Q (g2938), .QB (line23), .D(g16478), .CK(clk));
DFFX1 gate24(.Q (g2941), .QB (line24), .D(g16479), .CK(clk));
DFFX1 gate25(.Q (g2944), .QB (line25), .D(g16480), .CK(clk));
DFFX1 gate26(.Q (g2947), .QB (line26), .D(g16481), .CK(clk));
DFFX1 gate27(.Q (g2953), .QB (line27), .D(g16482), .CK(clk));
DFFX1 gate28(.Q (g2956), .QB (line28), .D(g16483), .CK(clk));
DFFX1 gate29(.Q (g2959), .QB (line29), .D(g16484), .CK(clk));
DFFX1 gate30(.Q (g2962), .QB (line30), .D(g16485), .CK(clk));
DFFX1 gate31(.Q (g2963), .QB (line31), .D(g16486), .CK(clk));
DFFX1 gate32(.Q (g2966), .QB (line32), .D(g16487), .CK(clk));
DFFX1 gate33(.Q (g2969), .QB (line33), .D(g16488), .CK(clk));
DFFX1 gate34(.Q (g2972), .QB (line34), .D(g16489), .CK(clk));
DFFX1 gate35(.Q (g2975), .QB (line35), .D(g16490), .CK(clk));
DFFX1 gate36(.Q (g2978), .QB (line36), .D(g16491), .CK(clk));
DFFX1 gate37(.Q (g2981), .QB (line37), .D(g16492), .CK(clk));
DFFX1 gate38(.Q (g2874), .QB (line38), .D(g16493), .CK(clk));
DFFX1 gate39(.Q (g1506), .QB (line39), .D(g20572), .CK(clk));
DFFX1 gate40(.Q (g1501), .QB (line40), .D(g20573), .CK(clk));
DFFX1 gate41(.Q (g1496), .QB (line41), .D(g20574), .CK(clk));
DFFX1 gate42(.Q (g1491), .QB (line42), .D(g20575), .CK(clk));
DFFX1 gate43(.Q (g1486), .QB (line43), .D(g20576), .CK(clk));
DFFX1 gate44(.Q (g1481), .QB (line44), .D(g20577), .CK(clk));
DFFX1 gate45(.Q (g1476), .QB (line45), .D(g20578), .CK(clk));
DFFX1 gate46(.Q (g1471), .QB (line46), .D(g20579), .CK(clk));
DFFX1 gate47(.Q (g2877), .QB (line47), .D(g23313), .CK(clk));
DFFX1 gate48(.Q (g2861), .QB (line48), .D(g21960), .CK(clk));
DFFX1 gate49(.Q (g813), .QB (line49), .D(g2861), .CK(clk));
DFFX1 gate50(.Q (g2864), .QB (line50), .D(g21961), .CK(clk));
DFFX1 gate51(.Q (g809), .QB (line51), .D(g2864), .CK(clk));
DFFX1 gate52(.Q (g2867), .QB (line52), .D(g21962), .CK(clk));
DFFX1 gate53(.Q (g805), .QB (line53), .D(g2867), .CK(clk));
DFFX1 gate54(.Q (g2870), .QB (line54), .D(g21963), .CK(clk));
DFFX1 gate55(.Q (g801), .QB (line55), .D(g2870), .CK(clk));
DFFX1 gate56(.Q (g2818), .QB (line56), .D(g21947), .CK(clk));
DFFX1 gate57(.Q (g797), .QB (line57), .D(g2818), .CK(clk));
DFFX1 gate58(.Q (g2821), .QB (line58), .D(g21948), .CK(clk));
DFFX1 gate59(.Q (g793), .QB (line59), .D(g2821), .CK(clk));
DFFX1 gate60(.Q (g2824), .QB (line60), .D(g21949), .CK(clk));
DFFX1 gate61(.Q (g789), .QB (line61), .D(g2824), .CK(clk));
DFFX1 gate62(.Q (g2827), .QB (line62), .D(g21950), .CK(clk));
DFFX1 gate63(.Q (g785), .QB (line63), .D(g2827), .CK(clk));
DFFX1 gate64(.Q (g2830), .QB (line64), .D(g23312), .CK(clk));
DFFX1 gate65(.Q (g2873), .QB (line65), .D(g2830), .CK(clk));
DFFX1 gate66(.Q (g2833), .QB (line66), .D(g21952), .CK(clk));
DFFX1 gate67(.Q (g125), .QB (line67), .D(g2833), .CK(clk));
DFFX1 gate68(.Q (g2836), .QB (line68), .D(g21953), .CK(clk));
DFFX1 gate69(.Q (g121), .QB (line69), .D(g2836), .CK(clk));
DFFX1 gate70(.Q (g2839), .QB (line70), .D(g21954), .CK(clk));
DFFX1 gate71(.Q (g117), .QB (line71), .D(g2839), .CK(clk));
DFFX1 gate72(.Q (g2842), .QB (line72), .D(g21955), .CK(clk));
DFFX1 gate73(.Q (g113), .QB (line73), .D(g2842), .CK(clk));
DFFX1 gate74(.Q (g2845), .QB (line74), .D(g21956), .CK(clk));
DFFX1 gate75(.Q (g109), .QB (line75), .D(g2845), .CK(clk));
DFFX1 gate76(.Q (g2848), .QB (line76), .D(g21957), .CK(clk));
DFFX1 gate77(.Q (g105), .QB (line77), .D(g2848), .CK(clk));
DFFX1 gate78(.Q (g2851), .QB (line78), .D(g21958), .CK(clk));
DFFX1 gate79(.Q (g101), .QB (line79), .D(g2851), .CK(clk));
DFFX1 gate80(.Q (g2854), .QB (line80), .D(g21959), .CK(clk));
DFFX1 gate81(.Q (g97), .QB (line81), .D(g2854), .CK(clk));
DFFX1 gate82(.Q (g2858), .QB (line82), .D(g23316), .CK(clk));
DFFX1 gate83(.Q (g2857), .QB (line83), .D(g2858), .CK(clk));
DFFX1 gate84(.Q (g2200), .QB (line84), .D(g20587), .CK(clk));
DFFX1 gate85(.Q (g2195), .QB (line85), .D(g20585), .CK(clk));
DFFX1 gate86(.Q (g2190), .QB (line86), .D(g20586), .CK(clk));
DFFX1 gate87(.Q (g2185), .QB (line87), .D(g20584), .CK(clk));
DFFX1 gate88(.Q (g2180), .QB (line88), .D(g20583), .CK(clk));
DFFX1 gate89(.Q (g2175), .QB (line89), .D(g20582), .CK(clk));
DFFX1 gate90(.Q (g2170), .QB (line90), .D(g20581), .CK(clk));
DFFX1 gate91(.Q (g2165), .QB (line91), .D(g20580), .CK(clk));
DFFX1 gate92(.Q (g2878), .QB (line92), .D(g23314), .CK(clk));
DFFX1 gate93(.Q (g3129), .QB (line93), .D(g13475), .CK(clk));
DFFX1 gate94(.Q (g3117), .QB (line94), .D(g3129), .CK(clk));
DFFX1 gate95(.Q (g3109), .QB (line95), .D(g3117), .CK(clk));
DFFX1 gate96(.Q (g3210), .QB (line96), .D(g20630), .CK(clk));
DFFX1 gate97(.Q (g3211), .QB (line97), .D(g20631), .CK(clk));
DFFX1 gate98(.Q (g3084), .QB (line98), .D(g20632), .CK(clk));
DFFX1 gate99(.Q (g3085), .QB (line99), .D(g20609), .CK(clk));
DFFX1 gate100(.Q (g3086), .QB (line100), .D(g20610), .CK(clk));
DFFX1 gate101(.Q (g3087), .QB (line101), .D(g20611), .CK(clk));
DFFX1 gate102(.Q (g3091), .QB (line102), .D(g20612), .CK(clk));
DFFX1 gate103(.Q (g3092), .QB (line103), .D(g20613), .CK(clk));
DFFX1 gate104(.Q (g3093), .QB (line104), .D(g20614), .CK(clk));
DFFX1 gate105(.Q (g3094), .QB (line105), .D(g20615), .CK(clk));
DFFX1 gate106(.Q (g3095), .QB (line106), .D(g20616), .CK(clk));
DFFX1 gate107(.Q (g3096), .QB (line107), .D(g20617), .CK(clk));
DFFX1 gate108(.Q (g3097), .QB (line108), .D(g26751), .CK(clk));
DFFX1 gate109(.Q (g3098), .QB (line109), .D(g26752), .CK(clk));
DFFX1 gate110(.Q (g3099), .QB (line110), .D(g26753), .CK(clk));
DFFX1 gate111(.Q (g3100), .QB (line111), .D(g29163), .CK(clk));
DFFX1 gate112(.Q (g3101), .QB (line112), .D(g29164), .CK(clk));
DFFX1 gate113(.Q (g3102), .QB (line113), .D(g29165), .CK(clk));
DFFX1 gate114(.Q (g3103), .QB (line114), .D(g30120), .CK(clk));
DFFX1 gate115(.Q (g3104), .QB (line115), .D(g30121), .CK(clk));
DFFX1 gate116(.Q (g3105), .QB (line116), .D(g30122), .CK(clk));
DFFX1 gate117(.Q (g3106), .QB (line117), .D(g30941), .CK(clk));
DFFX1 gate118(.Q (g3107), .QB (line118), .D(g30942), .CK(clk));
DFFX1 gate119(.Q (g3108), .QB (line119), .D(g30943), .CK(clk));
DFFX1 gate120(.Q (g3155), .QB (line120), .D(g20618), .CK(clk));
DFFX1 gate121(.Q (g3158), .QB (line121), .D(g20619), .CK(clk));
DFFX1 gate122(.Q (g3161), .QB (line122), .D(g20620), .CK(clk));
DFFX1 gate123(.Q (g3164), .QB (line123), .D(g20621), .CK(clk));
DFFX1 gate124(.Q (g3167), .QB (line124), .D(g20622), .CK(clk));
DFFX1 gate125(.Q (g3170), .QB (line125), .D(g20623), .CK(clk));
DFFX1 gate126(.Q (g3173), .QB (line126), .D(g20624), .CK(clk));
DFFX1 gate127(.Q (g3176), .QB (line127), .D(g20625), .CK(clk));
DFFX1 gate128(.Q (g3179), .QB (line128), .D(g20626), .CK(clk));
DFFX1 gate129(.Q (g3182), .QB (line129), .D(g20627), .CK(clk));
DFFX1 gate130(.Q (g3185), .QB (line130), .D(g20628), .CK(clk));
DFFX1 gate131(.Q (g3088), .QB (line131), .D(g20629), .CK(clk));
DFFX1 gate132(.Q (g3191), .QB (line132), .D(g27717), .CK(clk));
DFFX1 gate133(.Q (g3194), .QB (line133), .D(g28316), .CK(clk));
DFFX1 gate134(.Q (g3197), .QB (line134), .D(g28317), .CK(clk));
DFFX1 gate135(.Q (g3198), .QB (line135), .D(g28318), .CK(clk));
DFFX1 gate136(.Q (g3201), .QB (line136), .D(g28704), .CK(clk));
DFFX1 gate137(.Q (g3204), .QB (line137), .D(g28705), .CK(clk));
DFFX1 gate138(.Q (g3207), .QB (line138), .D(g28706), .CK(clk));
DFFX1 gate139(.Q (g3188), .QB (line139), .D(g29463), .CK(clk));
DFFX1 gate140(.Q (g3133), .QB (line140), .D(g29656), .CK(clk));
DFFX1 gate141(.Q (g3132), .QB (line141), .D(g28698), .CK(clk));
DFFX1 gate142(.Q (g3128), .QB (line142), .D(g29166), .CK(clk));
DFFX1 gate143(.Q (g3127), .QB (line143), .D(g28697), .CK(clk));
DFFX1 gate144(.Q (g3126), .QB (line144), .D(g28315), .CK(clk));
DFFX1 gate145(.Q (g3125), .QB (line145), .D(g28696), .CK(clk));
DFFX1 gate146(.Q (g3124), .QB (line146), .D(g28314), .CK(clk));
DFFX1 gate147(.Q (g3123), .QB (line147), .D(g28313), .CK(clk));
DFFX1 gate148(.Q (g3120), .QB (line148), .D(g28695), .CK(clk));
DFFX1 gate149(.Q (g3114), .QB (line149), .D(g28694), .CK(clk));
DFFX1 gate150(.Q (g3113), .QB (line150), .D(g28693), .CK(clk));
DFFX1 gate151(.Q (g3112), .QB (line151), .D(g28312), .CK(clk));
DFFX1 gate152(.Q (g3110), .QB (line152), .D(g28311), .CK(clk));
DFFX1 gate153(.Q (g3111), .QB (line153), .D(g28310), .CK(clk));
DFFX1 gate154(.Q (g3139), .QB (line154), .D(g29461), .CK(clk));
DFFX1 gate155(.Q (g3136), .QB (line155), .D(g28701), .CK(clk));
DFFX1 gate156(.Q (g3134), .QB (line156), .D(g28700), .CK(clk));
DFFX1 gate157(.Q (g3135), .QB (line157), .D(g28699), .CK(clk));
DFFX1 gate158(.Q (g3151), .QB (line158), .D(g29462), .CK(clk));
DFFX1 gate159(.Q (g3142), .QB (line159), .D(g28703), .CK(clk));
DFFX1 gate160(.Q (g3147), .QB (line160), .D(g28702), .CK(clk));
DFFX1 gate161(.Q (g185), .QB (line161), .D(g29657), .CK(clk));
DFFX1 gate162(.Q (g138), .QB (line162), .D(g13405), .CK(clk));
DFFX1 gate163(.Q (g135), .QB (line163), .D(g138), .CK(clk));
DFFX1 gate164(.Q (g165), .QB (line164), .D(g135), .CK(clk));
DFFX1 gate165(.Q (g130), .QB (line165), .D(g24259), .CK(clk));
DFFX1 gate166(.Q (g131), .QB (line166), .D(g24260), .CK(clk));
DFFX1 gate167(.Q (g129), .QB (line167), .D(g24261), .CK(clk));
DFFX1 gate168(.Q (g133), .QB (line168), .D(g24262), .CK(clk));
DFFX1 gate169(.Q (g134), .QB (line169), .D(g24263), .CK(clk));
DFFX1 gate170(.Q (g132), .QB (line170), .D(g24264), .CK(clk));
DFFX1 gate171(.Q (g142), .QB (line171), .D(g24265), .CK(clk));
DFFX1 gate172(.Q (g143), .QB (line172), .D(g24266), .CK(clk));
DFFX1 gate173(.Q (g141), .QB (line173), .D(g24267), .CK(clk));
DFFX1 gate174(.Q (g145), .QB (line174), .D(g24268), .CK(clk));
DFFX1 gate175(.Q (g146), .QB (line175), .D(g24269), .CK(clk));
DFFX1 gate176(.Q (g144), .QB (line176), .D(g24270), .CK(clk));
DFFX1 gate177(.Q (g148), .QB (line177), .D(g24271), .CK(clk));
DFFX1 gate178(.Q (g149), .QB (line178), .D(g24272), .CK(clk));
DFFX1 gate179(.Q (g147), .QB (line179), .D(g24273), .CK(clk));
DFFX1 gate180(.Q (g151), .QB (line180), .D(g24274), .CK(clk));
DFFX1 gate181(.Q (g152), .QB (line181), .D(g24275), .CK(clk));
DFFX1 gate182(.Q (g150), .QB (line182), .D(g24276), .CK(clk));
DFFX1 gate183(.Q (g154), .QB (line183), .D(g24277), .CK(clk));
DFFX1 gate184(.Q (g155), .QB (line184), .D(g24278), .CK(clk));
DFFX1 gate185(.Q (g153), .QB (line185), .D(g24279), .CK(clk));
DFFX1 gate186(.Q (g157), .QB (line186), .D(g24280), .CK(clk));
DFFX1 gate187(.Q (g158), .QB (line187), .D(g24281), .CK(clk));
DFFX1 gate188(.Q (g156), .QB (line188), .D(g24282), .CK(clk));
DFFX1 gate189(.Q (g160), .QB (line189), .D(g24283), .CK(clk));
DFFX1 gate190(.Q (g161), .QB (line190), .D(g24284), .CK(clk));
DFFX1 gate191(.Q (g159), .QB (line191), .D(g24285), .CK(clk));
DFFX1 gate192(.Q (g163), .QB (line192), .D(g24286), .CK(clk));
DFFX1 gate193(.Q (g164), .QB (line193), .D(g24287), .CK(clk));
DFFX1 gate194(.Q (g162), .QB (line194), .D(g24288), .CK(clk));
DFFX1 gate195(.Q (g169), .QB (line195), .D(g26679), .CK(clk));
DFFX1 gate196(.Q (g170), .QB (line196), .D(g26680), .CK(clk));
DFFX1 gate197(.Q (g168), .QB (line197), .D(g26681), .CK(clk));
DFFX1 gate198(.Q (g172), .QB (line198), .D(g26682), .CK(clk));
DFFX1 gate199(.Q (g173), .QB (line199), .D(g26683), .CK(clk));
DFFX1 gate200(.Q (g171), .QB (line200), .D(g26684), .CK(clk));
DFFX1 gate201(.Q (g175), .QB (line201), .D(g26685), .CK(clk));
DFFX1 gate202(.Q (g176), .QB (line202), .D(g26686), .CK(clk));
DFFX1 gate203(.Q (g174), .QB (line203), .D(g26687), .CK(clk));
DFFX1 gate204(.Q (g178), .QB (line204), .D(g26688), .CK(clk));
DFFX1 gate205(.Q (g179), .QB (line205), .D(g26689), .CK(clk));
DFFX1 gate206(.Q (g177), .QB (line206), .D(g26690), .CK(clk));
DFFX1 gate207(.Q (g186), .QB (line207), .D(g30506), .CK(clk));
DFFX1 gate208(.Q (g189), .QB (line208), .D(g30507), .CK(clk));
DFFX1 gate209(.Q (g192), .QB (line209), .D(g30508), .CK(clk));
DFFX1 gate210(.Q (g231), .QB (line210), .D(g30842), .CK(clk));
DFFX1 gate211(.Q (g234), .QB (line211), .D(g30843), .CK(clk));
DFFX1 gate212(.Q (g237), .QB (line212), .D(g30844), .CK(clk));
DFFX1 gate213(.Q (g195), .QB (line213), .D(g30836), .CK(clk));
DFFX1 gate214(.Q (g198), .QB (line214), .D(g30837), .CK(clk));
DFFX1 gate215(.Q (g201), .QB (line215), .D(g30838), .CK(clk));
DFFX1 gate216(.Q (g240), .QB (line216), .D(g30845), .CK(clk));
DFFX1 gate217(.Q (g243), .QB (line217), .D(g30846), .CK(clk));
DFFX1 gate218(.Q (g246), .QB (line218), .D(g30847), .CK(clk));
DFFX1 gate219(.Q (g204), .QB (line219), .D(g30509), .CK(clk));
DFFX1 gate220(.Q (g207), .QB (line220), .D(g30510), .CK(clk));
DFFX1 gate221(.Q (g210), .QB (line221), .D(g30511), .CK(clk));
DFFX1 gate222(.Q (g249), .QB (line222), .D(g30515), .CK(clk));
DFFX1 gate223(.Q (g252), .QB (line223), .D(g30516), .CK(clk));
DFFX1 gate224(.Q (g255), .QB (line224), .D(g30517), .CK(clk));
DFFX1 gate225(.Q (g213), .QB (line225), .D(g30512), .CK(clk));
DFFX1 gate226(.Q (g216), .QB (line226), .D(g30513), .CK(clk));
DFFX1 gate227(.Q (g219), .QB (line227), .D(g30514), .CK(clk));
DFFX1 gate228(.Q (g258), .QB (line228), .D(g30518), .CK(clk));
DFFX1 gate229(.Q (g261), .QB (line229), .D(g30519), .CK(clk));
DFFX1 gate230(.Q (g264), .QB (line230), .D(g30520), .CK(clk));
DFFX1 gate231(.Q (g222), .QB (line231), .D(g30839), .CK(clk));
DFFX1 gate232(.Q (g225), .QB (line232), .D(g30840), .CK(clk));
DFFX1 gate233(.Q (g228), .QB (line233), .D(g30841), .CK(clk));
DFFX1 gate234(.Q (g267), .QB (line234), .D(g30848), .CK(clk));
DFFX1 gate235(.Q (g270), .QB (line235), .D(g30849), .CK(clk));
DFFX1 gate236(.Q (g273), .QB (line236), .D(g30850), .CK(clk));
DFFX1 gate237(.Q (g92), .QB (line237), .D(g25983), .CK(clk));
DFFX1 gate238(.Q (g88), .QB (line238), .D(g26678), .CK(clk));
DFFX1 gate239(.Q (g83), .QB (line239), .D(g27189), .CK(clk));
DFFX1 gate240(.Q (g79), .QB (line240), .D(g27683), .CK(clk));
DFFX1 gate241(.Q (g74), .QB (line241), .D(g28206), .CK(clk));
DFFX1 gate242(.Q (g70), .QB (line242), .D(g28673), .CK(clk));
DFFX1 gate243(.Q (g65), .QB (line243), .D(g29131), .CK(clk));
DFFX1 gate244(.Q (g61), .QB (line244), .D(g29413), .CK(clk));
DFFX1 gate245(.Q (g56), .QB (line245), .D(g29627), .CK(clk));
DFFX1 gate246(.Q (g52), .QB (line246), .D(g29794), .CK(clk));
DFFX1 gate247(.Q (g180), .QB (line247), .D(g20555), .CK(clk));
DFFX1 gate248(.Q (g182), .QB (line248), .D(g180), .CK(clk));
DFFX1 gate249(.Q (g181), .QB (line249), .D(g182), .CK(clk));
DFFX1 gate250(.Q (g276), .QB (line250), .D(g13406), .CK(clk));
DFFX1 gate251(.Q (g405), .QB (line251), .D(g276), .CK(clk));
DFFX1 gate252(.Q (g401), .QB (line252), .D(g405), .CK(clk));
DFFX1 gate253(.Q (g309), .QB (line253), .D(g11496), .CK(clk));
DFFX1 gate254(.Q (g354), .QB (line254), .D(g28207), .CK(clk));
DFFX1 gate255(.Q (g343), .QB (line255), .D(g28208), .CK(clk));
DFFX1 gate256(.Q (g346), .QB (line256), .D(g28209), .CK(clk));
DFFX1 gate257(.Q (g369), .QB (line257), .D(g28210), .CK(clk));
DFFX1 gate258(.Q (g358), .QB (line258), .D(g28211), .CK(clk));
DFFX1 gate259(.Q (g361), .QB (line259), .D(g28212), .CK(clk));
DFFX1 gate260(.Q (g384), .QB (line260), .D(g28213), .CK(clk));
DFFX1 gate261(.Q (g373), .QB (line261), .D(g28214), .CK(clk));
DFFX1 gate262(.Q (g376), .QB (line262), .D(g28215), .CK(clk));
DFFX1 gate263(.Q (g398), .QB (line263), .D(g28216), .CK(clk));
DFFX1 gate264(.Q (g388), .QB (line264), .D(g28217), .CK(clk));
DFFX1 gate265(.Q (g391), .QB (line265), .D(g28218), .CK(clk));
DFFX1 gate266(.Q (g408), .QB (line266), .D(g29414), .CK(clk));
DFFX1 gate267(.Q (g411), .QB (line267), .D(g29415), .CK(clk));
DFFX1 gate268(.Q (g414), .QB (line268), .D(g29416), .CK(clk));
DFFX1 gate269(.Q (g417), .QB (line269), .D(g29631), .CK(clk));
DFFX1 gate270(.Q (g420), .QB (line270), .D(g29632), .CK(clk));
DFFX1 gate271(.Q (g423), .QB (line271), .D(g29633), .CK(clk));
DFFX1 gate272(.Q (g427), .QB (line272), .D(g29417), .CK(clk));
DFFX1 gate273(.Q (g428), .QB (line273), .D(g29418), .CK(clk));
DFFX1 gate274(.Q (g426), .QB (line274), .D(g29419), .CK(clk));
DFFX1 gate275(.Q (g429), .QB (line275), .D(g27684), .CK(clk));
DFFX1 gate276(.Q (g432), .QB (line276), .D(g27685), .CK(clk));
DFFX1 gate277(.Q (g435), .QB (line277), .D(g27686), .CK(clk));
DFFX1 gate278(.Q (g438), .QB (line278), .D(g27687), .CK(clk));
DFFX1 gate279(.Q (g441), .QB (line279), .D(g27688), .CK(clk));
DFFX1 gate280(.Q (g444), .QB (line280), .D(g27689), .CK(clk));
DFFX1 gate281(.Q (g448), .QB (line281), .D(g28674), .CK(clk));
DFFX1 gate282(.Q (g449), .QB (line282), .D(g28675), .CK(clk));
DFFX1 gate283(.Q (g447), .QB (line283), .D(g28676), .CK(clk));
DFFX1 gate284(.Q (g312), .QB (line284), .D(g29795), .CK(clk));
DFFX1 gate285(.Q (g313), .QB (line285), .D(g29796), .CK(clk));
DFFX1 gate286(.Q (g314), .QB (line286), .D(g29797), .CK(clk));
DFFX1 gate287(.Q (g315), .QB (line287), .D(g30851), .CK(clk));
DFFX1 gate288(.Q (g316), .QB (line288), .D(g30852), .CK(clk));
DFFX1 gate289(.Q (g317), .QB (line289), .D(g30853), .CK(clk));
DFFX1 gate290(.Q (g318), .QB (line290), .D(g30710), .CK(clk));
DFFX1 gate291(.Q (g319), .QB (line291), .D(g30711), .CK(clk));
DFFX1 gate292(.Q (g320), .QB (line292), .D(g30712), .CK(clk));
DFFX1 gate293(.Q (g322), .QB (line293), .D(g29628), .CK(clk));
DFFX1 gate294(.Q (g323), .QB (line294), .D(g29629), .CK(clk));
DFFX1 gate295(.Q (g321), .QB (line295), .D(g29630), .CK(clk));
DFFX1 gate296(.Q (g403), .QB (line296), .D(g27191), .CK(clk));
DFFX1 gate297(.Q (g404), .QB (line297), .D(g27192), .CK(clk));
DFFX1 gate298(.Q (g402), .QB (line298), .D(g27193), .CK(clk));
DFFX1 gate299(.Q (g450), .QB (line299), .D(g11509), .CK(clk));
DFFX1 gate300(.Q (g451), .QB (line300), .D(g450), .CK(clk));
DFFX1 gate301(.Q (g452), .QB (line301), .D(g11510), .CK(clk));
DFFX1 gate302(.Q (g453), .QB (line302), .D(g452), .CK(clk));
DFFX1 gate303(.Q (g454), .QB (line303), .D(g11511), .CK(clk));
DFFX1 gate304(.Q (g279), .QB (line304), .D(g454), .CK(clk));
DFFX1 gate305(.Q (g280), .QB (line305), .D(g11491), .CK(clk));
DFFX1 gate306(.Q (g281), .QB (line306), .D(g280), .CK(clk));
DFFX1 gate307(.Q (g282), .QB (line307), .D(g11492), .CK(clk));
DFFX1 gate308(.Q (g283), .QB (line308), .D(g282), .CK(clk));
DFFX1 gate309(.Q (g284), .QB (line309), .D(g11493), .CK(clk));
DFFX1 gate310(.Q (g285), .QB (line310), .D(g284), .CK(clk));
DFFX1 gate311(.Q (g286), .QB (line311), .D(g11494), .CK(clk));
DFFX1 gate312(.Q (g287), .QB (line312), .D(g286), .CK(clk));
DFFX1 gate313(.Q (g288), .QB (line313), .D(g11495), .CK(clk));
DFFX1 gate314(.Q (g289), .QB (line314), .D(g288), .CK(clk));
DFFX1 gate315(.Q (g290), .QB (line315), .D(g13407), .CK(clk));
DFFX1 gate316(.Q (g291), .QB (line316), .D(g290), .CK(clk));
DFFX1 gate317(.Q (g299), .QB (line317), .D(g19012), .CK(clk));
DFFX1 gate318(.Q (g305), .QB (line318), .D(g23148), .CK(clk));
DFFX1 gate319(.Q (g308), .QB (line319), .D(g23149), .CK(clk));
DFFX1 gate320(.Q (g297), .QB (line320), .D(g23150), .CK(clk));
DFFX1 gate321(.Q (g296), .QB (line321), .D(g23151), .CK(clk));
DFFX1 gate322(.Q (g295), .QB (line322), .D(g23152), .CK(clk));
DFFX1 gate323(.Q (g294), .QB (line323), .D(g23153), .CK(clk));
DFFX1 gate324(.Q (g304), .QB (line324), .D(g19016), .CK(clk));
DFFX1 gate325(.Q (g303), .QB (line325), .D(g19015), .CK(clk));
DFFX1 gate326(.Q (g302), .QB (line326), .D(g19014), .CK(clk));
DFFX1 gate327(.Q (g301), .QB (line327), .D(g19013), .CK(clk));
DFFX1 gate328(.Q (g300), .QB (line328), .D(g25130), .CK(clk));
DFFX1 gate329(.Q (g298), .QB (line329), .D(g27190), .CK(clk));
DFFX1 gate330(.Q (g342), .QB (line330), .D(g11497), .CK(clk));
DFFX1 gate331(.Q (g349), .QB (line331), .D(g342), .CK(clk));
DFFX1 gate332(.Q (g350), .QB (line332), .D(g11498), .CK(clk));
DFFX1 gate333(.Q (g351), .QB (line333), .D(g350), .CK(clk));
DFFX1 gate334(.Q (g352), .QB (line334), .D(g11499), .CK(clk));
DFFX1 gate335(.Q (g353), .QB (line335), .D(g352), .CK(clk));
DFFX1 gate336(.Q (g357), .QB (line336), .D(g11500), .CK(clk));
DFFX1 gate337(.Q (g364), .QB (line337), .D(g357), .CK(clk));
DFFX1 gate338(.Q (g365), .QB (line338), .D(g11501), .CK(clk));
DFFX1 gate339(.Q (g366), .QB (line339), .D(g365), .CK(clk));
DFFX1 gate340(.Q (g367), .QB (line340), .D(g11502), .CK(clk));
DFFX1 gate341(.Q (g368), .QB (line341), .D(g367), .CK(clk));
DFFX1 gate342(.Q (g372), .QB (line342), .D(g11503), .CK(clk));
DFFX1 gate343(.Q (g379), .QB (line343), .D(g372), .CK(clk));
DFFX1 gate344(.Q (g380), .QB (line344), .D(g11504), .CK(clk));
DFFX1 gate345(.Q (g381), .QB (line345), .D(g380), .CK(clk));
DFFX1 gate346(.Q (g382), .QB (line346), .D(g11505), .CK(clk));
DFFX1 gate347(.Q (g383), .QB (line347), .D(g382), .CK(clk));
DFFX1 gate348(.Q (g387), .QB (line348), .D(g11506), .CK(clk));
DFFX1 gate349(.Q (g394), .QB (line349), .D(g387), .CK(clk));
DFFX1 gate350(.Q (g395), .QB (line350), .D(g11507), .CK(clk));
DFFX1 gate351(.Q (g396), .QB (line351), .D(g395), .CK(clk));
DFFX1 gate352(.Q (g397), .QB (line352), .D(g11508), .CK(clk));
DFFX1 gate353(.Q (g324), .QB (line353), .D(g397), .CK(clk));
DFFX1 gate354(.Q (g325), .QB (line354), .D(g13408), .CK(clk));
DFFX1 gate355(.Q (g331), .QB (line355), .D(g325), .CK(clk));
DFFX1 gate356(.Q (g337), .QB (line356), .D(g331), .CK(clk));
DFFX1 gate357(.Q (g545), .QB (line357), .D(g13419), .CK(clk));
DFFX1 gate358(.Q (g551), .QB (line358), .D(g545), .CK(clk));
DFFX1 gate359(.Q (g550), .QB (line359), .D(g551), .CK(clk));
DFFX1 gate360(.Q (g554), .QB (line360), .D(g23160), .CK(clk));
DFFX1 gate361(.Q (g557), .QB (line361), .D(g20556), .CK(clk));
DFFX1 gate362(.Q (g510), .QB (line362), .D(g20557), .CK(clk));
DFFX1 gate363(.Q (g513), .QB (line363), .D(g16467), .CK(clk));
DFFX1 gate364(.Q (g523), .QB (line364), .D(g513), .CK(clk));
DFFX1 gate365(.Q (g524), .QB (line365), .D(g523), .CK(clk));
DFFX1 gate366(.Q (g564), .QB (line366), .D(g11512), .CK(clk));
DFFX1 gate367(.Q (g569), .QB (line367), .D(g564), .CK(clk));
DFFX1 gate368(.Q (g570), .QB (line368), .D(g11515), .CK(clk));
DFFX1 gate369(.Q (g571), .QB (line369), .D(g570), .CK(clk));
DFFX1 gate370(.Q (g572), .QB (line370), .D(g11516), .CK(clk));
DFFX1 gate371(.Q (g573), .QB (line371), .D(g572), .CK(clk));
DFFX1 gate372(.Q (g574), .QB (line372), .D(g11517), .CK(clk));
DFFX1 gate373(.Q (g565), .QB (line373), .D(g574), .CK(clk));
DFFX1 gate374(.Q (g566), .QB (line374), .D(g11513), .CK(clk));
DFFX1 gate375(.Q (g567), .QB (line375), .D(g566), .CK(clk));
DFFX1 gate376(.Q (g568), .QB (line376), .D(g11514), .CK(clk));
DFFX1 gate377(.Q (g489), .QB (line377), .D(g568), .CK(clk));
DFFX1 gate378(.Q (g474), .QB (line378), .D(g13409), .CK(clk));
DFFX1 gate379(.Q (g481), .QB (line379), .D(g474), .CK(clk));
DFFX1 gate380(.Q (g485), .QB (line380), .D(g481), .CK(clk));
DFFX1 gate381(.Q (g486), .QB (line381), .D(g24292), .CK(clk));
DFFX1 gate382(.Q (g487), .QB (line382), .D(g24293), .CK(clk));
DFFX1 gate383(.Q (g488), .QB (line383), .D(g24294), .CK(clk));
DFFX1 gate384(.Q (g455), .QB (line384), .D(g25139), .CK(clk));
DFFX1 gate385(.Q (g458), .QB (line385), .D(g25131), .CK(clk));
DFFX1 gate386(.Q (g461), .QB (line386), .D(g25132), .CK(clk));
DFFX1 gate387(.Q (g477), .QB (line387), .D(g25136), .CK(clk));
DFFX1 gate388(.Q (g478), .QB (line388), .D(g25137), .CK(clk));
DFFX1 gate389(.Q (g479), .QB (line389), .D(g25138), .CK(clk));
DFFX1 gate390(.Q (g480), .QB (line390), .D(g24289), .CK(clk));
DFFX1 gate391(.Q (g484), .QB (line391), .D(g24290), .CK(clk));
DFFX1 gate392(.Q (g464), .QB (line392), .D(g24291), .CK(clk));
DFFX1 gate393(.Q (g465), .QB (line393), .D(g25133), .CK(clk));
DFFX1 gate394(.Q (g468), .QB (line394), .D(g25134), .CK(clk));
DFFX1 gate395(.Q (g471), .QB (line395), .D(g25135), .CK(clk));
DFFX1 gate396(.Q (g528), .QB (line396), .D(g16468), .CK(clk));
DFFX1 gate397(.Q (g535), .QB (line397), .D(g528), .CK(clk));
DFFX1 gate398(.Q (g542), .QB (line398), .D(g535), .CK(clk));
DFFX1 gate399(.Q (g543), .QB (line399), .D(g19021), .CK(clk));
DFFX1 gate400(.Q (g544), .QB (line400), .D(g543), .CK(clk));
DFFX1 gate401(.Q (g548), .QB (line401), .D(g23159), .CK(clk));
DFFX1 gate402(.Q (g549), .QB (line402), .D(g19022), .CK(clk));
DFFX1 gate403(.Q (g499), .QB (line403), .D(g549), .CK(clk));
DFFX1 gate404(.Q (g558), .QB (line404), .D(g19023), .CK(clk));
DFFX1 gate405(.Q (g559), .QB (line405), .D(g558), .CK(clk));
DFFX1 gate406(.Q (g576), .QB (line406), .D(g28219), .CK(clk));
DFFX1 gate407(.Q (g577), .QB (line407), .D(g28220), .CK(clk));
DFFX1 gate408(.Q (g575), .QB (line408), .D(g28221), .CK(clk));
DFFX1 gate409(.Q (g579), .QB (line409), .D(g28222), .CK(clk));
DFFX1 gate410(.Q (g580), .QB (line410), .D(g28223), .CK(clk));
DFFX1 gate411(.Q (g578), .QB (line411), .D(g28224), .CK(clk));
DFFX1 gate412(.Q (g582), .QB (line412), .D(g28225), .CK(clk));
DFFX1 gate413(.Q (g583), .QB (line413), .D(g28226), .CK(clk));
DFFX1 gate414(.Q (g581), .QB (line414), .D(g28227), .CK(clk));
DFFX1 gate415(.Q (g585), .QB (line415), .D(g28228), .CK(clk));
DFFX1 gate416(.Q (g586), .QB (line416), .D(g28229), .CK(clk));
DFFX1 gate417(.Q (g584), .QB (line417), .D(g28230), .CK(clk));
DFFX1 gate418(.Q (g587), .QB (line418), .D(g25985), .CK(clk));
DFFX1 gate419(.Q (g590), .QB (line419), .D(g25986), .CK(clk));
DFFX1 gate420(.Q (g593), .QB (line420), .D(g25987), .CK(clk));
DFFX1 gate421(.Q (g596), .QB (line421), .D(g25988), .CK(clk));
DFFX1 gate422(.Q (g599), .QB (line422), .D(g25989), .CK(clk));
DFFX1 gate423(.Q (g602), .QB (line423), .D(g25990), .CK(clk));
DFFX1 gate424(.Q (g614), .QB (line424), .D(g29135), .CK(clk));
DFFX1 gate425(.Q (g617), .QB (line425), .D(g29136), .CK(clk));
DFFX1 gate426(.Q (g620), .QB (line426), .D(g29137), .CK(clk));
DFFX1 gate427(.Q (g605), .QB (line427), .D(g29132), .CK(clk));
DFFX1 gate428(.Q (g608), .QB (line428), .D(g29133), .CK(clk));
DFFX1 gate429(.Q (g611), .QB (line429), .D(g29134), .CK(clk));
DFFX1 gate430(.Q (g490), .QB (line430), .D(g27194), .CK(clk));
DFFX1 gate431(.Q (g493), .QB (line431), .D(g27195), .CK(clk));
DFFX1 gate432(.Q (g496), .QB (line432), .D(g27196), .CK(clk));
DFFX1 gate433(.Q (g506), .QB (line433), .D(g8284), .CK(clk));
DFFX1 gate434(.Q (g507), .QB (line434), .D(g24295), .CK(clk));
DFFX1 gate435(.Q (g508), .QB (line435), .D(g19017), .CK(clk));
DFFX1 gate436(.Q (g509), .QB (line436), .D(g19018), .CK(clk));
DFFX1 gate437(.Q (g514), .QB (line437), .D(g19019), .CK(clk));
DFFX1 gate438(.Q (g515), .QB (line438), .D(g19020), .CK(clk));
DFFX1 gate439(.Q (g516), .QB (line439), .D(g23158), .CK(clk));
DFFX1 gate440(.Q (g517), .QB (line440), .D(g23157), .CK(clk));
DFFX1 gate441(.Q (g518), .QB (line441), .D(g23156), .CK(clk));
DFFX1 gate442(.Q (g519), .QB (line442), .D(g23155), .CK(clk));
DFFX1 gate443(.Q (g520), .QB (line443), .D(g23154), .CK(clk));
DFFX1 gate444(.Q (g525), .QB (line444), .D(g520), .CK(clk));
DFFX1 gate445(.Q (g529), .QB (line445), .D(g13410), .CK(clk));
DFFX1 gate446(.Q (g530), .QB (line446), .D(g13411), .CK(clk));
DFFX1 gate447(.Q (g531), .QB (line447), .D(g13412), .CK(clk));
DFFX1 gate448(.Q (g532), .QB (line448), .D(g13413), .CK(clk));
DFFX1 gate449(.Q (g533), .QB (line449), .D(g13414), .CK(clk));
DFFX1 gate450(.Q (g534), .QB (line450), .D(g13415), .CK(clk));
DFFX1 gate451(.Q (g536), .QB (line451), .D(g13416), .CK(clk));
DFFX1 gate452(.Q (g537), .QB (line452), .D(g13417), .CK(clk));
DFFX1 gate453(.Q (g538), .QB (line453), .D(g25984), .CK(clk));
DFFX1 gate454(.Q (g541), .QB (line454), .D(g13418), .CK(clk));
DFFX1 gate455(.Q (g623), .QB (line455), .D(g13420), .CK(clk));
DFFX1 gate456(.Q (g626), .QB (line456), .D(g623), .CK(clk));
DFFX1 gate457(.Q (g629), .QB (line457), .D(g626), .CK(clk));
DFFX1 gate458(.Q (g630), .QB (line458), .D(g20558), .CK(clk));
DFFX1 gate459(.Q (g659), .QB (line459), .D(g21943), .CK(clk));
DFFX1 gate460(.Q (g640), .QB (line460), .D(g23161), .CK(clk));
DFFX1 gate461(.Q (g633), .QB (line461), .D(g24296), .CK(clk));
DFFX1 gate462(.Q (g653), .QB (line462), .D(g25140), .CK(clk));
DFFX1 gate463(.Q (g646), .QB (line463), .D(g25991), .CK(clk));
DFFX1 gate464(.Q (g660), .QB (line464), .D(g26691), .CK(clk));
DFFX1 gate465(.Q (g672), .QB (line465), .D(g27197), .CK(clk));
DFFX1 gate466(.Q (g666), .QB (line466), .D(g27690), .CK(clk));
DFFX1 gate467(.Q (g679), .QB (line467), .D(g28231), .CK(clk));
DFFX1 gate468(.Q (g686), .QB (line468), .D(g28677), .CK(clk));
DFFX1 gate469(.Q (g692), .QB (line469), .D(g29138), .CK(clk));
DFFX1 gate470(.Q (g699), .QB (line470), .D(g23162), .CK(clk));
DFFX1 gate471(.Q (g700), .QB (line471), .D(g23163), .CK(clk));
DFFX1 gate472(.Q (g698), .QB (line472), .D(g23164), .CK(clk));
DFFX1 gate473(.Q (g702), .QB (line473), .D(g23165), .CK(clk));
DFFX1 gate474(.Q (g703), .QB (line474), .D(g23166), .CK(clk));
DFFX1 gate475(.Q (g701), .QB (line475), .D(g23167), .CK(clk));
DFFX1 gate476(.Q (g705), .QB (line476), .D(g23168), .CK(clk));
DFFX1 gate477(.Q (g706), .QB (line477), .D(g23169), .CK(clk));
DFFX1 gate478(.Q (g704), .QB (line478), .D(g23170), .CK(clk));
DFFX1 gate479(.Q (g708), .QB (line479), .D(g23171), .CK(clk));
DFFX1 gate480(.Q (g709), .QB (line480), .D(g23172), .CK(clk));
DFFX1 gate481(.Q (g707), .QB (line481), .D(g23173), .CK(clk));
DFFX1 gate482(.Q (g711), .QB (line482), .D(g23174), .CK(clk));
DFFX1 gate483(.Q (g712), .QB (line483), .D(g23175), .CK(clk));
DFFX1 gate484(.Q (g710), .QB (line484), .D(g23176), .CK(clk));
DFFX1 gate485(.Q (g714), .QB (line485), .D(g23177), .CK(clk));
DFFX1 gate486(.Q (g715), .QB (line486), .D(g23178), .CK(clk));
DFFX1 gate487(.Q (g713), .QB (line487), .D(g23179), .CK(clk));
DFFX1 gate488(.Q (g717), .QB (line488), .D(g23180), .CK(clk));
DFFX1 gate489(.Q (g718), .QB (line489), .D(g23181), .CK(clk));
DFFX1 gate490(.Q (g716), .QB (line490), .D(g23182), .CK(clk));
DFFX1 gate491(.Q (g720), .QB (line491), .D(g23183), .CK(clk));
DFFX1 gate492(.Q (g721), .QB (line492), .D(g23184), .CK(clk));
DFFX1 gate493(.Q (g719), .QB (line493), .D(g23185), .CK(clk));
DFFX1 gate494(.Q (g723), .QB (line494), .D(g23186), .CK(clk));
DFFX1 gate495(.Q (g724), .QB (line495), .D(g23187), .CK(clk));
DFFX1 gate496(.Q (g722), .QB (line496), .D(g23188), .CK(clk));
DFFX1 gate497(.Q (g726), .QB (line497), .D(g23189), .CK(clk));
DFFX1 gate498(.Q (g727), .QB (line498), .D(g23190), .CK(clk));
DFFX1 gate499(.Q (g725), .QB (line499), .D(g23191), .CK(clk));
DFFX1 gate500(.Q (g729), .QB (line500), .D(g23192), .CK(clk));
DFFX1 gate501(.Q (g730), .QB (line501), .D(g23193), .CK(clk));
DFFX1 gate502(.Q (g728), .QB (line502), .D(g23194), .CK(clk));
DFFX1 gate503(.Q (g732), .QB (line503), .D(g23195), .CK(clk));
DFFX1 gate504(.Q (g733), .QB (line504), .D(g23196), .CK(clk));
DFFX1 gate505(.Q (g731), .QB (line505), .D(g23197), .CK(clk));
DFFX1 gate506(.Q (g735), .QB (line506), .D(g26692), .CK(clk));
DFFX1 gate507(.Q (g736), .QB (line507), .D(g26693), .CK(clk));
DFFX1 gate508(.Q (g734), .QB (line508), .D(g26694), .CK(clk));
DFFX1 gate509(.Q (g738), .QB (line509), .D(g24297), .CK(clk));
DFFX1 gate510(.Q (g739), .QB (line510), .D(g24298), .CK(clk));
DFFX1 gate511(.Q (g737), .QB (line511), .D(g24299), .CK(clk));
DFFX1 gate512(.Q (g826), .QB (line512), .D(g13421), .CK(clk));
DFFX1 gate513(.Q (g823), .QB (line513), .D(g826), .CK(clk));
DFFX1 gate514(.Q (g853), .QB (line514), .D(g823), .CK(clk));
DFFX1 gate515(.Q (g818), .QB (line515), .D(g24300), .CK(clk));
DFFX1 gate516(.Q (g819), .QB (line516), .D(g24301), .CK(clk));
DFFX1 gate517(.Q (g817), .QB (line517), .D(g24302), .CK(clk));
DFFX1 gate518(.Q (g821), .QB (line518), .D(g24303), .CK(clk));
DFFX1 gate519(.Q (g822), .QB (line519), .D(g24304), .CK(clk));
DFFX1 gate520(.Q (g820), .QB (line520), .D(g24305), .CK(clk));
DFFX1 gate521(.Q (g830), .QB (line521), .D(g24306), .CK(clk));
DFFX1 gate522(.Q (g831), .QB (line522), .D(g24307), .CK(clk));
DFFX1 gate523(.Q (g829), .QB (line523), .D(g24308), .CK(clk));
DFFX1 gate524(.Q (g833), .QB (line524), .D(g24309), .CK(clk));
DFFX1 gate525(.Q (g834), .QB (line525), .D(g24310), .CK(clk));
DFFX1 gate526(.Q (g832), .QB (line526), .D(g24311), .CK(clk));
DFFX1 gate527(.Q (g836), .QB (line527), .D(g24312), .CK(clk));
DFFX1 gate528(.Q (g837), .QB (line528), .D(g24313), .CK(clk));
DFFX1 gate529(.Q (g835), .QB (line529), .D(g24314), .CK(clk));
DFFX1 gate530(.Q (g839), .QB (line530), .D(g24315), .CK(clk));
DFFX1 gate531(.Q (g840), .QB (line531), .D(g24316), .CK(clk));
DFFX1 gate532(.Q (g838), .QB (line532), .D(g24317), .CK(clk));
DFFX1 gate533(.Q (g842), .QB (line533), .D(g24318), .CK(clk));
DFFX1 gate534(.Q (g843), .QB (line534), .D(g24319), .CK(clk));
DFFX1 gate535(.Q (g841), .QB (line535), .D(g24320), .CK(clk));
DFFX1 gate536(.Q (g845), .QB (line536), .D(g24321), .CK(clk));
DFFX1 gate537(.Q (g846), .QB (line537), .D(g24322), .CK(clk));
DFFX1 gate538(.Q (g844), .QB (line538), .D(g24323), .CK(clk));
DFFX1 gate539(.Q (g848), .QB (line539), .D(g24324), .CK(clk));
DFFX1 gate540(.Q (g849), .QB (line540), .D(g24325), .CK(clk));
DFFX1 gate541(.Q (g847), .QB (line541), .D(g24326), .CK(clk));
DFFX1 gate542(.Q (g851), .QB (line542), .D(g24327), .CK(clk));
DFFX1 gate543(.Q (g852), .QB (line543), .D(g24328), .CK(clk));
DFFX1 gate544(.Q (g850), .QB (line544), .D(g24329), .CK(clk));
DFFX1 gate545(.Q (g857), .QB (line545), .D(g26696), .CK(clk));
DFFX1 gate546(.Q (g858), .QB (line546), .D(g26697), .CK(clk));
DFFX1 gate547(.Q (g856), .QB (line547), .D(g26698), .CK(clk));
DFFX1 gate548(.Q (g860), .QB (line548), .D(g26699), .CK(clk));
DFFX1 gate549(.Q (g861), .QB (line549), .D(g26700), .CK(clk));
DFFX1 gate550(.Q (g859), .QB (line550), .D(g26701), .CK(clk));
DFFX1 gate551(.Q (g863), .QB (line551), .D(g26702), .CK(clk));
DFFX1 gate552(.Q (g864), .QB (line552), .D(g26703), .CK(clk));
DFFX1 gate553(.Q (g862), .QB (line553), .D(g26704), .CK(clk));
DFFX1 gate554(.Q (g866), .QB (line554), .D(g26705), .CK(clk));
DFFX1 gate555(.Q (g867), .QB (line555), .D(g26706), .CK(clk));
DFFX1 gate556(.Q (g865), .QB (line556), .D(g26707), .CK(clk));
DFFX1 gate557(.Q (g873), .QB (line557), .D(g30521), .CK(clk));
DFFX1 gate558(.Q (g876), .QB (line558), .D(g30522), .CK(clk));
DFFX1 gate559(.Q (g879), .QB (line559), .D(g30523), .CK(clk));
DFFX1 gate560(.Q (g918), .QB (line560), .D(g30860), .CK(clk));
DFFX1 gate561(.Q (g921), .QB (line561), .D(g30861), .CK(clk));
DFFX1 gate562(.Q (g924), .QB (line562), .D(g30862), .CK(clk));
DFFX1 gate563(.Q (g882), .QB (line563), .D(g30854), .CK(clk));
DFFX1 gate564(.Q (g885), .QB (line564), .D(g30855), .CK(clk));
DFFX1 gate565(.Q (g888), .QB (line565), .D(g30856), .CK(clk));
DFFX1 gate566(.Q (g927), .QB (line566), .D(g30863), .CK(clk));
DFFX1 gate567(.Q (g930), .QB (line567), .D(g30864), .CK(clk));
DFFX1 gate568(.Q (g933), .QB (line568), .D(g30865), .CK(clk));
DFFX1 gate569(.Q (g891), .QB (line569), .D(g30524), .CK(clk));
DFFX1 gate570(.Q (g894), .QB (line570), .D(g30525), .CK(clk));
DFFX1 gate571(.Q (g897), .QB (line571), .D(g30526), .CK(clk));
DFFX1 gate572(.Q (g936), .QB (line572), .D(g30530), .CK(clk));
DFFX1 gate573(.Q (g939), .QB (line573), .D(g30531), .CK(clk));
DFFX1 gate574(.Q (g942), .QB (line574), .D(g30532), .CK(clk));
DFFX1 gate575(.Q (g900), .QB (line575), .D(g30527), .CK(clk));
DFFX1 gate576(.Q (g903), .QB (line576), .D(g30528), .CK(clk));
DFFX1 gate577(.Q (g906), .QB (line577), .D(g30529), .CK(clk));
DFFX1 gate578(.Q (g945), .QB (line578), .D(g30533), .CK(clk));
DFFX1 gate579(.Q (g948), .QB (line579), .D(g30534), .CK(clk));
DFFX1 gate580(.Q (g951), .QB (line580), .D(g30535), .CK(clk));
DFFX1 gate581(.Q (g909), .QB (line581), .D(g30857), .CK(clk));
DFFX1 gate582(.Q (g912), .QB (line582), .D(g30858), .CK(clk));
DFFX1 gate583(.Q (g915), .QB (line583), .D(g30859), .CK(clk));
DFFX1 gate584(.Q (g954), .QB (line584), .D(g30866), .CK(clk));
DFFX1 gate585(.Q (g957), .QB (line585), .D(g30867), .CK(clk));
DFFX1 gate586(.Q (g960), .QB (line586), .D(g30868), .CK(clk));
DFFX1 gate587(.Q (g780), .QB (line587), .D(g25992), .CK(clk));
DFFX1 gate588(.Q (g776), .QB (line588), .D(g26695), .CK(clk));
DFFX1 gate589(.Q (g771), .QB (line589), .D(g27198), .CK(clk));
DFFX1 gate590(.Q (g767), .QB (line590), .D(g27691), .CK(clk));
DFFX1 gate591(.Q (g762), .QB (line591), .D(g28232), .CK(clk));
DFFX1 gate592(.Q (g758), .QB (line592), .D(g28678), .CK(clk));
DFFX1 gate593(.Q (g753), .QB (line593), .D(g29139), .CK(clk));
DFFX1 gate594(.Q (g749), .QB (line594), .D(g29420), .CK(clk));
DFFX1 gate595(.Q (g744), .QB (line595), .D(g29634), .CK(clk));
DFFX1 gate596(.Q (g740), .QB (line596), .D(g29798), .CK(clk));
DFFX1 gate597(.Q (g868), .QB (line597), .D(g20559), .CK(clk));
DFFX1 gate598(.Q (g870), .QB (line598), .D(g868), .CK(clk));
DFFX1 gate599(.Q (g869), .QB (line599), .D(g870), .CK(clk));
DFFX1 gate600(.Q (g963), .QB (line600), .D(g13422), .CK(clk));
DFFX1 gate601(.Q (g1092), .QB (line601), .D(g963), .CK(clk));
DFFX1 gate602(.Q (g1088), .QB (line602), .D(g1092), .CK(clk));
DFFX1 gate603(.Q (g996), .QB (line603), .D(g11523), .CK(clk));
DFFX1 gate604(.Q (g1041), .QB (line604), .D(g28233), .CK(clk));
DFFX1 gate605(.Q (g1030), .QB (line605), .D(g28234), .CK(clk));
DFFX1 gate606(.Q (g1033), .QB (line606), .D(g28235), .CK(clk));
DFFX1 gate607(.Q (g1056), .QB (line607), .D(g28236), .CK(clk));
DFFX1 gate608(.Q (g1045), .QB (line608), .D(g28237), .CK(clk));
DFFX1 gate609(.Q (g1048), .QB (line609), .D(g28238), .CK(clk));
DFFX1 gate610(.Q (g1071), .QB (line610), .D(g28239), .CK(clk));
DFFX1 gate611(.Q (g1060), .QB (line611), .D(g28240), .CK(clk));
DFFX1 gate612(.Q (g1063), .QB (line612), .D(g28241), .CK(clk));
DFFX1 gate613(.Q (g1085), .QB (line613), .D(g28242), .CK(clk));
DFFX1 gate614(.Q (g1075), .QB (line614), .D(g28243), .CK(clk));
DFFX1 gate615(.Q (g1078), .QB (line615), .D(g28244), .CK(clk));
DFFX1 gate616(.Q (g1095), .QB (line616), .D(g29421), .CK(clk));
DFFX1 gate617(.Q (g1098), .QB (line617), .D(g29422), .CK(clk));
DFFX1 gate618(.Q (g1101), .QB (line618), .D(g29423), .CK(clk));
DFFX1 gate619(.Q (g1104), .QB (line619), .D(g29638), .CK(clk));
DFFX1 gate620(.Q (g1107), .QB (line620), .D(g29639), .CK(clk));
DFFX1 gate621(.Q (g1110), .QB (line621), .D(g29640), .CK(clk));
DFFX1 gate622(.Q (g1114), .QB (line622), .D(g29424), .CK(clk));
DFFX1 gate623(.Q (g1115), .QB (line623), .D(g29425), .CK(clk));
DFFX1 gate624(.Q (g1113), .QB (line624), .D(g29426), .CK(clk));
DFFX1 gate625(.Q (g1116), .QB (line625), .D(g27692), .CK(clk));
DFFX1 gate626(.Q (g1119), .QB (line626), .D(g27693), .CK(clk));
DFFX1 gate627(.Q (g1122), .QB (line627), .D(g27694), .CK(clk));
DFFX1 gate628(.Q (g1125), .QB (line628), .D(g27695), .CK(clk));
DFFX1 gate629(.Q (g1128), .QB (line629), .D(g27696), .CK(clk));
DFFX1 gate630(.Q (g1131), .QB (line630), .D(g27697), .CK(clk));
DFFX1 gate631(.Q (g1135), .QB (line631), .D(g28679), .CK(clk));
DFFX1 gate632(.Q (g1136), .QB (line632), .D(g28680), .CK(clk));
DFFX1 gate633(.Q (g1134), .QB (line633), .D(g28681), .CK(clk));
DFFX1 gate634(.Q (g999), .QB (line634), .D(g29799), .CK(clk));
DFFX1 gate635(.Q (g1000), .QB (line635), .D(g29800), .CK(clk));
DFFX1 gate636(.Q (g1001), .QB (line636), .D(g29801), .CK(clk));
DFFX1 gate637(.Q (g1002), .QB (line637), .D(g30869), .CK(clk));
DFFX1 gate638(.Q (g1003), .QB (line638), .D(g30870), .CK(clk));
DFFX1 gate639(.Q (g1004), .QB (line639), .D(g30871), .CK(clk));
DFFX1 gate640(.Q (g1005), .QB (line640), .D(g30713), .CK(clk));
DFFX1 gate641(.Q (g1006), .QB (line641), .D(g30714), .CK(clk));
DFFX1 gate642(.Q (g1007), .QB (line642), .D(g30715), .CK(clk));
DFFX1 gate643(.Q (g1009), .QB (line643), .D(g29635), .CK(clk));
DFFX1 gate644(.Q (g1010), .QB (line644), .D(g29636), .CK(clk));
DFFX1 gate645(.Q (g1008), .QB (line645), .D(g29637), .CK(clk));
DFFX1 gate646(.Q (g1090), .QB (line646), .D(g27206), .CK(clk));
DFFX1 gate647(.Q (g1091), .QB (line647), .D(g27207), .CK(clk));
DFFX1 gate648(.Q (g1089), .QB (line648), .D(g27208), .CK(clk));
DFFX1 gate649(.Q (g1137), .QB (line649), .D(g11536), .CK(clk));
DFFX1 gate650(.Q (g1138), .QB (line650), .D(g1137), .CK(clk));
DFFX1 gate651(.Q (g1139), .QB (line651), .D(g11537), .CK(clk));
DFFX1 gate652(.Q (g1140), .QB (line652), .D(g1139), .CK(clk));
DFFX1 gate653(.Q (g1141), .QB (line653), .D(g11538), .CK(clk));
DFFX1 gate654(.Q (g966), .QB (line654), .D(g1141), .CK(clk));
DFFX1 gate655(.Q (g967), .QB (line655), .D(g11518), .CK(clk));
DFFX1 gate656(.Q (g968), .QB (line656), .D(g967), .CK(clk));
DFFX1 gate657(.Q (g969), .QB (line657), .D(g11519), .CK(clk));
DFFX1 gate658(.Q (g970), .QB (line658), .D(g969), .CK(clk));
DFFX1 gate659(.Q (g971), .QB (line659), .D(g11520), .CK(clk));
DFFX1 gate660(.Q (g972), .QB (line660), .D(g971), .CK(clk));
DFFX1 gate661(.Q (g973), .QB (line661), .D(g11521), .CK(clk));
DFFX1 gate662(.Q (g974), .QB (line662), .D(g973), .CK(clk));
DFFX1 gate663(.Q (g975), .QB (line663), .D(g11522), .CK(clk));
DFFX1 gate664(.Q (g976), .QB (line664), .D(g975), .CK(clk));
DFFX1 gate665(.Q (g977), .QB (line665), .D(g13423), .CK(clk));
DFFX1 gate666(.Q (g978), .QB (line666), .D(g977), .CK(clk));
DFFX1 gate667(.Q (g986), .QB (line667), .D(g19024), .CK(clk));
DFFX1 gate668(.Q (g992), .QB (line668), .D(g27200), .CK(clk));
DFFX1 gate669(.Q (g995), .QB (line669), .D(g27201), .CK(clk));
DFFX1 gate670(.Q (g984), .QB (line670), .D(g27202), .CK(clk));
DFFX1 gate671(.Q (g983), .QB (line671), .D(g27203), .CK(clk));
DFFX1 gate672(.Q (g982), .QB (line672), .D(g27204), .CK(clk));
DFFX1 gate673(.Q (g981), .QB (line673), .D(g27205), .CK(clk));
DFFX1 gate674(.Q (g991), .QB (line674), .D(g19028), .CK(clk));
DFFX1 gate675(.Q (g990), .QB (line675), .D(g19027), .CK(clk));
DFFX1 gate676(.Q (g989), .QB (line676), .D(g19026), .CK(clk));
DFFX1 gate677(.Q (g988), .QB (line677), .D(g19025), .CK(clk));
DFFX1 gate678(.Q (g987), .QB (line678), .D(g25141), .CK(clk));
DFFX1 gate679(.Q (g985), .QB (line679), .D(g27199), .CK(clk));
DFFX1 gate680(.Q (g1029), .QB (line680), .D(g11524), .CK(clk));
DFFX1 gate681(.Q (g1036), .QB (line681), .D(g1029), .CK(clk));
DFFX1 gate682(.Q (g1037), .QB (line682), .D(g11525), .CK(clk));
DFFX1 gate683(.Q (g1038), .QB (line683), .D(g1037), .CK(clk));
DFFX1 gate684(.Q (g1039), .QB (line684), .D(g11526), .CK(clk));
DFFX1 gate685(.Q (g1040), .QB (line685), .D(g1039), .CK(clk));
DFFX1 gate686(.Q (g1044), .QB (line686), .D(g11527), .CK(clk));
DFFX1 gate687(.Q (g1051), .QB (line687), .D(g1044), .CK(clk));
DFFX1 gate688(.Q (g1052), .QB (line688), .D(g11528), .CK(clk));
DFFX1 gate689(.Q (g1053), .QB (line689), .D(g1052), .CK(clk));
DFFX1 gate690(.Q (g1054), .QB (line690), .D(g11529), .CK(clk));
DFFX1 gate691(.Q (g1055), .QB (line691), .D(g1054), .CK(clk));
DFFX1 gate692(.Q (g1059), .QB (line692), .D(g11530), .CK(clk));
DFFX1 gate693(.Q (g1066), .QB (line693), .D(g1059), .CK(clk));
DFFX1 gate694(.Q (g1067), .QB (line694), .D(g11531), .CK(clk));
DFFX1 gate695(.Q (g1068), .QB (line695), .D(g1067), .CK(clk));
DFFX1 gate696(.Q (g1069), .QB (line696), .D(g11532), .CK(clk));
DFFX1 gate697(.Q (g1070), .QB (line697), .D(g1069), .CK(clk));
DFFX1 gate698(.Q (g1074), .QB (line698), .D(g11533), .CK(clk));
DFFX1 gate699(.Q (g1081), .QB (line699), .D(g1074), .CK(clk));
DFFX1 gate700(.Q (g1082), .QB (line700), .D(g11534), .CK(clk));
DFFX1 gate701(.Q (g1083), .QB (line701), .D(g1082), .CK(clk));
DFFX1 gate702(.Q (g1084), .QB (line702), .D(g11535), .CK(clk));
DFFX1 gate703(.Q (g1011), .QB (line703), .D(g1084), .CK(clk));
DFFX1 gate704(.Q (g1012), .QB (line704), .D(g13424), .CK(clk));
DFFX1 gate705(.Q (g1018), .QB (line705), .D(g1012), .CK(clk));
DFFX1 gate706(.Q (g1024), .QB (line706), .D(g1018), .CK(clk));
DFFX1 gate707(.Q (g1231), .QB (line707), .D(g13435), .CK(clk));
DFFX1 gate708(.Q (g1237), .QB (line708), .D(g1231), .CK(clk));
DFFX1 gate709(.Q (g1236), .QB (line709), .D(g1237), .CK(clk));
DFFX1 gate710(.Q (g1240), .QB (line710), .D(g23198), .CK(clk));
DFFX1 gate711(.Q (g1243), .QB (line711), .D(g20560), .CK(clk));
DFFX1 gate712(.Q (g1196), .QB (line712), .D(g20561), .CK(clk));
DFFX1 gate713(.Q (g1199), .QB (line713), .D(g16469), .CK(clk));
DFFX1 gate714(.Q (g1209), .QB (line714), .D(g1199), .CK(clk));
DFFX1 gate715(.Q (g1210), .QB (line715), .D(g1209), .CK(clk));
DFFX1 gate716(.Q (g1250), .QB (line716), .D(g11539), .CK(clk));
DFFX1 gate717(.Q (g1255), .QB (line717), .D(g1250), .CK(clk));
DFFX1 gate718(.Q (g1256), .QB (line718), .D(g11542), .CK(clk));
DFFX1 gate719(.Q (g1257), .QB (line719), .D(g1256), .CK(clk));
DFFX1 gate720(.Q (g1258), .QB (line720), .D(g11543), .CK(clk));
DFFX1 gate721(.Q (g1259), .QB (line721), .D(g1258), .CK(clk));
DFFX1 gate722(.Q (g1260), .QB (line722), .D(g11544), .CK(clk));
DFFX1 gate723(.Q (g1251), .QB (line723), .D(g1260), .CK(clk));
DFFX1 gate724(.Q (g1252), .QB (line724), .D(g11540), .CK(clk));
DFFX1 gate725(.Q (g1253), .QB (line725), .D(g1252), .CK(clk));
DFFX1 gate726(.Q (g1254), .QB (line726), .D(g11541), .CK(clk));
DFFX1 gate727(.Q (g1176), .QB (line727), .D(g1254), .CK(clk));
DFFX1 gate728(.Q (g1161), .QB (line728), .D(g13425), .CK(clk));
DFFX1 gate729(.Q (g1168), .QB (line729), .D(g1161), .CK(clk));
DFFX1 gate730(.Q (g1172), .QB (line730), .D(g1168), .CK(clk));
DFFX1 gate731(.Q (g1173), .QB (line731), .D(g24333), .CK(clk));
DFFX1 gate732(.Q (g1174), .QB (line732), .D(g24334), .CK(clk));
DFFX1 gate733(.Q (g1175), .QB (line733), .D(g24335), .CK(clk));
DFFX1 gate734(.Q (g1142), .QB (line734), .D(g25150), .CK(clk));
DFFX1 gate735(.Q (g1145), .QB (line735), .D(g25142), .CK(clk));
DFFX1 gate736(.Q (g1148), .QB (line736), .D(g25143), .CK(clk));
DFFX1 gate737(.Q (g1164), .QB (line737), .D(g25147), .CK(clk));
DFFX1 gate738(.Q (g1165), .QB (line738), .D(g25148), .CK(clk));
DFFX1 gate739(.Q (g1166), .QB (line739), .D(g25149), .CK(clk));
DFFX1 gate740(.Q (g1167), .QB (line740), .D(g24330), .CK(clk));
DFFX1 gate741(.Q (g1171), .QB (line741), .D(g24331), .CK(clk));
DFFX1 gate742(.Q (g1151), .QB (line742), .D(g24332), .CK(clk));
DFFX1 gate743(.Q (g1152), .QB (line743), .D(g25144), .CK(clk));
DFFX1 gate744(.Q (g1155), .QB (line744), .D(g25145), .CK(clk));
DFFX1 gate745(.Q (g1158), .QB (line745), .D(g25146), .CK(clk));
DFFX1 gate746(.Q (g1214), .QB (line746), .D(g16470), .CK(clk));
DFFX1 gate747(.Q (g1221), .QB (line747), .D(g1214), .CK(clk));
DFFX1 gate748(.Q (g1228), .QB (line748), .D(g1221), .CK(clk));
DFFX1 gate749(.Q (g1229), .QB (line749), .D(g19033), .CK(clk));
DFFX1 gate750(.Q (g1230), .QB (line750), .D(g1229), .CK(clk));
DFFX1 gate751(.Q (g1234), .QB (line751), .D(g27217), .CK(clk));
DFFX1 gate752(.Q (g1235), .QB (line752), .D(g19034), .CK(clk));
DFFX1 gate753(.Q (g1186), .QB (line753), .D(g1235), .CK(clk));
DFFX1 gate754(.Q (g1244), .QB (line754), .D(g19035), .CK(clk));
DFFX1 gate755(.Q (g1245), .QB (line755), .D(g1244), .CK(clk));
DFFX1 gate756(.Q (g1262), .QB (line756), .D(g28245), .CK(clk));
DFFX1 gate757(.Q (g1263), .QB (line757), .D(g28246), .CK(clk));
DFFX1 gate758(.Q (g1261), .QB (line758), .D(g28247), .CK(clk));
DFFX1 gate759(.Q (g1265), .QB (line759), .D(g28248), .CK(clk));
DFFX1 gate760(.Q (g1266), .QB (line760), .D(g28249), .CK(clk));
DFFX1 gate761(.Q (g1264), .QB (line761), .D(g28250), .CK(clk));
DFFX1 gate762(.Q (g1268), .QB (line762), .D(g28251), .CK(clk));
DFFX1 gate763(.Q (g1269), .QB (line763), .D(g28252), .CK(clk));
DFFX1 gate764(.Q (g1267), .QB (line764), .D(g28253), .CK(clk));
DFFX1 gate765(.Q (g1271), .QB (line765), .D(g28254), .CK(clk));
DFFX1 gate766(.Q (g1272), .QB (line766), .D(g28255), .CK(clk));
DFFX1 gate767(.Q (g1270), .QB (line767), .D(g28256), .CK(clk));
DFFX1 gate768(.Q (g1273), .QB (line768), .D(g25994), .CK(clk));
DFFX1 gate769(.Q (g1276), .QB (line769), .D(g25995), .CK(clk));
DFFX1 gate770(.Q (g1279), .QB (line770), .D(g25996), .CK(clk));
DFFX1 gate771(.Q (g1282), .QB (line771), .D(g25997), .CK(clk));
DFFX1 gate772(.Q (g1285), .QB (line772), .D(g25998), .CK(clk));
DFFX1 gate773(.Q (g1288), .QB (line773), .D(g25999), .CK(clk));
DFFX1 gate774(.Q (g1300), .QB (line774), .D(g29143), .CK(clk));
DFFX1 gate775(.Q (g1303), .QB (line775), .D(g29144), .CK(clk));
DFFX1 gate776(.Q (g1306), .QB (line776), .D(g29145), .CK(clk));
DFFX1 gate777(.Q (g1291), .QB (line777), .D(g29140), .CK(clk));
DFFX1 gate778(.Q (g1294), .QB (line778), .D(g29141), .CK(clk));
DFFX1 gate779(.Q (g1297), .QB (line779), .D(g29142), .CK(clk));
DFFX1 gate780(.Q (g1177), .QB (line780), .D(g27209), .CK(clk));
DFFX1 gate781(.Q (g1180), .QB (line781), .D(g27210), .CK(clk));
DFFX1 gate782(.Q (g1183), .QB (line782), .D(g27211), .CK(clk));
DFFX1 gate783(.Q (g1192), .QB (line783), .D(g8293), .CK(clk));
DFFX1 gate784(.Q (g1193), .QB (line784), .D(g24336), .CK(clk));
DFFX1 gate785(.Q (g1194), .QB (line785), .D(g19029), .CK(clk));
DFFX1 gate786(.Q (g1195), .QB (line786), .D(g19030), .CK(clk));
DFFX1 gate787(.Q (g1200), .QB (line787), .D(g19031), .CK(clk));
DFFX1 gate788(.Q (g1201), .QB (line788), .D(g19032), .CK(clk));
DFFX1 gate789(.Q (g1202), .QB (line789), .D(g27216), .CK(clk));
DFFX1 gate790(.Q (g1203), .QB (line790), .D(g27215), .CK(clk));
DFFX1 gate791(.Q (g1204), .QB (line791), .D(g27214), .CK(clk));
DFFX1 gate792(.Q (g1205), .QB (line792), .D(g27213), .CK(clk));
DFFX1 gate793(.Q (g1206), .QB (line793), .D(g27212), .CK(clk));
DFFX1 gate794(.Q (g1211), .QB (line794), .D(g1206), .CK(clk));
DFFX1 gate795(.Q (g1215), .QB (line795), .D(g13426), .CK(clk));
DFFX1 gate796(.Q (g1216), .QB (line796), .D(g13427), .CK(clk));
DFFX1 gate797(.Q (g1217), .QB (line797), .D(g13428), .CK(clk));
DFFX1 gate798(.Q (g1218), .QB (line798), .D(g13429), .CK(clk));
DFFX1 gate799(.Q (g1219), .QB (line799), .D(g13430), .CK(clk));
DFFX1 gate800(.Q (g1220), .QB (line800), .D(g13431), .CK(clk));
DFFX1 gate801(.Q (g1222), .QB (line801), .D(g13432), .CK(clk));
DFFX1 gate802(.Q (g1223), .QB (line802), .D(g13433), .CK(clk));
DFFX1 gate803(.Q (g1224), .QB (line803), .D(g25993), .CK(clk));
DFFX1 gate804(.Q (g1227), .QB (line804), .D(g13434), .CK(clk));
DFFX1 gate805(.Q (g1309), .QB (line805), .D(g13436), .CK(clk));
DFFX1 gate806(.Q (g1312), .QB (line806), .D(g1309), .CK(clk));
DFFX1 gate807(.Q (g1315), .QB (line807), .D(g1312), .CK(clk));
DFFX1 gate808(.Q (g1316), .QB (line808), .D(g20562), .CK(clk));
DFFX1 gate809(.Q (g1345), .QB (line809), .D(g21944), .CK(clk));
DFFX1 gate810(.Q (g1326), .QB (line810), .D(g23199), .CK(clk));
DFFX1 gate811(.Q (g1319), .QB (line811), .D(g24337), .CK(clk));
DFFX1 gate812(.Q (g1339), .QB (line812), .D(g25151), .CK(clk));
DFFX1 gate813(.Q (g1332), .QB (line813), .D(g26000), .CK(clk));
DFFX1 gate814(.Q (g1346), .QB (line814), .D(g26708), .CK(clk));
DFFX1 gate815(.Q (g1358), .QB (line815), .D(g27218), .CK(clk));
DFFX1 gate816(.Q (g1352), .QB (line816), .D(g27698), .CK(clk));
DFFX1 gate817(.Q (g1365), .QB (line817), .D(g28257), .CK(clk));
DFFX1 gate818(.Q (g1372), .QB (line818), .D(g28682), .CK(clk));
DFFX1 gate819(.Q (g1378), .QB (line819), .D(g29146), .CK(clk));
DFFX1 gate820(.Q (g1385), .QB (line820), .D(g23200), .CK(clk));
DFFX1 gate821(.Q (g1386), .QB (line821), .D(g23201), .CK(clk));
DFFX1 gate822(.Q (g1384), .QB (line822), .D(g23202), .CK(clk));
DFFX1 gate823(.Q (g1388), .QB (line823), .D(g23203), .CK(clk));
DFFX1 gate824(.Q (g1389), .QB (line824), .D(g23204), .CK(clk));
DFFX1 gate825(.Q (g1387), .QB (line825), .D(g23205), .CK(clk));
DFFX1 gate826(.Q (g1391), .QB (line826), .D(g23206), .CK(clk));
DFFX1 gate827(.Q (g1392), .QB (line827), .D(g23207), .CK(clk));
DFFX1 gate828(.Q (g1390), .QB (line828), .D(g23208), .CK(clk));
DFFX1 gate829(.Q (g1394), .QB (line829), .D(g23209), .CK(clk));
DFFX1 gate830(.Q (g1395), .QB (line830), .D(g23210), .CK(clk));
DFFX1 gate831(.Q (g1393), .QB (line831), .D(g23211), .CK(clk));
DFFX1 gate832(.Q (g1397), .QB (line832), .D(g23212), .CK(clk));
DFFX1 gate833(.Q (g1398), .QB (line833), .D(g23213), .CK(clk));
DFFX1 gate834(.Q (g1396), .QB (line834), .D(g23214), .CK(clk));
DFFX1 gate835(.Q (g1400), .QB (line835), .D(g23215), .CK(clk));
DFFX1 gate836(.Q (g1401), .QB (line836), .D(g23216), .CK(clk));
DFFX1 gate837(.Q (g1399), .QB (line837), .D(g23217), .CK(clk));
DFFX1 gate838(.Q (g1403), .QB (line838), .D(g23218), .CK(clk));
DFFX1 gate839(.Q (g1404), .QB (line839), .D(g23219), .CK(clk));
DFFX1 gate840(.Q (g1402), .QB (line840), .D(g23220), .CK(clk));
DFFX1 gate841(.Q (g1406), .QB (line841), .D(g23221), .CK(clk));
DFFX1 gate842(.Q (g1407), .QB (line842), .D(g23222), .CK(clk));
DFFX1 gate843(.Q (g1405), .QB (line843), .D(g23223), .CK(clk));
DFFX1 gate844(.Q (g1409), .QB (line844), .D(g23224), .CK(clk));
DFFX1 gate845(.Q (g1410), .QB (line845), .D(g23225), .CK(clk));
DFFX1 gate846(.Q (g1408), .QB (line846), .D(g23226), .CK(clk));
DFFX1 gate847(.Q (g1412), .QB (line847), .D(g23227), .CK(clk));
DFFX1 gate848(.Q (g1413), .QB (line848), .D(g23228), .CK(clk));
DFFX1 gate849(.Q (g1411), .QB (line849), .D(g23229), .CK(clk));
DFFX1 gate850(.Q (g1415), .QB (line850), .D(g23230), .CK(clk));
DFFX1 gate851(.Q (g1416), .QB (line851), .D(g23231), .CK(clk));
DFFX1 gate852(.Q (g1414), .QB (line852), .D(g23232), .CK(clk));
DFFX1 gate853(.Q (g1418), .QB (line853), .D(g23233), .CK(clk));
DFFX1 gate854(.Q (g1419), .QB (line854), .D(g23234), .CK(clk));
DFFX1 gate855(.Q (g1417), .QB (line855), .D(g23235), .CK(clk));
DFFX1 gate856(.Q (g1421), .QB (line856), .D(g26709), .CK(clk));
DFFX1 gate857(.Q (g1422), .QB (line857), .D(g26710), .CK(clk));
DFFX1 gate858(.Q (g1420), .QB (line858), .D(g26711), .CK(clk));
DFFX1 gate859(.Q (g1424), .QB (line859), .D(g24338), .CK(clk));
DFFX1 gate860(.Q (g1425), .QB (line860), .D(g24339), .CK(clk));
DFFX1 gate861(.Q (g1423), .QB (line861), .D(g24340), .CK(clk));
DFFX1 gate862(.Q (g1520), .QB (line862), .D(g13437), .CK(clk));
DFFX1 gate863(.Q (g1517), .QB (line863), .D(g1520), .CK(clk));
DFFX1 gate864(.Q (g1547), .QB (line864), .D(g1517), .CK(clk));
DFFX1 gate865(.Q (g1512), .QB (line865), .D(g24341), .CK(clk));
DFFX1 gate866(.Q (g1513), .QB (line866), .D(g24342), .CK(clk));
DFFX1 gate867(.Q (g1511), .QB (line867), .D(g24343), .CK(clk));
DFFX1 gate868(.Q (g1515), .QB (line868), .D(g24344), .CK(clk));
DFFX1 gate869(.Q (g1516), .QB (line869), .D(g24345), .CK(clk));
DFFX1 gate870(.Q (g1514), .QB (line870), .D(g24346), .CK(clk));
DFFX1 gate871(.Q (g1524), .QB (line871), .D(g24347), .CK(clk));
DFFX1 gate872(.Q (g1525), .QB (line872), .D(g24348), .CK(clk));
DFFX1 gate873(.Q (g1523), .QB (line873), .D(g24349), .CK(clk));
DFFX1 gate874(.Q (g1527), .QB (line874), .D(g24350), .CK(clk));
DFFX1 gate875(.Q (g1528), .QB (line875), .D(g24351), .CK(clk));
DFFX1 gate876(.Q (g1526), .QB (line876), .D(g24352), .CK(clk));
DFFX1 gate877(.Q (g1530), .QB (line877), .D(g24353), .CK(clk));
DFFX1 gate878(.Q (g1531), .QB (line878), .D(g24354), .CK(clk));
DFFX1 gate879(.Q (g1529), .QB (line879), .D(g24355), .CK(clk));
DFFX1 gate880(.Q (g1533), .QB (line880), .D(g24356), .CK(clk));
DFFX1 gate881(.Q (g1534), .QB (line881), .D(g24357), .CK(clk));
DFFX1 gate882(.Q (g1532), .QB (line882), .D(g24358), .CK(clk));
DFFX1 gate883(.Q (g1536), .QB (line883), .D(g24359), .CK(clk));
DFFX1 gate884(.Q (g1537), .QB (line884), .D(g24360), .CK(clk));
DFFX1 gate885(.Q (g1535), .QB (line885), .D(g24361), .CK(clk));
DFFX1 gate886(.Q (g1539), .QB (line886), .D(g24362), .CK(clk));
DFFX1 gate887(.Q (g1540), .QB (line887), .D(g24363), .CK(clk));
DFFX1 gate888(.Q (g1538), .QB (line888), .D(g24364), .CK(clk));
DFFX1 gate889(.Q (g1542), .QB (line889), .D(g24365), .CK(clk));
DFFX1 gate890(.Q (g1543), .QB (line890), .D(g24366), .CK(clk));
DFFX1 gate891(.Q (g1541), .QB (line891), .D(g24367), .CK(clk));
DFFX1 gate892(.Q (g1545), .QB (line892), .D(g24368), .CK(clk));
DFFX1 gate893(.Q (g1546), .QB (line893), .D(g24369), .CK(clk));
DFFX1 gate894(.Q (g1544), .QB (line894), .D(g24370), .CK(clk));
DFFX1 gate895(.Q (g1551), .QB (line895), .D(g26713), .CK(clk));
DFFX1 gate896(.Q (g1552), .QB (line896), .D(g26714), .CK(clk));
DFFX1 gate897(.Q (g1550), .QB (line897), .D(g26715), .CK(clk));
DFFX1 gate898(.Q (g1554), .QB (line898), .D(g26716), .CK(clk));
DFFX1 gate899(.Q (g1555), .QB (line899), .D(g26717), .CK(clk));
DFFX1 gate900(.Q (g1553), .QB (line900), .D(g26718), .CK(clk));
DFFX1 gate901(.Q (g1557), .QB (line901), .D(g26719), .CK(clk));
DFFX1 gate902(.Q (g1558), .QB (line902), .D(g26720), .CK(clk));
DFFX1 gate903(.Q (g1556), .QB (line903), .D(g26721), .CK(clk));
DFFX1 gate904(.Q (g1560), .QB (line904), .D(g26722), .CK(clk));
DFFX1 gate905(.Q (g1561), .QB (line905), .D(g26723), .CK(clk));
DFFX1 gate906(.Q (g1559), .QB (line906), .D(g26724), .CK(clk));
DFFX1 gate907(.Q (g1567), .QB (line907), .D(g30536), .CK(clk));
DFFX1 gate908(.Q (g1570), .QB (line908), .D(g30537), .CK(clk));
DFFX1 gate909(.Q (g1573), .QB (line909), .D(g30538), .CK(clk));
DFFX1 gate910(.Q (g1612), .QB (line910), .D(g30878), .CK(clk));
DFFX1 gate911(.Q (g1615), .QB (line911), .D(g30879), .CK(clk));
DFFX1 gate912(.Q (g1618), .QB (line912), .D(g30880), .CK(clk));
DFFX1 gate913(.Q (g1576), .QB (line913), .D(g30872), .CK(clk));
DFFX1 gate914(.Q (g1579), .QB (line914), .D(g30873), .CK(clk));
DFFX1 gate915(.Q (g1582), .QB (line915), .D(g30874), .CK(clk));
DFFX1 gate916(.Q (g1621), .QB (line916), .D(g30881), .CK(clk));
DFFX1 gate917(.Q (g1624), .QB (line917), .D(g30882), .CK(clk));
DFFX1 gate918(.Q (g1627), .QB (line918), .D(g30883), .CK(clk));
DFFX1 gate919(.Q (g1585), .QB (line919), .D(g30539), .CK(clk));
DFFX1 gate920(.Q (g1588), .QB (line920), .D(g30540), .CK(clk));
DFFX1 gate921(.Q (g1591), .QB (line921), .D(g30541), .CK(clk));
DFFX1 gate922(.Q (g1630), .QB (line922), .D(g30545), .CK(clk));
DFFX1 gate923(.Q (g1633), .QB (line923), .D(g30546), .CK(clk));
DFFX1 gate924(.Q (g1636), .QB (line924), .D(g30547), .CK(clk));
DFFX1 gate925(.Q (g1594), .QB (line925), .D(g30542), .CK(clk));
DFFX1 gate926(.Q (g1597), .QB (line926), .D(g30543), .CK(clk));
DFFX1 gate927(.Q (g1600), .QB (line927), .D(g30544), .CK(clk));
DFFX1 gate928(.Q (g1639), .QB (line928), .D(g30548), .CK(clk));
DFFX1 gate929(.Q (g1642), .QB (line929), .D(g30549), .CK(clk));
DFFX1 gate930(.Q (g1645), .QB (line930), .D(g30550), .CK(clk));
DFFX1 gate931(.Q (g1603), .QB (line931), .D(g30875), .CK(clk));
DFFX1 gate932(.Q (g1606), .QB (line932), .D(g30876), .CK(clk));
DFFX1 gate933(.Q (g1609), .QB (line933), .D(g30877), .CK(clk));
DFFX1 gate934(.Q (g1648), .QB (line934), .D(g30884), .CK(clk));
DFFX1 gate935(.Q (g1651), .QB (line935), .D(g30885), .CK(clk));
DFFX1 gate936(.Q (g1654), .QB (line936), .D(g30886), .CK(clk));
DFFX1 gate937(.Q (g1466), .QB (line937), .D(g26001), .CK(clk));
DFFX1 gate938(.Q (g1462), .QB (line938), .D(g26712), .CK(clk));
DFFX1 gate939(.Q (g1457), .QB (line939), .D(g27219), .CK(clk));
DFFX1 gate940(.Q (g1453), .QB (line940), .D(g27699), .CK(clk));
DFFX1 gate941(.Q (g1448), .QB (line941), .D(g28258), .CK(clk));
DFFX1 gate942(.Q (g1444), .QB (line942), .D(g28683), .CK(clk));
DFFX1 gate943(.Q (g1439), .QB (line943), .D(g29147), .CK(clk));
DFFX1 gate944(.Q (g1435), .QB (line944), .D(g29427), .CK(clk));
DFFX1 gate945(.Q (g1430), .QB (line945), .D(g29641), .CK(clk));
DFFX1 gate946(.Q (g1426), .QB (line946), .D(g29802), .CK(clk));
DFFX1 gate947(.Q (g1562), .QB (line947), .D(g20563), .CK(clk));
DFFX1 gate948(.Q (g1564), .QB (line948), .D(g1562), .CK(clk));
DFFX1 gate949(.Q (g1563), .QB (line949), .D(g1564), .CK(clk));
DFFX1 gate950(.Q (g1657), .QB (line950), .D(g13438), .CK(clk));
DFFX1 gate951(.Q (g1786), .QB (line951), .D(g1657), .CK(clk));
DFFX1 gate952(.Q (g1782), .QB (line952), .D(g1786), .CK(clk));
DFFX1 gate953(.Q (g1690), .QB (line953), .D(g11550), .CK(clk));
DFFX1 gate954(.Q (g1735), .QB (line954), .D(g28259), .CK(clk));
DFFX1 gate955(.Q (g1724), .QB (line955), .D(g28260), .CK(clk));
DFFX1 gate956(.Q (g1727), .QB (line956), .D(g28261), .CK(clk));
DFFX1 gate957(.Q (g1750), .QB (line957), .D(g28262), .CK(clk));
DFFX1 gate958(.Q (g1739), .QB (line958), .D(g28263), .CK(clk));
DFFX1 gate959(.Q (g1742), .QB (line959), .D(g28264), .CK(clk));
DFFX1 gate960(.Q (g1765), .QB (line960), .D(g28265), .CK(clk));
DFFX1 gate961(.Q (g1754), .QB (line961), .D(g28266), .CK(clk));
DFFX1 gate962(.Q (g1757), .QB (line962), .D(g28267), .CK(clk));
DFFX1 gate963(.Q (g1779), .QB (line963), .D(g28268), .CK(clk));
DFFX1 gate964(.Q (g1769), .QB (line964), .D(g28269), .CK(clk));
DFFX1 gate965(.Q (g1772), .QB (line965), .D(g28270), .CK(clk));
DFFX1 gate966(.Q (g1789), .QB (line966), .D(g29434), .CK(clk));
DFFX1 gate967(.Q (g1792), .QB (line967), .D(g29435), .CK(clk));
DFFX1 gate968(.Q (g1795), .QB (line968), .D(g29436), .CK(clk));
DFFX1 gate969(.Q (g1798), .QB (line969), .D(g29645), .CK(clk));
DFFX1 gate970(.Q (g1801), .QB (line970), .D(g29646), .CK(clk));
DFFX1 gate971(.Q (g1804), .QB (line971), .D(g29647), .CK(clk));
DFFX1 gate972(.Q (g1808), .QB (line972), .D(g29437), .CK(clk));
DFFX1 gate973(.Q (g1809), .QB (line973), .D(g29438), .CK(clk));
DFFX1 gate974(.Q (g1807), .QB (line974), .D(g29439), .CK(clk));
DFFX1 gate975(.Q (g1810), .QB (line975), .D(g27700), .CK(clk));
DFFX1 gate976(.Q (g1813), .QB (line976), .D(g27701), .CK(clk));
DFFX1 gate977(.Q (g1816), .QB (line977), .D(g27702), .CK(clk));
DFFX1 gate978(.Q (g1819), .QB (line978), .D(g27703), .CK(clk));
DFFX1 gate979(.Q (g1822), .QB (line979), .D(g27704), .CK(clk));
DFFX1 gate980(.Q (g1825), .QB (line980), .D(g27705), .CK(clk));
DFFX1 gate981(.Q (g1829), .QB (line981), .D(g28684), .CK(clk));
DFFX1 gate982(.Q (g1830), .QB (line982), .D(g28685), .CK(clk));
DFFX1 gate983(.Q (g1828), .QB (line983), .D(g28686), .CK(clk));
DFFX1 gate984(.Q (g1693), .QB (line984), .D(g29803), .CK(clk));
DFFX1 gate985(.Q (g1694), .QB (line985), .D(g29804), .CK(clk));
DFFX1 gate986(.Q (g1695), .QB (line986), .D(g29805), .CK(clk));
DFFX1 gate987(.Q (g1696), .QB (line987), .D(g30887), .CK(clk));
DFFX1 gate988(.Q (g1697), .QB (line988), .D(g30888), .CK(clk));
DFFX1 gate989(.Q (g1698), .QB (line989), .D(g30889), .CK(clk));
DFFX1 gate990(.Q (g1699), .QB (line990), .D(g30716), .CK(clk));
DFFX1 gate991(.Q (g1700), .QB (line991), .D(g30717), .CK(clk));
DFFX1 gate992(.Q (g1701), .QB (line992), .D(g30718), .CK(clk));
DFFX1 gate993(.Q (g1703), .QB (line993), .D(g29642), .CK(clk));
DFFX1 gate994(.Q (g1704), .QB (line994), .D(g29643), .CK(clk));
DFFX1 gate995(.Q (g1702), .QB (line995), .D(g29644), .CK(clk));
DFFX1 gate996(.Q (g1784), .QB (line996), .D(g27221), .CK(clk));
DFFX1 gate997(.Q (g1785), .QB (line997), .D(g27222), .CK(clk));
DFFX1 gate998(.Q (g1783), .QB (line998), .D(g27223), .CK(clk));
DFFX1 gate999(.Q (g1831), .QB (line999), .D(g11563), .CK(clk));
DFFX1 gate1000(.Q (g1832), .QB (line1000), .D(g1831), .CK(clk));
DFFX1 gate1001(.Q (g1833), .QB (line1001), .D(g11564), .CK(clk));
DFFX1 gate1002(.Q (g1834), .QB (line1002), .D(g1833), .CK(clk));
DFFX1 gate1003(.Q (g1835), .QB (line1003), .D(g11565), .CK(clk));
DFFX1 gate1004(.Q (g1660), .QB (line1004), .D(g1835), .CK(clk));
DFFX1 gate1005(.Q (g1661), .QB (line1005), .D(g11545), .CK(clk));
DFFX1 gate1006(.Q (g1662), .QB (line1006), .D(g1661), .CK(clk));
DFFX1 gate1007(.Q (g1663), .QB (line1007), .D(g11546), .CK(clk));
DFFX1 gate1008(.Q (g1664), .QB (line1008), .D(g1663), .CK(clk));
DFFX1 gate1009(.Q (g1665), .QB (line1009), .D(g11547), .CK(clk));
DFFX1 gate1010(.Q (g1666), .QB (line1010), .D(g1665), .CK(clk));
DFFX1 gate1011(.Q (g1667), .QB (line1011), .D(g11548), .CK(clk));
DFFX1 gate1012(.Q (g1668), .QB (line1012), .D(g1667), .CK(clk));
DFFX1 gate1013(.Q (g1669), .QB (line1013), .D(g11549), .CK(clk));
DFFX1 gate1014(.Q (g1670), .QB (line1014), .D(g1669), .CK(clk));
DFFX1 gate1015(.Q (g1671), .QB (line1015), .D(g13439), .CK(clk));
DFFX1 gate1016(.Q (g1672), .QB (line1016), .D(g1671), .CK(clk));
DFFX1 gate1017(.Q (g1680), .QB (line1017), .D(g19036), .CK(clk));
DFFX1 gate1018(.Q (g1686), .QB (line1018), .D(g29428), .CK(clk));
DFFX1 gate1019(.Q (g1689), .QB (line1019), .D(g29429), .CK(clk));
DFFX1 gate1020(.Q (g1678), .QB (line1020), .D(g29430), .CK(clk));
DFFX1 gate1021(.Q (g1677), .QB (line1021), .D(g29431), .CK(clk));
DFFX1 gate1022(.Q (g1676), .QB (line1022), .D(g29432), .CK(clk));
DFFX1 gate1023(.Q (g1675), .QB (line1023), .D(g29433), .CK(clk));
DFFX1 gate1024(.Q (g1685), .QB (line1024), .D(g19040), .CK(clk));
DFFX1 gate1025(.Q (g1684), .QB (line1025), .D(g19039), .CK(clk));
DFFX1 gate1026(.Q (g1683), .QB (line1026), .D(g19038), .CK(clk));
DFFX1 gate1027(.Q (g1682), .QB (line1027), .D(g19037), .CK(clk));
DFFX1 gate1028(.Q (g1681), .QB (line1028), .D(g25152), .CK(clk));
DFFX1 gate1029(.Q (g1679), .QB (line1029), .D(g27220), .CK(clk));
DFFX1 gate1030(.Q (g1723), .QB (line1030), .D(g11551), .CK(clk));
DFFX1 gate1031(.Q (g1730), .QB (line1031), .D(g1723), .CK(clk));
DFFX1 gate1032(.Q (g1731), .QB (line1032), .D(g11552), .CK(clk));
DFFX1 gate1033(.Q (g1732), .QB (line1033), .D(g1731), .CK(clk));
DFFX1 gate1034(.Q (g1733), .QB (line1034), .D(g11553), .CK(clk));
DFFX1 gate1035(.Q (g1734), .QB (line1035), .D(g1733), .CK(clk));
DFFX1 gate1036(.Q (g1738), .QB (line1036), .D(g11554), .CK(clk));
DFFX1 gate1037(.Q (g1745), .QB (line1037), .D(g1738), .CK(clk));
DFFX1 gate1038(.Q (g1746), .QB (line1038), .D(g11555), .CK(clk));
DFFX1 gate1039(.Q (g1747), .QB (line1039), .D(g1746), .CK(clk));
DFFX1 gate1040(.Q (g1748), .QB (line1040), .D(g11556), .CK(clk));
DFFX1 gate1041(.Q (g1749), .QB (line1041), .D(g1748), .CK(clk));
DFFX1 gate1042(.Q (g1753), .QB (line1042), .D(g11557), .CK(clk));
DFFX1 gate1043(.Q (g1760), .QB (line1043), .D(g1753), .CK(clk));
DFFX1 gate1044(.Q (g1761), .QB (line1044), .D(g11558), .CK(clk));
DFFX1 gate1045(.Q (g1762), .QB (line1045), .D(g1761), .CK(clk));
DFFX1 gate1046(.Q (g1763), .QB (line1046), .D(g11559), .CK(clk));
DFFX1 gate1047(.Q (g1764), .QB (line1047), .D(g1763), .CK(clk));
DFFX1 gate1048(.Q (g1768), .QB (line1048), .D(g11560), .CK(clk));
DFFX1 gate1049(.Q (g1775), .QB (line1049), .D(g1768), .CK(clk));
DFFX1 gate1050(.Q (g1776), .QB (line1050), .D(g11561), .CK(clk));
DFFX1 gate1051(.Q (g1777), .QB (line1051), .D(g1776), .CK(clk));
DFFX1 gate1052(.Q (g1778), .QB (line1052), .D(g11562), .CK(clk));
DFFX1 gate1053(.Q (g1705), .QB (line1053), .D(g1778), .CK(clk));
DFFX1 gate1054(.Q (g1706), .QB (line1054), .D(g13440), .CK(clk));
DFFX1 gate1055(.Q (g1712), .QB (line1055), .D(g1706), .CK(clk));
DFFX1 gate1056(.Q (g1718), .QB (line1056), .D(g1712), .CK(clk));
DFFX1 gate1057(.Q (g1925), .QB (line1057), .D(g13451), .CK(clk));
DFFX1 gate1058(.Q (g1931), .QB (line1058), .D(g1925), .CK(clk));
DFFX1 gate1059(.Q (g1930), .QB (line1059), .D(g1931), .CK(clk));
DFFX1 gate1060(.Q (g1934), .QB (line1060), .D(g23236), .CK(clk));
DFFX1 gate1061(.Q (g1937), .QB (line1061), .D(g20564), .CK(clk));
DFFX1 gate1062(.Q (g1890), .QB (line1062), .D(g20565), .CK(clk));
DFFX1 gate1063(.Q (g1893), .QB (line1063), .D(g16471), .CK(clk));
DFFX1 gate1064(.Q (g1903), .QB (line1064), .D(g1893), .CK(clk));
DFFX1 gate1065(.Q (g1904), .QB (line1065), .D(g1903), .CK(clk));
DFFX1 gate1066(.Q (g1944), .QB (line1066), .D(g11566), .CK(clk));
DFFX1 gate1067(.Q (g1949), .QB (line1067), .D(g1944), .CK(clk));
DFFX1 gate1068(.Q (g1950), .QB (line1068), .D(g11569), .CK(clk));
DFFX1 gate1069(.Q (g1951), .QB (line1069), .D(g1950), .CK(clk));
DFFX1 gate1070(.Q (g1952), .QB (line1070), .D(g11570), .CK(clk));
DFFX1 gate1071(.Q (g1953), .QB (line1071), .D(g1952), .CK(clk));
DFFX1 gate1072(.Q (g1954), .QB (line1072), .D(g11571), .CK(clk));
DFFX1 gate1073(.Q (g1945), .QB (line1073), .D(g1954), .CK(clk));
DFFX1 gate1074(.Q (g1946), .QB (line1074), .D(g11567), .CK(clk));
DFFX1 gate1075(.Q (g1947), .QB (line1075), .D(g1946), .CK(clk));
DFFX1 gate1076(.Q (g1948), .QB (line1076), .D(g11568), .CK(clk));
DFFX1 gate1077(.Q (g1870), .QB (line1077), .D(g1948), .CK(clk));
DFFX1 gate1078(.Q (g1855), .QB (line1078), .D(g13441), .CK(clk));
DFFX1 gate1079(.Q (g1862), .QB (line1079), .D(g1855), .CK(clk));
DFFX1 gate1080(.Q (g1866), .QB (line1080), .D(g1862), .CK(clk));
DFFX1 gate1081(.Q (g1867), .QB (line1081), .D(g24374), .CK(clk));
DFFX1 gate1082(.Q (g1868), .QB (line1082), .D(g24375), .CK(clk));
DFFX1 gate1083(.Q (g1869), .QB (line1083), .D(g24376), .CK(clk));
DFFX1 gate1084(.Q (g1836), .QB (line1084), .D(g25161), .CK(clk));
DFFX1 gate1085(.Q (g1839), .QB (line1085), .D(g25153), .CK(clk));
DFFX1 gate1086(.Q (g1842), .QB (line1086), .D(g25154), .CK(clk));
DFFX1 gate1087(.Q (g1858), .QB (line1087), .D(g25158), .CK(clk));
DFFX1 gate1088(.Q (g1859), .QB (line1088), .D(g25159), .CK(clk));
DFFX1 gate1089(.Q (g1860), .QB (line1089), .D(g25160), .CK(clk));
DFFX1 gate1090(.Q (g1861), .QB (line1090), .D(g24371), .CK(clk));
DFFX1 gate1091(.Q (g1865), .QB (line1091), .D(g24372), .CK(clk));
DFFX1 gate1092(.Q (g1845), .QB (line1092), .D(g24373), .CK(clk));
DFFX1 gate1093(.Q (g1846), .QB (line1093), .D(g25155), .CK(clk));
DFFX1 gate1094(.Q (g1849), .QB (line1094), .D(g25156), .CK(clk));
DFFX1 gate1095(.Q (g1852), .QB (line1095), .D(g25157), .CK(clk));
DFFX1 gate1096(.Q (g1908), .QB (line1096), .D(g16472), .CK(clk));
DFFX1 gate1097(.Q (g1915), .QB (line1097), .D(g1908), .CK(clk));
DFFX1 gate1098(.Q (g1922), .QB (line1098), .D(g1915), .CK(clk));
DFFX1 gate1099(.Q (g1923), .QB (line1099), .D(g19045), .CK(clk));
DFFX1 gate1100(.Q (g1924), .QB (line1100), .D(g1923), .CK(clk));
DFFX1 gate1101(.Q (g1928), .QB (line1101), .D(g29445), .CK(clk));
DFFX1 gate1102(.Q (g1929), .QB (line1102), .D(g19046), .CK(clk));
DFFX1 gate1103(.Q (g1880), .QB (line1103), .D(g1929), .CK(clk));
DFFX1 gate1104(.Q (g1938), .QB (line1104), .D(g19047), .CK(clk));
DFFX1 gate1105(.Q (g1939), .QB (line1105), .D(g1938), .CK(clk));
DFFX1 gate1106(.Q (g1956), .QB (line1106), .D(g28271), .CK(clk));
DFFX1 gate1107(.Q (g1957), .QB (line1107), .D(g28272), .CK(clk));
DFFX1 gate1108(.Q (g1955), .QB (line1108), .D(g28273), .CK(clk));
DFFX1 gate1109(.Q (g1959), .QB (line1109), .D(g28274), .CK(clk));
DFFX1 gate1110(.Q (g1960), .QB (line1110), .D(g28275), .CK(clk));
DFFX1 gate1111(.Q (g1958), .QB (line1111), .D(g28276), .CK(clk));
DFFX1 gate1112(.Q (g1962), .QB (line1112), .D(g28277), .CK(clk));
DFFX1 gate1113(.Q (g1963), .QB (line1113), .D(g28278), .CK(clk));
DFFX1 gate1114(.Q (g1961), .QB (line1114), .D(g28279), .CK(clk));
DFFX1 gate1115(.Q (g1965), .QB (line1115), .D(g28280), .CK(clk));
DFFX1 gate1116(.Q (g1966), .QB (line1116), .D(g28281), .CK(clk));
DFFX1 gate1117(.Q (g1964), .QB (line1117), .D(g28282), .CK(clk));
DFFX1 gate1118(.Q (g1967), .QB (line1118), .D(g26003), .CK(clk));
DFFX1 gate1119(.Q (g1970), .QB (line1119), .D(g26004), .CK(clk));
DFFX1 gate1120(.Q (g1973), .QB (line1120), .D(g26005), .CK(clk));
DFFX1 gate1121(.Q (g1976), .QB (line1121), .D(g26006), .CK(clk));
DFFX1 gate1122(.Q (g1979), .QB (line1122), .D(g26007), .CK(clk));
DFFX1 gate1123(.Q (g1982), .QB (line1123), .D(g26008), .CK(clk));
DFFX1 gate1124(.Q (g1994), .QB (line1124), .D(g29151), .CK(clk));
DFFX1 gate1125(.Q (g1997), .QB (line1125), .D(g29152), .CK(clk));
DFFX1 gate1126(.Q (g2000), .QB (line1126), .D(g29153), .CK(clk));
DFFX1 gate1127(.Q (g1985), .QB (line1127), .D(g29148), .CK(clk));
DFFX1 gate1128(.Q (g1988), .QB (line1128), .D(g29149), .CK(clk));
DFFX1 gate1129(.Q (g1991), .QB (line1129), .D(g29150), .CK(clk));
DFFX1 gate1130(.Q (g1871), .QB (line1130), .D(g27224), .CK(clk));
DFFX1 gate1131(.Q (g1874), .QB (line1131), .D(g27225), .CK(clk));
DFFX1 gate1132(.Q (g1877), .QB (line1132), .D(g27226), .CK(clk));
DFFX1 gate1133(.Q (g1886), .QB (line1133), .D(g8302), .CK(clk));
DFFX1 gate1134(.Q (g1887), .QB (line1134), .D(g24377), .CK(clk));
DFFX1 gate1135(.Q (g1888), .QB (line1135), .D(g19041), .CK(clk));
DFFX1 gate1136(.Q (g1889), .QB (line1136), .D(g19042), .CK(clk));
DFFX1 gate1137(.Q (g1894), .QB (line1137), .D(g19043), .CK(clk));
DFFX1 gate1138(.Q (g1895), .QB (line1138), .D(g19044), .CK(clk));
DFFX1 gate1139(.Q (g1896), .QB (line1139), .D(g29444), .CK(clk));
DFFX1 gate1140(.Q (g1897), .QB (line1140), .D(g29443), .CK(clk));
DFFX1 gate1141(.Q (g1898), .QB (line1141), .D(g29442), .CK(clk));
DFFX1 gate1142(.Q (g1899), .QB (line1142), .D(g29441), .CK(clk));
DFFX1 gate1143(.Q (g1900), .QB (line1143), .D(g29440), .CK(clk));
DFFX1 gate1144(.Q (g1905), .QB (line1144), .D(g1900), .CK(clk));
DFFX1 gate1145(.Q (g1909), .QB (line1145), .D(g13442), .CK(clk));
DFFX1 gate1146(.Q (g1910), .QB (line1146), .D(g13443), .CK(clk));
DFFX1 gate1147(.Q (g1911), .QB (line1147), .D(g13444), .CK(clk));
DFFX1 gate1148(.Q (g1912), .QB (line1148), .D(g13445), .CK(clk));
DFFX1 gate1149(.Q (g1913), .QB (line1149), .D(g13446), .CK(clk));
DFFX1 gate1150(.Q (g1914), .QB (line1150), .D(g13447), .CK(clk));
DFFX1 gate1151(.Q (g1916), .QB (line1151), .D(g13448), .CK(clk));
DFFX1 gate1152(.Q (g1917), .QB (line1152), .D(g13449), .CK(clk));
DFFX1 gate1153(.Q (g1918), .QB (line1153), .D(g26002), .CK(clk));
DFFX1 gate1154(.Q (g1921), .QB (line1154), .D(g13450), .CK(clk));
DFFX1 gate1155(.Q (g2003), .QB (line1155), .D(g13452), .CK(clk));
DFFX1 gate1156(.Q (g2006), .QB (line1156), .D(g2003), .CK(clk));
DFFX1 gate1157(.Q (g2009), .QB (line1157), .D(g2006), .CK(clk));
DFFX1 gate1158(.Q (g2010), .QB (line1158), .D(g20566), .CK(clk));
DFFX1 gate1159(.Q (g2039), .QB (line1159), .D(g21945), .CK(clk));
DFFX1 gate1160(.Q (g2020), .QB (line1160), .D(g23237), .CK(clk));
DFFX1 gate1161(.Q (g2013), .QB (line1161), .D(g24378), .CK(clk));
DFFX1 gate1162(.Q (g2033), .QB (line1162), .D(g25162), .CK(clk));
DFFX1 gate1163(.Q (g2026), .QB (line1163), .D(g26009), .CK(clk));
DFFX1 gate1164(.Q (g2040), .QB (line1164), .D(g26725), .CK(clk));
DFFX1 gate1165(.Q (g2052), .QB (line1165), .D(g27227), .CK(clk));
DFFX1 gate1166(.Q (g2046), .QB (line1166), .D(g27706), .CK(clk));
DFFX1 gate1167(.Q (g2059), .QB (line1167), .D(g28283), .CK(clk));
DFFX1 gate1168(.Q (g2066), .QB (line1168), .D(g28687), .CK(clk));
DFFX1 gate1169(.Q (g2072), .QB (line1169), .D(g29154), .CK(clk));
DFFX1 gate1170(.Q (g2079), .QB (line1170), .D(g23238), .CK(clk));
DFFX1 gate1171(.Q (g2080), .QB (line1171), .D(g23239), .CK(clk));
DFFX1 gate1172(.Q (g2078), .QB (line1172), .D(g23240), .CK(clk));
DFFX1 gate1173(.Q (g2082), .QB (line1173), .D(g23241), .CK(clk));
DFFX1 gate1174(.Q (g2083), .QB (line1174), .D(g23242), .CK(clk));
DFFX1 gate1175(.Q (g2081), .QB (line1175), .D(g23243), .CK(clk));
DFFX1 gate1176(.Q (g2085), .QB (line1176), .D(g23244), .CK(clk));
DFFX1 gate1177(.Q (g2086), .QB (line1177), .D(g23245), .CK(clk));
DFFX1 gate1178(.Q (g2084), .QB (line1178), .D(g23246), .CK(clk));
DFFX1 gate1179(.Q (g2088), .QB (line1179), .D(g23247), .CK(clk));
DFFX1 gate1180(.Q (g2089), .QB (line1180), .D(g23248), .CK(clk));
DFFX1 gate1181(.Q (g2087), .QB (line1181), .D(g23249), .CK(clk));
DFFX1 gate1182(.Q (g2091), .QB (line1182), .D(g23250), .CK(clk));
DFFX1 gate1183(.Q (g2092), .QB (line1183), .D(g23251), .CK(clk));
DFFX1 gate1184(.Q (g2090), .QB (line1184), .D(g23252), .CK(clk));
DFFX1 gate1185(.Q (g2094), .QB (line1185), .D(g23253), .CK(clk));
DFFX1 gate1186(.Q (g2095), .QB (line1186), .D(g23254), .CK(clk));
DFFX1 gate1187(.Q (g2093), .QB (line1187), .D(g23255), .CK(clk));
DFFX1 gate1188(.Q (g2097), .QB (line1188), .D(g23256), .CK(clk));
DFFX1 gate1189(.Q (g2098), .QB (line1189), .D(g23257), .CK(clk));
DFFX1 gate1190(.Q (g2096), .QB (line1190), .D(g23258), .CK(clk));
DFFX1 gate1191(.Q (g2100), .QB (line1191), .D(g23259), .CK(clk));
DFFX1 gate1192(.Q (g2101), .QB (line1192), .D(g23260), .CK(clk));
DFFX1 gate1193(.Q (g2099), .QB (line1193), .D(g23261), .CK(clk));
DFFX1 gate1194(.Q (g2103), .QB (line1194), .D(g23262), .CK(clk));
DFFX1 gate1195(.Q (g2104), .QB (line1195), .D(g23263), .CK(clk));
DFFX1 gate1196(.Q (g2102), .QB (line1196), .D(g23264), .CK(clk));
DFFX1 gate1197(.Q (g2106), .QB (line1197), .D(g23265), .CK(clk));
DFFX1 gate1198(.Q (g2107), .QB (line1198), .D(g23266), .CK(clk));
DFFX1 gate1199(.Q (g2105), .QB (line1199), .D(g23267), .CK(clk));
DFFX1 gate1200(.Q (g2109), .QB (line1200), .D(g23268), .CK(clk));
DFFX1 gate1201(.Q (g2110), .QB (line1201), .D(g23269), .CK(clk));
DFFX1 gate1202(.Q (g2108), .QB (line1202), .D(g23270), .CK(clk));
DFFX1 gate1203(.Q (g2112), .QB (line1203), .D(g23271), .CK(clk));
DFFX1 gate1204(.Q (g2113), .QB (line1204), .D(g23272), .CK(clk));
DFFX1 gate1205(.Q (g2111), .QB (line1205), .D(g23273), .CK(clk));
DFFX1 gate1206(.Q (g2115), .QB (line1206), .D(g26726), .CK(clk));
DFFX1 gate1207(.Q (g2116), .QB (line1207), .D(g26727), .CK(clk));
DFFX1 gate1208(.Q (g2114), .QB (line1208), .D(g26728), .CK(clk));
DFFX1 gate1209(.Q (g2118), .QB (line1209), .D(g24379), .CK(clk));
DFFX1 gate1210(.Q (g2119), .QB (line1210), .D(g24380), .CK(clk));
DFFX1 gate1211(.Q (g2117), .QB (line1211), .D(g24381), .CK(clk));
DFFX1 gate1212(.Q (g2214), .QB (line1212), .D(g13453), .CK(clk));
DFFX1 gate1213(.Q (g2211), .QB (line1213), .D(g2214), .CK(clk));
DFFX1 gate1214(.Q (g2241), .QB (line1214), .D(g2211), .CK(clk));
DFFX1 gate1215(.Q (g2206), .QB (line1215), .D(g24382), .CK(clk));
DFFX1 gate1216(.Q (g2207), .QB (line1216), .D(g24383), .CK(clk));
DFFX1 gate1217(.Q (g2205), .QB (line1217), .D(g24384), .CK(clk));
DFFX1 gate1218(.Q (g2209), .QB (line1218), .D(g24385), .CK(clk));
DFFX1 gate1219(.Q (g2210), .QB (line1219), .D(g24386), .CK(clk));
DFFX1 gate1220(.Q (g2208), .QB (line1220), .D(g24387), .CK(clk));
DFFX1 gate1221(.Q (g2218), .QB (line1221), .D(g24388), .CK(clk));
DFFX1 gate1222(.Q (g2219), .QB (line1222), .D(g24389), .CK(clk));
DFFX1 gate1223(.Q (g2217), .QB (line1223), .D(g24390), .CK(clk));
DFFX1 gate1224(.Q (g2221), .QB (line1224), .D(g24391), .CK(clk));
DFFX1 gate1225(.Q (g2222), .QB (line1225), .D(g24392), .CK(clk));
DFFX1 gate1226(.Q (g2220), .QB (line1226), .D(g24393), .CK(clk));
DFFX1 gate1227(.Q (g2224), .QB (line1227), .D(g24394), .CK(clk));
DFFX1 gate1228(.Q (g2225), .QB (line1228), .D(g24395), .CK(clk));
DFFX1 gate1229(.Q (g2223), .QB (line1229), .D(g24396), .CK(clk));
DFFX1 gate1230(.Q (g2227), .QB (line1230), .D(g24397), .CK(clk));
DFFX1 gate1231(.Q (g2228), .QB (line1231), .D(g24398), .CK(clk));
DFFX1 gate1232(.Q (g2226), .QB (line1232), .D(g24399), .CK(clk));
DFFX1 gate1233(.Q (g2230), .QB (line1233), .D(g24400), .CK(clk));
DFFX1 gate1234(.Q (g2231), .QB (line1234), .D(g24401), .CK(clk));
DFFX1 gate1235(.Q (g2229), .QB (line1235), .D(g24402), .CK(clk));
DFFX1 gate1236(.Q (g2233), .QB (line1236), .D(g24403), .CK(clk));
DFFX1 gate1237(.Q (g2234), .QB (line1237), .D(g24404), .CK(clk));
DFFX1 gate1238(.Q (g2232), .QB (line1238), .D(g24405), .CK(clk));
DFFX1 gate1239(.Q (g2236), .QB (line1239), .D(g24406), .CK(clk));
DFFX1 gate1240(.Q (g2237), .QB (line1240), .D(g24407), .CK(clk));
DFFX1 gate1241(.Q (g2235), .QB (line1241), .D(g24408), .CK(clk));
DFFX1 gate1242(.Q (g2239), .QB (line1242), .D(g24409), .CK(clk));
DFFX1 gate1243(.Q (g2240), .QB (line1243), .D(g24410), .CK(clk));
DFFX1 gate1244(.Q (g2238), .QB (line1244), .D(g24411), .CK(clk));
DFFX1 gate1245(.Q (g2245), .QB (line1245), .D(g26730), .CK(clk));
DFFX1 gate1246(.Q (g2246), .QB (line1246), .D(g26731), .CK(clk));
DFFX1 gate1247(.Q (g2244), .QB (line1247), .D(g26732), .CK(clk));
DFFX1 gate1248(.Q (g2248), .QB (line1248), .D(g26733), .CK(clk));
DFFX1 gate1249(.Q (g2249), .QB (line1249), .D(g26734), .CK(clk));
DFFX1 gate1250(.Q (g2247), .QB (line1250), .D(g26735), .CK(clk));
DFFX1 gate1251(.Q (g2251), .QB (line1251), .D(g26736), .CK(clk));
DFFX1 gate1252(.Q (g2252), .QB (line1252), .D(g26737), .CK(clk));
DFFX1 gate1253(.Q (g2250), .QB (line1253), .D(g26738), .CK(clk));
DFFX1 gate1254(.Q (g2254), .QB (line1254), .D(g26739), .CK(clk));
DFFX1 gate1255(.Q (g2255), .QB (line1255), .D(g26740), .CK(clk));
DFFX1 gate1256(.Q (g2253), .QB (line1256), .D(g26741), .CK(clk));
DFFX1 gate1257(.Q (g2261), .QB (line1257), .D(g30551), .CK(clk));
DFFX1 gate1258(.Q (g2264), .QB (line1258), .D(g30552), .CK(clk));
DFFX1 gate1259(.Q (g2267), .QB (line1259), .D(g30553), .CK(clk));
DFFX1 gate1260(.Q (g2306), .QB (line1260), .D(g30896), .CK(clk));
DFFX1 gate1261(.Q (g2309), .QB (line1261), .D(g30897), .CK(clk));
DFFX1 gate1262(.Q (g2312), .QB (line1262), .D(g30898), .CK(clk));
DFFX1 gate1263(.Q (g2270), .QB (line1263), .D(g30890), .CK(clk));
DFFX1 gate1264(.Q (g2273), .QB (line1264), .D(g30891), .CK(clk));
DFFX1 gate1265(.Q (g2276), .QB (line1265), .D(g30892), .CK(clk));
DFFX1 gate1266(.Q (g2315), .QB (line1266), .D(g30899), .CK(clk));
DFFX1 gate1267(.Q (g2318), .QB (line1267), .D(g30900), .CK(clk));
DFFX1 gate1268(.Q (g2321), .QB (line1268), .D(g30901), .CK(clk));
DFFX1 gate1269(.Q (g2279), .QB (line1269), .D(g30554), .CK(clk));
DFFX1 gate1270(.Q (g2282), .QB (line1270), .D(g30555), .CK(clk));
DFFX1 gate1271(.Q (g2285), .QB (line1271), .D(g30556), .CK(clk));
DFFX1 gate1272(.Q (g2324), .QB (line1272), .D(g30560), .CK(clk));
DFFX1 gate1273(.Q (g2327), .QB (line1273), .D(g30561), .CK(clk));
DFFX1 gate1274(.Q (g2330), .QB (line1274), .D(g30562), .CK(clk));
DFFX1 gate1275(.Q (g2288), .QB (line1275), .D(g30557), .CK(clk));
DFFX1 gate1276(.Q (g2291), .QB (line1276), .D(g30558), .CK(clk));
DFFX1 gate1277(.Q (g2294), .QB (line1277), .D(g30559), .CK(clk));
DFFX1 gate1278(.Q (g2333), .QB (line1278), .D(g30563), .CK(clk));
DFFX1 gate1279(.Q (g2336), .QB (line1279), .D(g30564), .CK(clk));
DFFX1 gate1280(.Q (g2339), .QB (line1280), .D(g30565), .CK(clk));
DFFX1 gate1281(.Q (g2297), .QB (line1281), .D(g30893), .CK(clk));
DFFX1 gate1282(.Q (g2300), .QB (line1282), .D(g30894), .CK(clk));
DFFX1 gate1283(.Q (g2303), .QB (line1283), .D(g30895), .CK(clk));
DFFX1 gate1284(.Q (g2342), .QB (line1284), .D(g30902), .CK(clk));
DFFX1 gate1285(.Q (g2345), .QB (line1285), .D(g30903), .CK(clk));
DFFX1 gate1286(.Q (g2348), .QB (line1286), .D(g30904), .CK(clk));
DFFX1 gate1287(.Q (g2160), .QB (line1287), .D(g26010), .CK(clk));
DFFX1 gate1288(.Q (g2156), .QB (line1288), .D(g26729), .CK(clk));
DFFX1 gate1289(.Q (g2151), .QB (line1289), .D(g27228), .CK(clk));
DFFX1 gate1290(.Q (g2147), .QB (line1290), .D(g27707), .CK(clk));
DFFX1 gate1291(.Q (g2142), .QB (line1291), .D(g28284), .CK(clk));
DFFX1 gate1292(.Q (g2138), .QB (line1292), .D(g28688), .CK(clk));
DFFX1 gate1293(.Q (g2133), .QB (line1293), .D(g29155), .CK(clk));
DFFX1 gate1294(.Q (g2129), .QB (line1294), .D(g29446), .CK(clk));
DFFX1 gate1295(.Q (g2124), .QB (line1295), .D(g29648), .CK(clk));
DFFX1 gate1296(.Q (g2120), .QB (line1296), .D(g29806), .CK(clk));
DFFX1 gate1297(.Q (g2256), .QB (line1297), .D(g20567), .CK(clk));
DFFX1 gate1298(.Q (g2258), .QB (line1298), .D(g2256), .CK(clk));
DFFX1 gate1299(.Q (g2257), .QB (line1299), .D(g2258), .CK(clk));
DFFX1 gate1300(.Q (g2351), .QB (line1300), .D(g13454), .CK(clk));
DFFX1 gate1301(.Q (g2480), .QB (line1301), .D(g2351), .CK(clk));
DFFX1 gate1302(.Q (g2476), .QB (line1302), .D(g2480), .CK(clk));
DFFX1 gate1303(.Q (g2384), .QB (line1303), .D(g11577), .CK(clk));
DFFX1 gate1304(.Q (g2429), .QB (line1304), .D(g28285), .CK(clk));
DFFX1 gate1305(.Q (g2418), .QB (line1305), .D(g28286), .CK(clk));
DFFX1 gate1306(.Q (g2421), .QB (line1306), .D(g28287), .CK(clk));
DFFX1 gate1307(.Q (g2444), .QB (line1307), .D(g28288), .CK(clk));
DFFX1 gate1308(.Q (g2433), .QB (line1308), .D(g28289), .CK(clk));
DFFX1 gate1309(.Q (g2436), .QB (line1309), .D(g28290), .CK(clk));
DFFX1 gate1310(.Q (g2459), .QB (line1310), .D(g28291), .CK(clk));
DFFX1 gate1311(.Q (g2448), .QB (line1311), .D(g28292), .CK(clk));
DFFX1 gate1312(.Q (g2451), .QB (line1312), .D(g28293), .CK(clk));
DFFX1 gate1313(.Q (g2473), .QB (line1313), .D(g28294), .CK(clk));
DFFX1 gate1314(.Q (g2463), .QB (line1314), .D(g28295), .CK(clk));
DFFX1 gate1315(.Q (g2466), .QB (line1315), .D(g28296), .CK(clk));
DFFX1 gate1316(.Q (g2483), .QB (line1316), .D(g29447), .CK(clk));
DFFX1 gate1317(.Q (g2486), .QB (line1317), .D(g29448), .CK(clk));
DFFX1 gate1318(.Q (g2489), .QB (line1318), .D(g29449), .CK(clk));
DFFX1 gate1319(.Q (g2492), .QB (line1319), .D(g29652), .CK(clk));
DFFX1 gate1320(.Q (g2495), .QB (line1320), .D(g29653), .CK(clk));
DFFX1 gate1321(.Q (g2498), .QB (line1321), .D(g29654), .CK(clk));
DFFX1 gate1322(.Q (g2502), .QB (line1322), .D(g29450), .CK(clk));
DFFX1 gate1323(.Q (g2503), .QB (line1323), .D(g29451), .CK(clk));
DFFX1 gate1324(.Q (g2501), .QB (line1324), .D(g29452), .CK(clk));
DFFX1 gate1325(.Q (g2504), .QB (line1325), .D(g27708), .CK(clk));
DFFX1 gate1326(.Q (g2507), .QB (line1326), .D(g27709), .CK(clk));
DFFX1 gate1327(.Q (g2510), .QB (line1327), .D(g27710), .CK(clk));
DFFX1 gate1328(.Q (g2513), .QB (line1328), .D(g27711), .CK(clk));
DFFX1 gate1329(.Q (g2516), .QB (line1329), .D(g27712), .CK(clk));
DFFX1 gate1330(.Q (g2519), .QB (line1330), .D(g27713), .CK(clk));
DFFX1 gate1331(.Q (g2523), .QB (line1331), .D(g28689), .CK(clk));
DFFX1 gate1332(.Q (g2524), .QB (line1332), .D(g28690), .CK(clk));
DFFX1 gate1333(.Q (g2522), .QB (line1333), .D(g28691), .CK(clk));
DFFX1 gate1334(.Q (g2387), .QB (line1334), .D(g29807), .CK(clk));
DFFX1 gate1335(.Q (g2388), .QB (line1335), .D(g29808), .CK(clk));
DFFX1 gate1336(.Q (g2389), .QB (line1336), .D(g29809), .CK(clk));
DFFX1 gate1337(.Q (g2390), .QB (line1337), .D(g30905), .CK(clk));
DFFX1 gate1338(.Q (g2391), .QB (line1338), .D(g30906), .CK(clk));
DFFX1 gate1339(.Q (g2392), .QB (line1339), .D(g30907), .CK(clk));
DFFX1 gate1340(.Q (g2393), .QB (line1340), .D(g30719), .CK(clk));
DFFX1 gate1341(.Q (g2394), .QB (line1341), .D(g30720), .CK(clk));
DFFX1 gate1342(.Q (g2395), .QB (line1342), .D(g30721), .CK(clk));
DFFX1 gate1343(.Q (g2397), .QB (line1343), .D(g29649), .CK(clk));
DFFX1 gate1344(.Q (g2398), .QB (line1344), .D(g29650), .CK(clk));
DFFX1 gate1345(.Q (g2396), .QB (line1345), .D(g29651), .CK(clk));
DFFX1 gate1346(.Q (g2478), .QB (line1346), .D(g27230), .CK(clk));
DFFX1 gate1347(.Q (g2479), .QB (line1347), .D(g27231), .CK(clk));
DFFX1 gate1348(.Q (g2477), .QB (line1348), .D(g27232), .CK(clk));
DFFX1 gate1349(.Q (g2525), .QB (line1349), .D(g11590), .CK(clk));
DFFX1 gate1350(.Q (g2526), .QB (line1350), .D(g2525), .CK(clk));
DFFX1 gate1351(.Q (g2527), .QB (line1351), .D(g11591), .CK(clk));
DFFX1 gate1352(.Q (g2528), .QB (line1352), .D(g2527), .CK(clk));
DFFX1 gate1353(.Q (g2529), .QB (line1353), .D(g11592), .CK(clk));
DFFX1 gate1354(.Q (g2354), .QB (line1354), .D(g2529), .CK(clk));
DFFX1 gate1355(.Q (g2355), .QB (line1355), .D(g11572), .CK(clk));
DFFX1 gate1356(.Q (g2356), .QB (line1356), .D(g2355), .CK(clk));
DFFX1 gate1357(.Q (g2357), .QB (line1357), .D(g11573), .CK(clk));
DFFX1 gate1358(.Q (g2358), .QB (line1358), .D(g2357), .CK(clk));
DFFX1 gate1359(.Q (g2359), .QB (line1359), .D(g11574), .CK(clk));
DFFX1 gate1360(.Q (g2360), .QB (line1360), .D(g2359), .CK(clk));
DFFX1 gate1361(.Q (g2361), .QB (line1361), .D(g11575), .CK(clk));
DFFX1 gate1362(.Q (g2362), .QB (line1362), .D(g2361), .CK(clk));
DFFX1 gate1363(.Q (g2363), .QB (line1363), .D(g11576), .CK(clk));
DFFX1 gate1364(.Q (g2364), .QB (line1364), .D(g2363), .CK(clk));
DFFX1 gate1365(.Q (g2365), .QB (line1365), .D(g13455), .CK(clk));
DFFX1 gate1366(.Q (g2366), .QB (line1366), .D(g2365), .CK(clk));
DFFX1 gate1367(.Q (g2374), .QB (line1367), .D(g19048), .CK(clk));
DFFX1 gate1368(.Q (g2380), .QB (line1368), .D(g30314), .CK(clk));
DFFX1 gate1369(.Q (g2383), .QB (line1369), .D(g30315), .CK(clk));
DFFX1 gate1370(.Q (g2372), .QB (line1370), .D(g30316), .CK(clk));
DFFX1 gate1371(.Q (g2371), .QB (line1371), .D(g30317), .CK(clk));
DFFX1 gate1372(.Q (g2370), .QB (line1372), .D(g30318), .CK(clk));
DFFX1 gate1373(.Q (g2369), .QB (line1373), .D(g30319), .CK(clk));
DFFX1 gate1374(.Q (g2379), .QB (line1374), .D(g19052), .CK(clk));
DFFX1 gate1375(.Q (g2378), .QB (line1375), .D(g19051), .CK(clk));
DFFX1 gate1376(.Q (g2377), .QB (line1376), .D(g19050), .CK(clk));
DFFX1 gate1377(.Q (g2376), .QB (line1377), .D(g19049), .CK(clk));
DFFX1 gate1378(.Q (g2375), .QB (line1378), .D(g25163), .CK(clk));
DFFX1 gate1379(.Q (g2373), .QB (line1379), .D(g27229), .CK(clk));
DFFX1 gate1380(.Q (g2417), .QB (line1380), .D(g11578), .CK(clk));
DFFX1 gate1381(.Q (g2424), .QB (line1381), .D(g2417), .CK(clk));
DFFX1 gate1382(.Q (g2425), .QB (line1382), .D(g11579), .CK(clk));
DFFX1 gate1383(.Q (g2426), .QB (line1383), .D(g2425), .CK(clk));
DFFX1 gate1384(.Q (g2427), .QB (line1384), .D(g11580), .CK(clk));
DFFX1 gate1385(.Q (g2428), .QB (line1385), .D(g2427), .CK(clk));
DFFX1 gate1386(.Q (g2432), .QB (line1386), .D(g11581), .CK(clk));
DFFX1 gate1387(.Q (g2439), .QB (line1387), .D(g2432), .CK(clk));
DFFX1 gate1388(.Q (g2440), .QB (line1388), .D(g11582), .CK(clk));
DFFX1 gate1389(.Q (g2441), .QB (line1389), .D(g2440), .CK(clk));
DFFX1 gate1390(.Q (g2442), .QB (line1390), .D(g11583), .CK(clk));
DFFX1 gate1391(.Q (g2443), .QB (line1391), .D(g2442), .CK(clk));
DFFX1 gate1392(.Q (g2447), .QB (line1392), .D(g11584), .CK(clk));
DFFX1 gate1393(.Q (g2454), .QB (line1393), .D(g2447), .CK(clk));
DFFX1 gate1394(.Q (g2455), .QB (line1394), .D(g11585), .CK(clk));
DFFX1 gate1395(.Q (g2456), .QB (line1395), .D(g2455), .CK(clk));
DFFX1 gate1396(.Q (g2457), .QB (line1396), .D(g11586), .CK(clk));
DFFX1 gate1397(.Q (g2458), .QB (line1397), .D(g2457), .CK(clk));
DFFX1 gate1398(.Q (g2462), .QB (line1398), .D(g11587), .CK(clk));
DFFX1 gate1399(.Q (g2469), .QB (line1399), .D(g2462), .CK(clk));
DFFX1 gate1400(.Q (g2470), .QB (line1400), .D(g11588), .CK(clk));
DFFX1 gate1401(.Q (g2471), .QB (line1401), .D(g2470), .CK(clk));
DFFX1 gate1402(.Q (g2472), .QB (line1402), .D(g11589), .CK(clk));
DFFX1 gate1403(.Q (g2399), .QB (line1403), .D(g2472), .CK(clk));
DFFX1 gate1404(.Q (g2400), .QB (line1404), .D(g13456), .CK(clk));
DFFX1 gate1405(.Q (g2406), .QB (line1405), .D(g2400), .CK(clk));
DFFX1 gate1406(.Q (g2412), .QB (line1406), .D(g2406), .CK(clk));
DFFX1 gate1407(.Q (g2619), .QB (line1407), .D(g13467), .CK(clk));
DFFX1 gate1408(.Q (g2625), .QB (line1408), .D(g2619), .CK(clk));
DFFX1 gate1409(.Q (g2624), .QB (line1409), .D(g2625), .CK(clk));
DFFX1 gate1410(.Q (g2628), .QB (line1410), .D(g23274), .CK(clk));
DFFX1 gate1411(.Q (g2631), .QB (line1411), .D(g20568), .CK(clk));
DFFX1 gate1412(.Q (g2584), .QB (line1412), .D(g20569), .CK(clk));
DFFX1 gate1413(.Q (g2587), .QB (line1413), .D(g16473), .CK(clk));
DFFX1 gate1414(.Q (g2597), .QB (line1414), .D(g2587), .CK(clk));
DFFX1 gate1415(.Q (g2598), .QB (line1415), .D(g2597), .CK(clk));
DFFX1 gate1416(.Q (g2638), .QB (line1416), .D(g11593), .CK(clk));
DFFX1 gate1417(.Q (g2643), .QB (line1417), .D(g2638), .CK(clk));
DFFX1 gate1418(.Q (g2644), .QB (line1418), .D(g11596), .CK(clk));
DFFX1 gate1419(.Q (g2645), .QB (line1419), .D(g2644), .CK(clk));
DFFX1 gate1420(.Q (g2646), .QB (line1420), .D(g11597), .CK(clk));
DFFX1 gate1421(.Q (g2647), .QB (line1421), .D(g2646), .CK(clk));
DFFX1 gate1422(.Q (g2648), .QB (line1422), .D(g11598), .CK(clk));
DFFX1 gate1423(.Q (g2639), .QB (line1423), .D(g2648), .CK(clk));
DFFX1 gate1424(.Q (g2640), .QB (line1424), .D(g11594), .CK(clk));
DFFX1 gate1425(.Q (g2641), .QB (line1425), .D(g2640), .CK(clk));
DFFX1 gate1426(.Q (g2642), .QB (line1426), .D(g11595), .CK(clk));
DFFX1 gate1427(.Q (g2564), .QB (line1427), .D(g2642), .CK(clk));
DFFX1 gate1428(.Q (g2549), .QB (line1428), .D(g13457), .CK(clk));
DFFX1 gate1429(.Q (g2556), .QB (line1429), .D(g2549), .CK(clk));
DFFX1 gate1430(.Q (g2560), .QB (line1430), .D(g2556), .CK(clk));
DFFX1 gate1431(.Q (g2561), .QB (line1431), .D(g24415), .CK(clk));
DFFX1 gate1432(.Q (g2562), .QB (line1432), .D(g24416), .CK(clk));
DFFX1 gate1433(.Q (g2563), .QB (line1433), .D(g24417), .CK(clk));
DFFX1 gate1434(.Q (g2530), .QB (line1434), .D(g25172), .CK(clk));
DFFX1 gate1435(.Q (g2533), .QB (line1435), .D(g25164), .CK(clk));
DFFX1 gate1436(.Q (g2536), .QB (line1436), .D(g25165), .CK(clk));
DFFX1 gate1437(.Q (g2552), .QB (line1437), .D(g25169), .CK(clk));
DFFX1 gate1438(.Q (g2553), .QB (line1438), .D(g25170), .CK(clk));
DFFX1 gate1439(.Q (g2554), .QB (line1439), .D(g25171), .CK(clk));
DFFX1 gate1440(.Q (g2555), .QB (line1440), .D(g24412), .CK(clk));
DFFX1 gate1441(.Q (g2559), .QB (line1441), .D(g24413), .CK(clk));
DFFX1 gate1442(.Q (g2539), .QB (line1442), .D(g24414), .CK(clk));
DFFX1 gate1443(.Q (g2540), .QB (line1443), .D(g25166), .CK(clk));
DFFX1 gate1444(.Q (g2543), .QB (line1444), .D(g25167), .CK(clk));
DFFX1 gate1445(.Q (g2546), .QB (line1445), .D(g25168), .CK(clk));
DFFX1 gate1446(.Q (g2602), .QB (line1446), .D(g16474), .CK(clk));
DFFX1 gate1447(.Q (g2609), .QB (line1447), .D(g2602), .CK(clk));
DFFX1 gate1448(.Q (g2616), .QB (line1448), .D(g2609), .CK(clk));
DFFX1 gate1449(.Q (g2617), .QB (line1449), .D(g19057), .CK(clk));
DFFX1 gate1450(.Q (g2618), .QB (line1450), .D(g2617), .CK(clk));
DFFX1 gate1451(.Q (g2622), .QB (line1451), .D(g30325), .CK(clk));
DFFX1 gate1452(.Q (g2623), .QB (line1452), .D(g19058), .CK(clk));
DFFX1 gate1453(.Q (g2574), .QB (line1453), .D(g2623), .CK(clk));
DFFX1 gate1454(.Q (g2632), .QB (line1454), .D(g19059), .CK(clk));
DFFX1 gate1455(.Q (g2633), .QB (line1455), .D(g2632), .CK(clk));
DFFX1 gate1456(.Q (g2650), .QB (line1456), .D(g28297), .CK(clk));
DFFX1 gate1457(.Q (g2651), .QB (line1457), .D(g28298), .CK(clk));
DFFX1 gate1458(.Q (g2649), .QB (line1458), .D(g28299), .CK(clk));
DFFX1 gate1459(.Q (g2653), .QB (line1459), .D(g28300), .CK(clk));
DFFX1 gate1460(.Q (g2654), .QB (line1460), .D(g28301), .CK(clk));
DFFX1 gate1461(.Q (g2652), .QB (line1461), .D(g28302), .CK(clk));
DFFX1 gate1462(.Q (g2656), .QB (line1462), .D(g28303), .CK(clk));
DFFX1 gate1463(.Q (g2657), .QB (line1463), .D(g28304), .CK(clk));
DFFX1 gate1464(.Q (g2655), .QB (line1464), .D(g28305), .CK(clk));
DFFX1 gate1465(.Q (g2659), .QB (line1465), .D(g28306), .CK(clk));
DFFX1 gate1466(.Q (g2660), .QB (line1466), .D(g28307), .CK(clk));
DFFX1 gate1467(.Q (g2658), .QB (line1467), .D(g28308), .CK(clk));
DFFX1 gate1468(.Q (g2661), .QB (line1468), .D(g26012), .CK(clk));
DFFX1 gate1469(.Q (g2664), .QB (line1469), .D(g26013), .CK(clk));
DFFX1 gate1470(.Q (g2667), .QB (line1470), .D(g26014), .CK(clk));
DFFX1 gate1471(.Q (g2670), .QB (line1471), .D(g26015), .CK(clk));
DFFX1 gate1472(.Q (g2673), .QB (line1472), .D(g26016), .CK(clk));
DFFX1 gate1473(.Q (g2676), .QB (line1473), .D(g26017), .CK(clk));
DFFX1 gate1474(.Q (g2688), .QB (line1474), .D(g29159), .CK(clk));
DFFX1 gate1475(.Q (g2691), .QB (line1475), .D(g29160), .CK(clk));
DFFX1 gate1476(.Q (g2694), .QB (line1476), .D(g29161), .CK(clk));
DFFX1 gate1477(.Q (g2679), .QB (line1477), .D(g29156), .CK(clk));
DFFX1 gate1478(.Q (g2682), .QB (line1478), .D(g29157), .CK(clk));
DFFX1 gate1479(.Q (g2685), .QB (line1479), .D(g29158), .CK(clk));
DFFX1 gate1480(.Q (g2565), .QB (line1480), .D(g27233), .CK(clk));
DFFX1 gate1481(.Q (g2568), .QB (line1481), .D(g27234), .CK(clk));
DFFX1 gate1482(.Q (g2571), .QB (line1482), .D(g27235), .CK(clk));
DFFX1 gate1483(.Q (g2580), .QB (line1483), .D(g8311), .CK(clk));
DFFX1 gate1484(.Q (g2581), .QB (line1484), .D(g24418), .CK(clk));
DFFX1 gate1485(.Q (g2582), .QB (line1485), .D(g19053), .CK(clk));
DFFX1 gate1486(.Q (g2583), .QB (line1486), .D(g19054), .CK(clk));
DFFX1 gate1487(.Q (g2588), .QB (line1487), .D(g19055), .CK(clk));
DFFX1 gate1488(.Q (g2589), .QB (line1488), .D(g19056), .CK(clk));
DFFX1 gate1489(.Q (g2590), .QB (line1489), .D(g30324), .CK(clk));
DFFX1 gate1490(.Q (g2591), .QB (line1490), .D(g30323), .CK(clk));
DFFX1 gate1491(.Q (g2592), .QB (line1491), .D(g30322), .CK(clk));
DFFX1 gate1492(.Q (g2593), .QB (line1492), .D(g30321), .CK(clk));
DFFX1 gate1493(.Q (g2594), .QB (line1493), .D(g30320), .CK(clk));
DFFX1 gate1494(.Q (g2599), .QB (line1494), .D(g2594), .CK(clk));
DFFX1 gate1495(.Q (g2603), .QB (line1495), .D(g13458), .CK(clk));
DFFX1 gate1496(.Q (g2604), .QB (line1496), .D(g13459), .CK(clk));
DFFX1 gate1497(.Q (g2605), .QB (line1497), .D(g13460), .CK(clk));
DFFX1 gate1498(.Q (g2606), .QB (line1498), .D(g13461), .CK(clk));
DFFX1 gate1499(.Q (g2607), .QB (line1499), .D(g13462), .CK(clk));
DFFX1 gate1500(.Q (g2608), .QB (line1500), .D(g13463), .CK(clk));
DFFX1 gate1501(.Q (g2610), .QB (line1501), .D(g13464), .CK(clk));
DFFX1 gate1502(.Q (g2611), .QB (line1502), .D(g13465), .CK(clk));
DFFX1 gate1503(.Q (g2612), .QB (line1503), .D(g26011), .CK(clk));
DFFX1 gate1504(.Q (g2615), .QB (line1504), .D(g13466), .CK(clk));
DFFX1 gate1505(.Q (g2697), .QB (line1505), .D(g13468), .CK(clk));
DFFX1 gate1506(.Q (g2700), .QB (line1506), .D(g2697), .CK(clk));
DFFX1 gate1507(.Q (g2703), .QB (line1507), .D(g2700), .CK(clk));
DFFX1 gate1508(.Q (g2704), .QB (line1508), .D(g20570), .CK(clk));
DFFX1 gate1509(.Q (g2733), .QB (line1509), .D(g21946), .CK(clk));
DFFX1 gate1510(.Q (g2714), .QB (line1510), .D(g23275), .CK(clk));
DFFX1 gate1511(.Q (g2707), .QB (line1511), .D(g24419), .CK(clk));
DFFX1 gate1512(.Q (g2727), .QB (line1512), .D(g25173), .CK(clk));
DFFX1 gate1513(.Q (g2720), .QB (line1513), .D(g26018), .CK(clk));
DFFX1 gate1514(.Q (g2734), .QB (line1514), .D(g26742), .CK(clk));
DFFX1 gate1515(.Q (g2746), .QB (line1515), .D(g27236), .CK(clk));
DFFX1 gate1516(.Q (g2740), .QB (line1516), .D(g27714), .CK(clk));
DFFX1 gate1517(.Q (g2753), .QB (line1517), .D(g28309), .CK(clk));
DFFX1 gate1518(.Q (g2760), .QB (line1518), .D(g28692), .CK(clk));
DFFX1 gate1519(.Q (g2766), .QB (line1519), .D(g29162), .CK(clk));
DFFX1 gate1520(.Q (g2773), .QB (line1520), .D(g23276), .CK(clk));
DFFX1 gate1521(.Q (g2774), .QB (line1521), .D(g23277), .CK(clk));
DFFX1 gate1522(.Q (g2772), .QB (line1522), .D(g23278), .CK(clk));
DFFX1 gate1523(.Q (g2776), .QB (line1523), .D(g23279), .CK(clk));
DFFX1 gate1524(.Q (g2777), .QB (line1524), .D(g23280), .CK(clk));
DFFX1 gate1525(.Q (g2775), .QB (line1525), .D(g23281), .CK(clk));
DFFX1 gate1526(.Q (g2779), .QB (line1526), .D(g23282), .CK(clk));
DFFX1 gate1527(.Q (g2780), .QB (line1527), .D(g23283), .CK(clk));
DFFX1 gate1528(.Q (g2778), .QB (line1528), .D(g23284), .CK(clk));
DFFX1 gate1529(.Q (g2782), .QB (line1529), .D(g23285), .CK(clk));
DFFX1 gate1530(.Q (g2783), .QB (line1530), .D(g23286), .CK(clk));
DFFX1 gate1531(.Q (g2781), .QB (line1531), .D(g23287), .CK(clk));
DFFX1 gate1532(.Q (g2785), .QB (line1532), .D(g23288), .CK(clk));
DFFX1 gate1533(.Q (g2786), .QB (line1533), .D(g23289), .CK(clk));
DFFX1 gate1534(.Q (g2784), .QB (line1534), .D(g23290), .CK(clk));
DFFX1 gate1535(.Q (g2788), .QB (line1535), .D(g23291), .CK(clk));
DFFX1 gate1536(.Q (g2789), .QB (line1536), .D(g23292), .CK(clk));
DFFX1 gate1537(.Q (g2787), .QB (line1537), .D(g23293), .CK(clk));
DFFX1 gate1538(.Q (g2791), .QB (line1538), .D(g23294), .CK(clk));
DFFX1 gate1539(.Q (g2792), .QB (line1539), .D(g23295), .CK(clk));
DFFX1 gate1540(.Q (g2790), .QB (line1540), .D(g23296), .CK(clk));
DFFX1 gate1541(.Q (g2794), .QB (line1541), .D(g23297), .CK(clk));
DFFX1 gate1542(.Q (g2795), .QB (line1542), .D(g23298), .CK(clk));
DFFX1 gate1543(.Q (g2793), .QB (line1543), .D(g23299), .CK(clk));
DFFX1 gate1544(.Q (g2797), .QB (line1544), .D(g23300), .CK(clk));
DFFX1 gate1545(.Q (g2798), .QB (line1545), .D(g23301), .CK(clk));
DFFX1 gate1546(.Q (g2796), .QB (line1546), .D(g23302), .CK(clk));
DFFX1 gate1547(.Q (g2800), .QB (line1547), .D(g23303), .CK(clk));
DFFX1 gate1548(.Q (g2801), .QB (line1548), .D(g23304), .CK(clk));
DFFX1 gate1549(.Q (g2799), .QB (line1549), .D(g23305), .CK(clk));
DFFX1 gate1550(.Q (g2803), .QB (line1550), .D(g23306), .CK(clk));
DFFX1 gate1551(.Q (g2804), .QB (line1551), .D(g23307), .CK(clk));
DFFX1 gate1552(.Q (g2802), .QB (line1552), .D(g23308), .CK(clk));
DFFX1 gate1553(.Q (g2806), .QB (line1553), .D(g23309), .CK(clk));
DFFX1 gate1554(.Q (g2807), .QB (line1554), .D(g23310), .CK(clk));
DFFX1 gate1555(.Q (g2805), .QB (line1555), .D(g23311), .CK(clk));
DFFX1 gate1556(.Q (g2809), .QB (line1556), .D(g26743), .CK(clk));
DFFX1 gate1557(.Q (g2810), .QB (line1557), .D(g26744), .CK(clk));
DFFX1 gate1558(.Q (g2808), .QB (line1558), .D(g26745), .CK(clk));
DFFX1 gate1559(.Q (g2812), .QB (line1559), .D(g24420), .CK(clk));
DFFX1 gate1560(.Q (g2813), .QB (line1560), .D(g24421), .CK(clk));
DFFX1 gate1561(.Q (g2811), .QB (line1561), .D(g24422), .CK(clk));
DFFX1 gate1562(.Q (g3054), .QB (line1562), .D(g23317), .CK(clk));
DFFX1 gate1563(.Q (g3079), .QB (line1563), .D(g23318), .CK(clk));
DFFX1 gate1564(.Q (g3080), .QB (line1564), .D(g21965), .CK(clk));
DFFX1 gate1565(.Q (g3043), .QB (line1565), .D(g29453), .CK(clk));
DFFX1 gate1566(.Q (g3044), .QB (line1566), .D(g29454), .CK(clk));
DFFX1 gate1567(.Q (g3045), .QB (line1567), .D(g29455), .CK(clk));
DFFX1 gate1568(.Q (g3046), .QB (line1568), .D(g29456), .CK(clk));
DFFX1 gate1569(.Q (g3047), .QB (line1569), .D(g29457), .CK(clk));
DFFX1 gate1570(.Q (g3048), .QB (line1570), .D(g29458), .CK(clk));
DFFX1 gate1571(.Q (g3049), .QB (line1571), .D(g29459), .CK(clk));
DFFX1 gate1572(.Q (g3050), .QB (line1572), .D(g29460), .CK(clk));
DFFX1 gate1573(.Q (g3051), .QB (line1573), .D(g29655), .CK(clk));
DFFX1 gate1574(.Q (g3052), .QB (line1574), .D(g29972), .CK(clk));
DFFX1 gate1575(.Q (g3053), .QB (line1575), .D(g29973), .CK(clk));
DFFX1 gate1576(.Q (g3055), .QB (line1576), .D(g29974), .CK(clk));
DFFX1 gate1577(.Q (g3056), .QB (line1577), .D(g29975), .CK(clk));
DFFX1 gate1578(.Q (g3057), .QB (line1578), .D(g29976), .CK(clk));
DFFX1 gate1579(.Q (g3058), .QB (line1579), .D(g29977), .CK(clk));
DFFX1 gate1580(.Q (g3059), .QB (line1580), .D(g29978), .CK(clk));
DFFX1 gate1581(.Q (g3060), .QB (line1581), .D(g29979), .CK(clk));
DFFX1 gate1582(.Q (g3061), .QB (line1582), .D(g30119), .CK(clk));
DFFX1 gate1583(.Q (g3062), .QB (line1583), .D(g30908), .CK(clk));
DFFX1 gate1584(.Q (g3063), .QB (line1584), .D(g30909), .CK(clk));
DFFX1 gate1585(.Q (g3064), .QB (line1585), .D(g30910), .CK(clk));
DFFX1 gate1586(.Q (g3065), .QB (line1586), .D(g30911), .CK(clk));
DFFX1 gate1587(.Q (g3066), .QB (line1587), .D(g30912), .CK(clk));
DFFX1 gate1588(.Q (g3067), .QB (line1588), .D(g30913), .CK(clk));
DFFX1 gate1589(.Q (g3068), .QB (line1589), .D(g30914), .CK(clk));
DFFX1 gate1590(.Q (g3069), .QB (line1590), .D(g30915), .CK(clk));
DFFX1 gate1591(.Q (g3070), .QB (line1591), .D(g30940), .CK(clk));
DFFX1 gate1592(.Q (g3071), .QB (line1592), .D(g30980), .CK(clk));
DFFX1 gate1593(.Q (g3072), .QB (line1593), .D(g30981), .CK(clk));
DFFX1 gate1594(.Q (g3073), .QB (line1594), .D(g30982), .CK(clk));
DFFX1 gate1595(.Q (g3074), .QB (line1595), .D(g30983), .CK(clk));
DFFX1 gate1596(.Q (g3075), .QB (line1596), .D(g30984), .CK(clk));
DFFX1 gate1597(.Q (g3076), .QB (line1597), .D(g30985), .CK(clk));
DFFX1 gate1598(.Q (g3077), .QB (line1598), .D(g30986), .CK(clk));
DFFX1 gate1599(.Q (g3078), .QB (line1599), .D(g30987), .CK(clk));
DFFX1 gate1600(.Q (g2997), .QB (line1600), .D(g30989), .CK(clk));
DFFX1 gate1601(.Q (g2993), .QB (line1601), .D(g26748), .CK(clk));
DFFX1 gate1602(.Q (g2998), .QB (line1602), .D(g27238), .CK(clk));
DFFX1 gate1603(.Q (g3006), .QB (line1603), .D(g25177), .CK(clk));
DFFX1 gate1604(.Q (g3002), .QB (line1604), .D(g26021), .CK(clk));
DFFX1 gate1605(.Q (g3013), .QB (line1605), .D(g26750), .CK(clk));
DFFX1 gate1606(.Q (g3010), .QB (line1606), .D(g27239), .CK(clk));
DFFX1 gate1607(.Q (g3024), .QB (line1607), .D(g27716), .CK(clk));
DFFX1 gate1608(.Q (g3018), .QB (line1608), .D(g24425), .CK(clk));
DFFX1 gate1609(.Q (g3028), .QB (line1609), .D(g25176), .CK(clk));
DFFX1 gate1610(.Q (g3036), .QB (line1610), .D(g26022), .CK(clk));
DFFX1 gate1611(.Q (g3032), .QB (line1611), .D(g26749), .CK(clk));
DFFX1 gate1612(.Q (g3040), .QB (line1612), .D(g16497), .CK(clk));
DFFX1 gate1613(.Q (g2986), .QB (line1613), .D(g3040), .CK(clk));
DFFX1 gate1614(.Q (g2987), .QB (line1614), .D(g16495), .CK(clk));
DFFX1 gate1615(.Q (g48), .QB (line1615), .D(g20595), .CK(clk));
DFFX1 gate1616(.Q (g45), .QB (line1616), .D(g20596), .CK(clk));
DFFX1 gate1617(.Q (g42), .QB (line1617), .D(g20597), .CK(clk));
DFFX1 gate1618(.Q (g39), .QB (line1618), .D(g20598), .CK(clk));
DFFX1 gate1619(.Q (g27), .QB (line1619), .D(g20599), .CK(clk));
DFFX1 gate1620(.Q (g30), .QB (line1620), .D(g20600), .CK(clk));
DFFX1 gate1621(.Q (g33), .QB (line1621), .D(g20601), .CK(clk));
DFFX1 gate1622(.Q (g36), .QB (line1622), .D(g20602), .CK(clk));
DFFX1 gate1623(.Q (g3083), .QB (line1623), .D(g20603), .CK(clk));
DFFX1 gate1624(.Q (g26), .QB (line1624), .D(g20604), .CK(clk));
DFFX1 gate1625(.Q (g2992), .QB (line1625), .D(g21966), .CK(clk));
DFFX1 gate1626(.Q (g23), .QB (line1626), .D(g20605), .CK(clk));
DFFX1 gate1627(.Q (g20), .QB (line1627), .D(g20606), .CK(clk));
DFFX1 gate1628(.Q (g17), .QB (line1628), .D(g20607), .CK(clk));
DFFX1 gate1629(.Q (g11), .QB (line1629), .D(g20608), .CK(clk));
DFFX1 gate1630(.Q (g14), .QB (line1630), .D(g20589), .CK(clk));
DFFX1 gate1631(.Q (g5), .QB (line1631), .D(g20590), .CK(clk));
DFFX1 gate1632(.Q (g8), .QB (line1632), .D(g20591), .CK(clk));
DFFX1 gate1633(.Q (g2), .QB (line1633), .D(g20592), .CK(clk));
DFFX1 gate1634(.Q (g2990), .QB (line1634), .D(g20593), .CK(clk));
DFFX1 gate1635(.Q (g2991), .QB (line1635), .D(g21964), .CK(clk));
DFFX1 gate1636(.Q (g1), .QB (line1636), .D(g20594), .CK(clk));
INVX1 gate1637(.O (I13089), .I (g563));
INVX1 gate1638(.O (g562), .I (I13089));
INVX1 gate1639(.O (I13092), .I (g1249));
INVX1 gate1640(.O (g1248), .I (I13092));
INVX1 gate1641(.O (I13095), .I (g1943));
INVX1 gate1642(.O (g1942), .I (I13095));
INVX1 gate1643(.O (I13098), .I (g2637));
INVX1 gate1644(.O (g2636), .I (I13098));
INVX1 gate1645(.O (I13101), .I (g1));
INVX1 gate1646(.O (g3235), .I (I13101));
INVX1 gate1647(.O (I13104), .I (g2));
INVX1 gate1648(.O (g3236), .I (I13104));
INVX1 gate1649(.O (I13107), .I (g5));
INVX1 gate1650(.O (g3237), .I (I13107));
INVX1 gate1651(.O (I13110), .I (g8));
INVX1 gate1652(.O (g3238), .I (I13110));
INVX1 gate1653(.O (I13113), .I (g11));
INVX1 gate1654(.O (g3239), .I (I13113));
INVX1 gate1655(.O (I13116), .I (g14));
INVX1 gate1656(.O (g3240), .I (I13116));
INVX1 gate1657(.O (I13119), .I (g17));
INVX1 gate1658(.O (g3241), .I (I13119));
INVX1 gate1659(.O (I13122), .I (g20));
INVX1 gate1660(.O (g3242), .I (I13122));
INVX1 gate1661(.O (I13125), .I (g23));
INVX1 gate1662(.O (g3243), .I (I13125));
INVX1 gate1663(.O (I13128), .I (g26));
INVX1 gate1664(.O (g3244), .I (I13128));
INVX1 gate1665(.O (I13131), .I (g27));
INVX1 gate1666(.O (g3245), .I (I13131));
INVX1 gate1667(.O (I13134), .I (g30));
INVX1 gate1668(.O (g3246), .I (I13134));
INVX1 gate1669(.O (I13137), .I (g33));
INVX1 gate1670(.O (g3247), .I (I13137));
INVX1 gate1671(.O (I13140), .I (g36));
INVX1 gate1672(.O (g3248), .I (I13140));
INVX1 gate1673(.O (I13143), .I (g39));
INVX1 gate1674(.O (g3249), .I (I13143));
INVX1 gate1675(.O (I13146), .I (g42));
INVX1 gate1676(.O (g3250), .I (I13146));
INVX1 gate1677(.O (I13149), .I (g45));
INVX1 gate1678(.O (g3251), .I (I13149));
INVX1 gate1679(.O (I13152), .I (g48));
INVX1 gate1680(.O (g3252), .I (I13152));
INVX1 gate1681(.O (I13155), .I (g51));
INVX1 gate1682(.O (g3253), .I (I13155));
INVX1 gate1683(.O (I13158), .I (g165));
INVX1 gate1684(.O (g3254), .I (I13158));
INVX1 gate1685(.O (I13161), .I (g308));
INVX1 gate1686(.O (g3304), .I (I13161));
INVX1 gate1687(.O (g3305), .I (g305));
INVX1 gate1688(.O (I13165), .I (g401));
INVX1 gate1689(.O (g3306), .I (I13165));
INVX1 gate1690(.O (g3337), .I (g309));
INVX1 gate1691(.O (I13169), .I (g550));
INVX1 gate1692(.O (g3338), .I (I13169));
INVX1 gate1693(.O (g3365), .I (g499));
INVX1 gate1694(.O (I13173), .I (g629));
INVX1 gate1695(.O (g3366), .I (I13173));
INVX1 gate1696(.O (I13176), .I (g630));
INVX1 gate1697(.O (g3398), .I (I13176));
INVX1 gate1698(.O (I13179), .I (g853));
INVX1 gate1699(.O (g3410), .I (I13179));
INVX1 gate1700(.O (I13182), .I (g995));
INVX1 gate1701(.O (g3460), .I (I13182));
INVX1 gate1702(.O (g3461), .I (g992));
INVX1 gate1703(.O (I13186), .I (g1088));
INVX1 gate1704(.O (g3462), .I (I13186));
INVX1 gate1705(.O (g3493), .I (g996));
INVX1 gate1706(.O (I13190), .I (g1236));
INVX1 gate1707(.O (g3494), .I (I13190));
INVX1 gate1708(.O (g3521), .I (g1186));
INVX1 gate1709(.O (I13194), .I (g1315));
INVX1 gate1710(.O (g3522), .I (I13194));
INVX1 gate1711(.O (I13197), .I (g1316));
INVX1 gate1712(.O (g3554), .I (I13197));
INVX1 gate1713(.O (I13200), .I (g1547));
INVX1 gate1714(.O (g3566), .I (I13200));
INVX1 gate1715(.O (I13203), .I (g1689));
INVX1 gate1716(.O (g3616), .I (I13203));
INVX1 gate1717(.O (g3617), .I (g1686));
INVX1 gate1718(.O (I13207), .I (g1782));
INVX1 gate1719(.O (g3618), .I (I13207));
INVX1 gate1720(.O (g3649), .I (g1690));
INVX1 gate1721(.O (I13211), .I (g1930));
INVX1 gate1722(.O (g3650), .I (I13211));
INVX1 gate1723(.O (g3677), .I (g1880));
INVX1 gate1724(.O (I13215), .I (g2009));
INVX1 gate1725(.O (g3678), .I (I13215));
INVX1 gate1726(.O (I13218), .I (g2010));
INVX1 gate1727(.O (g3710), .I (I13218));
INVX1 gate1728(.O (I13221), .I (g2241));
INVX1 gate1729(.O (g3722), .I (I13221));
INVX1 gate1730(.O (I13224), .I (g2383));
INVX1 gate1731(.O (g3772), .I (I13224));
INVX1 gate1732(.O (g3773), .I (g2380));
INVX1 gate1733(.O (I13228), .I (g2476));
INVX1 gate1734(.O (g3774), .I (I13228));
INVX1 gate1735(.O (g3805), .I (g2384));
INVX1 gate1736(.O (I13232), .I (g2624));
INVX1 gate1737(.O (g3806), .I (I13232));
INVX1 gate1738(.O (g3833), .I (g2574));
INVX1 gate1739(.O (I13236), .I (g2703));
INVX1 gate1740(.O (g3834), .I (I13236));
INVX1 gate1741(.O (I13239), .I (g2704));
INVX1 gate1742(.O (g3866), .I (I13239));
INVX1 gate1743(.O (I13242), .I (g2879));
INVX1 gate1744(.O (g3878), .I (I13242));
INVX1 gate1745(.O (g3897), .I (g2950));
INVX1 gate1746(.O (I13246), .I (g2987));
INVX1 gate1747(.O (g3900), .I (I13246));
INVX1 gate1748(.O (g3919), .I (g3080));
INVX1 gate1749(.O (g3922), .I (g150));
INVX1 gate1750(.O (g3925), .I (g155));
INVX1 gate1751(.O (g3928), .I (g157));
INVX1 gate1752(.O (g3931), .I (g171));
INVX1 gate1753(.O (g3934), .I (g176));
INVX1 gate1754(.O (g3937), .I (g178));
INVX1 gate1755(.O (g3940), .I (g408));
INVX1 gate1756(.O (g3941), .I (g455));
INVX1 gate1757(.O (g3942), .I (g699));
INVX1 gate1758(.O (g3945), .I (g726));
INVX1 gate1759(.O (g3948), .I (g835));
INVX1 gate1760(.O (g3951), .I (g840));
INVX1 gate1761(.O (g3954), .I (g842));
INVX1 gate1762(.O (g3957), .I (g856));
INVX1 gate1763(.O (g3960), .I (g861));
INVX1 gate1764(.O (g3963), .I (g863));
INVX1 gate1765(.O (g3966), .I (g1526));
INVX1 gate1766(.O (g3969), .I (g1531));
INVX1 gate1767(.O (g3972), .I (g1533));
INVX1 gate1768(.O (g3975), .I (g1552));
INVX1 gate1769(.O (g3978), .I (g1554));
INVX1 gate1770(.O (g3981), .I (g2217));
INVX1 gate1771(.O (g3984), .I (g2222));
INVX1 gate1772(.O (g3987), .I (g2224));
INVX1 gate1773(.O (g3990), .I (g2245));
INVX1 gate1774(.O (I13275), .I (g2848));
INVX1 gate1775(.O (g3993), .I (I13275));
INVX1 gate1776(.O (g3994), .I (g2848));
INVX1 gate1777(.O (g3995), .I (g3064));
INVX1 gate1778(.O (g3996), .I (g3073));
INVX1 gate1779(.O (g3997), .I (g45));
INVX1 gate1780(.O (g3998), .I (g23));
INVX1 gate1781(.O (g3999), .I (g3204));
INVX1 gate1782(.O (g4000), .I (g153));
INVX1 gate1783(.O (g4003), .I (g158));
INVX1 gate1784(.O (g4006), .I (g160));
INVX1 gate1785(.O (g4009), .I (g174));
INVX1 gate1786(.O (g4012), .I (g179));
INVX1 gate1787(.O (g4015), .I (g411));
INVX1 gate1788(.O (g4016), .I (g417));
INVX1 gate1789(.O (g4017), .I (g427));
INVX1 gate1790(.O (g4020), .I (g700));
INVX1 gate1791(.O (g4023), .I (g702));
INVX1 gate1792(.O (g4026), .I (g727));
INVX1 gate1793(.O (g4029), .I (g838));
INVX1 gate1794(.O (g4032), .I (g843));
INVX1 gate1795(.O (g4035), .I (g845));
INVX1 gate1796(.O (g4038), .I (g859));
INVX1 gate1797(.O (g4041), .I (g864));
INVX1 gate1798(.O (g4044), .I (g866));
INVX1 gate1799(.O (g4047), .I (g1095));
INVX1 gate1800(.O (g4048), .I (g1142));
INVX1 gate1801(.O (g4049), .I (g1385));
INVX1 gate1802(.O (g4052), .I (g1412));
INVX1 gate1803(.O (g4055), .I (g1529));
INVX1 gate1804(.O (g4058), .I (g1534));
INVX1 gate1805(.O (g4061), .I (g1536));
INVX1 gate1806(.O (g4064), .I (g1550));
INVX1 gate1807(.O (g4067), .I (g1555));
INVX1 gate1808(.O (g4070), .I (g1557));
INVX1 gate1809(.O (g4073), .I (g2220));
INVX1 gate1810(.O (g4076), .I (g2225));
INVX1 gate1811(.O (g4079), .I (g2227));
INVX1 gate1812(.O (g4082), .I (g2246));
INVX1 gate1813(.O (g4085), .I (g2248));
INVX1 gate1814(.O (I13316), .I (g2836));
INVX1 gate1815(.O (g4088), .I (I13316));
INVX1 gate1816(.O (g4089), .I (g2836));
INVX1 gate1817(.O (I13320), .I (g2864));
INVX1 gate1818(.O (g4090), .I (I13320));
INVX1 gate1819(.O (g4091), .I (g2864));
INVX1 gate1820(.O (g4092), .I (g3074));
INVX1 gate1821(.O (g4093), .I (g33));
INVX1 gate1822(.O (g4094), .I (g3207));
INVX1 gate1823(.O (g4095), .I (g130));
INVX1 gate1824(.O (g4098), .I (g156));
INVX1 gate1825(.O (g4101), .I (g161));
INVX1 gate1826(.O (g4104), .I (g163));
INVX1 gate1827(.O (g4107), .I (g177));
INVX1 gate1828(.O (g4110), .I (g414));
INVX1 gate1829(.O (g4111), .I (g420));
INVX1 gate1830(.O (g4112), .I (g428));
INVX1 gate1831(.O (g4115), .I (g698));
INVX1 gate1832(.O (g4118), .I (g703));
INVX1 gate1833(.O (g4121), .I (g705));
INVX1 gate1834(.O (g4124), .I (g725));
INVX1 gate1835(.O (g4127), .I (g841));
INVX1 gate1836(.O (g4130), .I (g846));
INVX1 gate1837(.O (g4133), .I (g848));
INVX1 gate1838(.O (g4136), .I (g862));
INVX1 gate1839(.O (g4139), .I (g867));
INVX1 gate1840(.O (g4142), .I (g1098));
INVX1 gate1841(.O (g4143), .I (g1104));
INVX1 gate1842(.O (g4144), .I (g1114));
INVX1 gate1843(.O (g4147), .I (g1386));
INVX1 gate1844(.O (g4150), .I (g1388));
INVX1 gate1845(.O (g4153), .I (g1413));
INVX1 gate1846(.O (g4156), .I (g1532));
INVX1 gate1847(.O (g4159), .I (g1537));
INVX1 gate1848(.O (g4162), .I (g1539));
INVX1 gate1849(.O (g4165), .I (g1553));
INVX1 gate1850(.O (g4168), .I (g1558));
INVX1 gate1851(.O (g4171), .I (g1560));
INVX1 gate1852(.O (g4174), .I (g1789));
INVX1 gate1853(.O (g4175), .I (g1836));
INVX1 gate1854(.O (g4176), .I (g2079));
INVX1 gate1855(.O (g4179), .I (g2106));
INVX1 gate1856(.O (g4182), .I (g2223));
INVX1 gate1857(.O (g4185), .I (g2228));
INVX1 gate1858(.O (g4188), .I (g2230));
INVX1 gate1859(.O (g4191), .I (g2244));
INVX1 gate1860(.O (g4194), .I (g2249));
INVX1 gate1861(.O (g4197), .I (g2251));
INVX1 gate1862(.O (I13366), .I (g2851));
INVX1 gate1863(.O (g4200), .I (I13366));
INVX1 gate1864(.O (g4201), .I (g2851));
INVX1 gate1865(.O (g4202), .I (g42));
INVX1 gate1866(.O (g4203), .I (g20));
INVX1 gate1867(.O (g4204), .I (g3188));
INVX1 gate1868(.O (g4205), .I (g131));
INVX1 gate1869(.O (g4208), .I (g133));
INVX1 gate1870(.O (g4211), .I (g159));
INVX1 gate1871(.O (g4214), .I (g164));
INVX1 gate1872(.O (g4217), .I (g354));
INVX1 gate1873(.O (g4220), .I (g423));
INVX1 gate1874(.O (g4221), .I (g426));
INVX1 gate1875(.O (g4224), .I (g429));
INVX1 gate1876(.O (g4225), .I (g701));
INVX1 gate1877(.O (g4228), .I (g706));
INVX1 gate1878(.O (g4231), .I (g708));
INVX1 gate1879(.O (g4234), .I (g818));
INVX1 gate1880(.O (g4237), .I (g844));
INVX1 gate1881(.O (g4240), .I (g849));
INVX1 gate1882(.O (g4243), .I (g851));
INVX1 gate1883(.O (g4246), .I (g865));
INVX1 gate1884(.O (g4249), .I (g1101));
INVX1 gate1885(.O (g4250), .I (g1107));
INVX1 gate1886(.O (g4251), .I (g1115));
INVX1 gate1887(.O (g4254), .I (g1384));
INVX1 gate1888(.O (g4257), .I (g1389));
INVX1 gate1889(.O (g4260), .I (g1391));
INVX1 gate1890(.O (g4263), .I (g1411));
INVX1 gate1891(.O (g4266), .I (g1535));
INVX1 gate1892(.O (g4269), .I (g1540));
INVX1 gate1893(.O (g4272), .I (g1542));
INVX1 gate1894(.O (g4275), .I (g1556));
INVX1 gate1895(.O (g4278), .I (g1561));
INVX1 gate1896(.O (g4281), .I (g1792));
INVX1 gate1897(.O (g4282), .I (g1798));
INVX1 gate1898(.O (g4283), .I (g1808));
INVX1 gate1899(.O (g4286), .I (g2080));
INVX1 gate1900(.O (g4289), .I (g2082));
INVX1 gate1901(.O (g4292), .I (g2107));
INVX1 gate1902(.O (g4295), .I (g2226));
INVX1 gate1903(.O (g4298), .I (g2231));
INVX1 gate1904(.O (g4301), .I (g2233));
INVX1 gate1905(.O (g4304), .I (g2247));
INVX1 gate1906(.O (g4307), .I (g2252));
INVX1 gate1907(.O (g4310), .I (g2254));
INVX1 gate1908(.O (g4313), .I (g2483));
INVX1 gate1909(.O (g4314), .I (g2530));
INVX1 gate1910(.O (g4315), .I (g2773));
INVX1 gate1911(.O (g4318), .I (g2800));
INVX1 gate1912(.O (I13417), .I (g2839));
INVX1 gate1913(.O (g4321), .I (I13417));
INVX1 gate1914(.O (g4322), .I (g2839));
INVX1 gate1915(.O (I13421), .I (g2867));
INVX1 gate1916(.O (g4323), .I (I13421));
INVX1 gate1917(.O (g4324), .I (g2867));
INVX1 gate1918(.O (g4325), .I (g36));
INVX1 gate1919(.O (g4326), .I (g181));
INVX1 gate1920(.O (g4329), .I (g129));
INVX1 gate1921(.O (g4332), .I (g134));
INVX1 gate1922(.O (g4335), .I (g162));
INVX1 gate1923(.O (I13430), .I (g101));
INVX1 gate1924(.O (g4338), .I (I13430));
INVX1 gate1925(.O (I13433), .I (g105));
INVX1 gate1926(.O (g4339), .I (I13433));
INVX1 gate1927(.O (g4340), .I (g343));
INVX1 gate1928(.O (g4343), .I (g369));
INVX1 gate1929(.O (g4346), .I (g432));
INVX1 gate1930(.O (g4347), .I (g438));
INVX1 gate1931(.O (g4348), .I (g704));
INVX1 gate1932(.O (g4351), .I (g709));
INVX1 gate1933(.O (g4354), .I (g711));
INVX1 gate1934(.O (g4357), .I (g729));
INVX1 gate1935(.O (g4360), .I (g819));
INVX1 gate1936(.O (g4363), .I (g821));
INVX1 gate1937(.O (g4366), .I (g847));
INVX1 gate1938(.O (g4369), .I (g852));
INVX1 gate1939(.O (g4372), .I (g1041));
INVX1 gate1940(.O (g4375), .I (g1110));
INVX1 gate1941(.O (g4376), .I (g1113));
INVX1 gate1942(.O (g4379), .I (g1116));
INVX1 gate1943(.O (g4380), .I (g1387));
INVX1 gate1944(.O (g4383), .I (g1392));
INVX1 gate1945(.O (g4386), .I (g1394));
INVX1 gate1946(.O (g4389), .I (g1512));
INVX1 gate1947(.O (g4392), .I (g1538));
INVX1 gate1948(.O (g4395), .I (g1543));
INVX1 gate1949(.O (g4398), .I (g1545));
INVX1 gate1950(.O (g4401), .I (g1559));
INVX1 gate1951(.O (g4404), .I (g1795));
INVX1 gate1952(.O (g4405), .I (g1801));
INVX1 gate1953(.O (g4406), .I (g1809));
INVX1 gate1954(.O (g4409), .I (g2078));
INVX1 gate1955(.O (g4412), .I (g2083));
INVX1 gate1956(.O (g4415), .I (g2085));
INVX1 gate1957(.O (g4418), .I (g2105));
INVX1 gate1958(.O (g4421), .I (g2229));
INVX1 gate1959(.O (g4424), .I (g2234));
INVX1 gate1960(.O (g4427), .I (g2236));
INVX1 gate1961(.O (g4430), .I (g2250));
INVX1 gate1962(.O (g4433), .I (g2255));
INVX1 gate1963(.O (g4436), .I (g2486));
INVX1 gate1964(.O (g4437), .I (g2492));
INVX1 gate1965(.O (g4438), .I (g2502));
INVX1 gate1966(.O (g4441), .I (g2774));
INVX1 gate1967(.O (g4444), .I (g2776));
INVX1 gate1968(.O (g4447), .I (g2801));
INVX1 gate1969(.O (I13478), .I (g2854));
INVX1 gate1970(.O (g4450), .I (I13478));
INVX1 gate1971(.O (g4451), .I (g2854));
INVX1 gate1972(.O (g4452), .I (g17));
INVX1 gate1973(.O (g4453), .I (g132));
INVX1 gate1974(.O (g4456), .I (g309));
INVX1 gate1975(.O (g4465), .I (g346));
INVX1 gate1976(.O (g4468), .I (g358));
INVX1 gate1977(.O (g4471), .I (g384));
INVX1 gate1978(.O (g4474), .I (g435));
INVX1 gate1979(.O (g4475), .I (g441));
INVX1 gate1980(.O (g4476), .I (g576));
INVX1 gate1981(.O (g4479), .I (g587));
INVX1 gate1982(.O (g4480), .I (g707));
INVX1 gate1983(.O (g4483), .I (g712));
INVX1 gate1984(.O (g4486), .I (g714));
INVX1 gate1985(.O (g4489), .I (g730));
INVX1 gate1986(.O (g4492), .I (g732));
INVX1 gate1987(.O (g4495), .I (g869));
INVX1 gate1988(.O (g4498), .I (g817));
INVX1 gate1989(.O (g4501), .I (g822));
INVX1 gate1990(.O (g4504), .I (g850));
INVX1 gate1991(.O (I13501), .I (g789));
INVX1 gate1992(.O (g4507), .I (I13501));
INVX1 gate1993(.O (I13504), .I (g793));
INVX1 gate1994(.O (g4508), .I (I13504));
INVX1 gate1995(.O (g4509), .I (g1030));
INVX1 gate1996(.O (g4512), .I (g1056));
INVX1 gate1997(.O (g4515), .I (g1119));
INVX1 gate1998(.O (g4516), .I (g1125));
INVX1 gate1999(.O (g4517), .I (g1390));
INVX1 gate2000(.O (g4520), .I (g1395));
INVX1 gate2001(.O (g4523), .I (g1397));
INVX1 gate2002(.O (g4526), .I (g1415));
INVX1 gate2003(.O (g4529), .I (g1513));
INVX1 gate2004(.O (g4532), .I (g1515));
INVX1 gate2005(.O (g4535), .I (g1541));
INVX1 gate2006(.O (g4538), .I (g1546));
INVX1 gate2007(.O (g4541), .I (g1735));
INVX1 gate2008(.O (g4544), .I (g1804));
INVX1 gate2009(.O (g4545), .I (g1807));
INVX1 gate2010(.O (g4548), .I (g1810));
INVX1 gate2011(.O (g4549), .I (g2081));
INVX1 gate2012(.O (g4552), .I (g2086));
INVX1 gate2013(.O (g4555), .I (g2088));
INVX1 gate2014(.O (g4558), .I (g2206));
INVX1 gate2015(.O (g4561), .I (g2232));
INVX1 gate2016(.O (g4564), .I (g2237));
INVX1 gate2017(.O (g4567), .I (g2239));
INVX1 gate2018(.O (g4570), .I (g2253));
INVX1 gate2019(.O (g4573), .I (g2489));
INVX1 gate2020(.O (g4574), .I (g2495));
INVX1 gate2021(.O (g4575), .I (g2503));
INVX1 gate2022(.O (g4578), .I (g2772));
INVX1 gate2023(.O (g4581), .I (g2777));
INVX1 gate2024(.O (g4584), .I (g2779));
INVX1 gate2025(.O (g4587), .I (g2799));
INVX1 gate2026(.O (I13538), .I (g2870));
INVX1 gate2027(.O (g4590), .I (I13538));
INVX1 gate2028(.O (g4591), .I (g2870));
INVX1 gate2029(.O (g4592), .I (g361));
INVX1 gate2030(.O (g4595), .I (g373));
INVX1 gate2031(.O (g4598), .I (g398));
INVX1 gate2032(.O (g4601), .I (g444));
INVX1 gate2033(.O (g4602), .I (g525));
INVX1 gate2034(.O (g4603), .I (g577));
INVX1 gate2035(.O (g4606), .I (g579));
INVX1 gate2036(.O (g4609), .I (g590));
INVX1 gate2037(.O (g4610), .I (g596));
INVX1 gate2038(.O (g4611), .I (g710));
INVX1 gate2039(.O (g4614), .I (g715));
INVX1 gate2040(.O (g4617), .I (g717));
INVX1 gate2041(.O (g4620), .I (g728));
INVX1 gate2042(.O (g4623), .I (g733));
INVX1 gate2043(.O (g4626), .I (g735));
INVX1 gate2044(.O (g4629), .I (g820));
INVX1 gate2045(.O (g4632), .I (g996));
INVX1 gate2046(.O (g4641), .I (g1033));
INVX1 gate2047(.O (g4644), .I (g1045));
INVX1 gate2048(.O (g4647), .I (g1071));
INVX1 gate2049(.O (g4650), .I (g1122));
INVX1 gate2050(.O (g4651), .I (g1128));
INVX1 gate2051(.O (g4652), .I (g1262));
INVX1 gate2052(.O (g4655), .I (g1273));
INVX1 gate2053(.O (g4656), .I (g1393));
INVX1 gate2054(.O (g4659), .I (g1398));
INVX1 gate2055(.O (g4662), .I (g1400));
INVX1 gate2056(.O (g4665), .I (g1416));
INVX1 gate2057(.O (g4668), .I (g1418));
INVX1 gate2058(.O (g4671), .I (g1563));
INVX1 gate2059(.O (g4674), .I (g1511));
INVX1 gate2060(.O (g4677), .I (g1516));
INVX1 gate2061(.O (g4680), .I (g1544));
INVX1 gate2062(.O (I13575), .I (g1476));
INVX1 gate2063(.O (g4683), .I (I13575));
INVX1 gate2064(.O (I13578), .I (g1481));
INVX1 gate2065(.O (g4684), .I (I13578));
INVX1 gate2066(.O (g4685), .I (g1724));
INVX1 gate2067(.O (g4688), .I (g1750));
INVX1 gate2068(.O (g4691), .I (g1813));
INVX1 gate2069(.O (g4692), .I (g1819));
INVX1 gate2070(.O (g4693), .I (g2084));
INVX1 gate2071(.O (g4696), .I (g2089));
INVX1 gate2072(.O (g4699), .I (g2091));
INVX1 gate2073(.O (g4702), .I (g2109));
INVX1 gate2074(.O (g4705), .I (g2207));
INVX1 gate2075(.O (g4708), .I (g2209));
INVX1 gate2076(.O (g4711), .I (g2235));
INVX1 gate2077(.O (g4714), .I (g2240));
INVX1 gate2078(.O (g4717), .I (g2429));
INVX1 gate2079(.O (g4720), .I (g2498));
INVX1 gate2080(.O (g4721), .I (g2501));
INVX1 gate2081(.O (g4724), .I (g2504));
INVX1 gate2082(.O (g4725), .I (g2775));
INVX1 gate2083(.O (g4728), .I (g2780));
INVX1 gate2084(.O (g4731), .I (g2782));
INVX1 gate2085(.O (g4734), .I (g11));
INVX1 gate2086(.O (I13601), .I (g121));
INVX1 gate2087(.O (g4735), .I (I13601));
INVX1 gate2088(.O (I13604), .I (g125));
INVX1 gate2089(.O (g4736), .I (I13604));
INVX1 gate2090(.O (g4737), .I (g376));
INVX1 gate2091(.O (g4740), .I (g388));
INVX1 gate2092(.O (g4743), .I (g575));
INVX1 gate2093(.O (g4746), .I (g580));
INVX1 gate2094(.O (g4749), .I (g582));
INVX1 gate2095(.O (g4752), .I (g593));
INVX1 gate2096(.O (g4753), .I (g599));
INVX1 gate2097(.O (g4754), .I (g713));
INVX1 gate2098(.O (g4757), .I (g718));
INVX1 gate2099(.O (g4760), .I (g720));
INVX1 gate2100(.O (g4763), .I (g731));
INVX1 gate2101(.O (g4766), .I (g736));
INVX1 gate2102(.O (g4769), .I (g1048));
INVX1 gate2103(.O (g4772), .I (g1060));
INVX1 gate2104(.O (g4775), .I (g1085));
INVX1 gate2105(.O (g4778), .I (g1131));
INVX1 gate2106(.O (g4779), .I (g1211));
INVX1 gate2107(.O (g4780), .I (g1263));
INVX1 gate2108(.O (g4783), .I (g1265));
INVX1 gate2109(.O (g4786), .I (g1276));
INVX1 gate2110(.O (g4787), .I (g1282));
INVX1 gate2111(.O (g4788), .I (g1396));
INVX1 gate2112(.O (g4791), .I (g1401));
INVX1 gate2113(.O (g4794), .I (g1403));
INVX1 gate2114(.O (g4797), .I (g1414));
INVX1 gate2115(.O (g4800), .I (g1419));
INVX1 gate2116(.O (g4803), .I (g1421));
INVX1 gate2117(.O (g4806), .I (g1514));
INVX1 gate2118(.O (g4809), .I (g1690));
INVX1 gate2119(.O (g4818), .I (g1727));
INVX1 gate2120(.O (g4821), .I (g1739));
INVX1 gate2121(.O (g4824), .I (g1765));
INVX1 gate2122(.O (g4827), .I (g1816));
INVX1 gate2123(.O (g4828), .I (g1822));
INVX1 gate2124(.O (g4829), .I (g1956));
INVX1 gate2125(.O (g4832), .I (g1967));
INVX1 gate2126(.O (g4833), .I (g2087));
INVX1 gate2127(.O (g4836), .I (g2092));
INVX1 gate2128(.O (g4839), .I (g2094));
INVX1 gate2129(.O (g4842), .I (g2110));
INVX1 gate2130(.O (g4845), .I (g2112));
INVX1 gate2131(.O (g4848), .I (g2257));
INVX1 gate2132(.O (g4851), .I (g2205));
INVX1 gate2133(.O (g4854), .I (g2210));
INVX1 gate2134(.O (g4857), .I (g2238));
INVX1 gate2135(.O (I13652), .I (g2170));
INVX1 gate2136(.O (g4860), .I (I13652));
INVX1 gate2137(.O (I13655), .I (g2175));
INVX1 gate2138(.O (g4861), .I (I13655));
INVX1 gate2139(.O (g4862), .I (g2418));
INVX1 gate2140(.O (g4865), .I (g2444));
INVX1 gate2141(.O (g4868), .I (g2507));
INVX1 gate2142(.O (g4869), .I (g2513));
INVX1 gate2143(.O (g4870), .I (g2778));
INVX1 gate2144(.O (g4873), .I (g2783));
INVX1 gate2145(.O (g4876), .I (g2785));
INVX1 gate2146(.O (g4879), .I (g2803));
INVX1 gate2147(.O (g4882), .I (g391));
INVX1 gate2148(.O (g4885), .I (g448));
INVX1 gate2149(.O (g4888), .I (g578));
INVX1 gate2150(.O (g4891), .I (g583));
INVX1 gate2151(.O (g4894), .I (g585));
INVX1 gate2152(.O (g4897), .I (g602));
INVX1 gate2153(.O (g4898), .I (g605));
INVX1 gate2154(.O (g4899), .I (g716));
INVX1 gate2155(.O (g4902), .I (g721));
INVX1 gate2156(.O (g4905), .I (g723));
INVX1 gate2157(.O (g4908), .I (g734));
INVX1 gate2158(.O (I13677), .I (g809));
INVX1 gate2159(.O (g4911), .I (I13677));
INVX1 gate2160(.O (I13680), .I (g813));
INVX1 gate2161(.O (g4912), .I (I13680));
INVX1 gate2162(.O (g4913), .I (g1063));
INVX1 gate2163(.O (g4916), .I (g1075));
INVX1 gate2164(.O (g4919), .I (g1261));
INVX1 gate2165(.O (g4922), .I (g1266));
INVX1 gate2166(.O (g4925), .I (g1268));
INVX1 gate2167(.O (g4928), .I (g1279));
INVX1 gate2168(.O (g4929), .I (g1285));
INVX1 gate2169(.O (g4930), .I (g1399));
INVX1 gate2170(.O (g4933), .I (g1404));
INVX1 gate2171(.O (g4936), .I (g1406));
INVX1 gate2172(.O (g4939), .I (g1417));
INVX1 gate2173(.O (g4942), .I (g1422));
INVX1 gate2174(.O (g4945), .I (g1742));
INVX1 gate2175(.O (g4948), .I (g1754));
INVX1 gate2176(.O (g4951), .I (g1779));
INVX1 gate2177(.O (g4954), .I (g1825));
INVX1 gate2178(.O (g4955), .I (g1905));
INVX1 gate2179(.O (g4956), .I (g1957));
INVX1 gate2180(.O (g4959), .I (g1959));
INVX1 gate2181(.O (g4962), .I (g1970));
INVX1 gate2182(.O (g4963), .I (g1976));
INVX1 gate2183(.O (g4964), .I (g2090));
INVX1 gate2184(.O (g4967), .I (g2095));
INVX1 gate2185(.O (g4970), .I (g2097));
INVX1 gate2186(.O (g4973), .I (g2108));
INVX1 gate2187(.O (g4976), .I (g2113));
INVX1 gate2188(.O (g4979), .I (g2115));
INVX1 gate2189(.O (g4982), .I (g2208));
INVX1 gate2190(.O (g4985), .I (g2384));
INVX1 gate2191(.O (g4994), .I (g2421));
INVX1 gate2192(.O (g4997), .I (g2433));
INVX1 gate2193(.O (g5000), .I (g2459));
INVX1 gate2194(.O (g5003), .I (g2510));
INVX1 gate2195(.O (g5004), .I (g2516));
INVX1 gate2196(.O (g5005), .I (g2650));
INVX1 gate2197(.O (g5008), .I (g2661));
INVX1 gate2198(.O (g5009), .I (g2781));
INVX1 gate2199(.O (g5012), .I (g2786));
INVX1 gate2200(.O (g5015), .I (g2788));
INVX1 gate2201(.O (g5018), .I (g2804));
INVX1 gate2202(.O (g5021), .I (g2806));
INVX1 gate2203(.O (g5024), .I (g449));
INVX1 gate2204(.O (g5027), .I (g581));
INVX1 gate2205(.O (g5030), .I (g586));
INVX1 gate2206(.O (g5033), .I (g608));
INVX1 gate2207(.O (g5034), .I (g614));
INVX1 gate2208(.O (g5035), .I (g719));
INVX1 gate2209(.O (g5038), .I (g724));
INVX1 gate2210(.O (g5041), .I (g1078));
INVX1 gate2211(.O (g5044), .I (g1135));
INVX1 gate2212(.O (g5047), .I (g1264));
INVX1 gate2213(.O (g5050), .I (g1269));
INVX1 gate2214(.O (g5053), .I (g1271));
INVX1 gate2215(.O (g5056), .I (g1288));
INVX1 gate2216(.O (g5057), .I (g1291));
INVX1 gate2217(.O (g5058), .I (g1402));
INVX1 gate2218(.O (g5061), .I (g1407));
INVX1 gate2219(.O (g5064), .I (g1409));
INVX1 gate2220(.O (g5067), .I (g1420));
INVX1 gate2221(.O (I13742), .I (g1501));
INVX1 gate2222(.O (g5070), .I (I13742));
INVX1 gate2223(.O (I13745), .I (g1506));
INVX1 gate2224(.O (g5071), .I (I13745));
INVX1 gate2225(.O (g5072), .I (g1757));
INVX1 gate2226(.O (g5075), .I (g1769));
INVX1 gate2227(.O (g5078), .I (g1955));
INVX1 gate2228(.O (g5081), .I (g1960));
INVX1 gate2229(.O (g5084), .I (g1962));
INVX1 gate2230(.O (g5087), .I (g1973));
INVX1 gate2231(.O (g5088), .I (g1979));
INVX1 gate2232(.O (g5089), .I (g2093));
INVX1 gate2233(.O (g5092), .I (g2098));
INVX1 gate2234(.O (g5095), .I (g2100));
INVX1 gate2235(.O (g5098), .I (g2111));
INVX1 gate2236(.O (g5101), .I (g2116));
INVX1 gate2237(.O (g5104), .I (g2436));
INVX1 gate2238(.O (g5107), .I (g2448));
INVX1 gate2239(.O (g5110), .I (g2473));
INVX1 gate2240(.O (g5113), .I (g2519));
INVX1 gate2241(.O (g5114), .I (g2599));
INVX1 gate2242(.O (g5115), .I (g2651));
INVX1 gate2243(.O (g5118), .I (g2653));
INVX1 gate2244(.O (g5121), .I (g2664));
INVX1 gate2245(.O (g5122), .I (g2670));
INVX1 gate2246(.O (g5123), .I (g2784));
INVX1 gate2247(.O (g5126), .I (g2789));
INVX1 gate2248(.O (g5129), .I (g2791));
INVX1 gate2249(.O (g5132), .I (g2802));
INVX1 gate2250(.O (g5135), .I (g2807));
INVX1 gate2251(.O (g5138), .I (g2809));
INVX1 gate2252(.O (I13775), .I (g109));
INVX1 gate2253(.O (g5141), .I (I13775));
INVX1 gate2254(.O (g5142), .I (g447));
INVX1 gate2255(.O (g5145), .I (g584));
INVX1 gate2256(.O (g5148), .I (g611));
INVX1 gate2257(.O (g5149), .I (g617));
INVX1 gate2258(.O (g5150), .I (g722));
INVX1 gate2259(.O (g5153), .I (g1136));
INVX1 gate2260(.O (g5156), .I (g1267));
INVX1 gate2261(.O (g5159), .I (g1272));
INVX1 gate2262(.O (g5162), .I (g1294));
INVX1 gate2263(.O (g5163), .I (g1300));
INVX1 gate2264(.O (g5164), .I (g1405));
INVX1 gate2265(.O (g5167), .I (g1410));
INVX1 gate2266(.O (g5170), .I (g1772));
INVX1 gate2267(.O (g5173), .I (g1829));
INVX1 gate2268(.O (g5176), .I (g1958));
INVX1 gate2269(.O (g5179), .I (g1963));
INVX1 gate2270(.O (g5182), .I (g1965));
INVX1 gate2271(.O (g5185), .I (g1982));
INVX1 gate2272(.O (g5186), .I (g1985));
INVX1 gate2273(.O (g5187), .I (g2096));
INVX1 gate2274(.O (g5190), .I (g2101));
INVX1 gate2275(.O (g5193), .I (g2103));
INVX1 gate2276(.O (g5196), .I (g2114));
INVX1 gate2277(.O (I13801), .I (g2195));
INVX1 gate2278(.O (g5199), .I (I13801));
INVX1 gate2279(.O (I13804), .I (g2200));
INVX1 gate2280(.O (g5200), .I (I13804));
INVX1 gate2281(.O (g5201), .I (g2451));
INVX1 gate2282(.O (g5204), .I (g2463));
INVX1 gate2283(.O (g5207), .I (g2649));
INVX1 gate2284(.O (g5210), .I (g2654));
INVX1 gate2285(.O (g5213), .I (g2656));
INVX1 gate2286(.O (g5216), .I (g2667));
INVX1 gate2287(.O (g5217), .I (g2673));
INVX1 gate2288(.O (g5218), .I (g2787));
INVX1 gate2289(.O (g5221), .I (g2792));
INVX1 gate2290(.O (g5224), .I (g2794));
INVX1 gate2291(.O (g5227), .I (g2805));
INVX1 gate2292(.O (g5230), .I (g2810));
INVX1 gate2293(.O (g5233), .I (g620));
INVX1 gate2294(.O (I13820), .I (g797));
INVX1 gate2295(.O (g5234), .I (I13820));
INVX1 gate2296(.O (g5235), .I (g1134));
INVX1 gate2297(.O (g5238), .I (g1270));
INVX1 gate2298(.O (g5241), .I (g1297));
INVX1 gate2299(.O (g5242), .I (g1303));
INVX1 gate2300(.O (g5243), .I (g1408));
INVX1 gate2301(.O (g5246), .I (g1830));
INVX1 gate2302(.O (g5249), .I (g1961));
INVX1 gate2303(.O (g5252), .I (g1966));
INVX1 gate2304(.O (g5255), .I (g1988));
INVX1 gate2305(.O (g5256), .I (g1994));
INVX1 gate2306(.O (g5257), .I (g2099));
INVX1 gate2307(.O (g5260), .I (g2104));
INVX1 gate2308(.O (g5263), .I (g2466));
INVX1 gate2309(.O (g5266), .I (g2523));
INVX1 gate2310(.O (g5269), .I (g2652));
INVX1 gate2311(.O (g5272), .I (g2657));
INVX1 gate2312(.O (g5275), .I (g2659));
INVX1 gate2313(.O (g5278), .I (g2676));
INVX1 gate2314(.O (g5279), .I (g2679));
INVX1 gate2315(.O (g5280), .I (g2790));
INVX1 gate2316(.O (g5283), .I (g2795));
INVX1 gate2317(.O (g5286), .I (g2797));
INVX1 gate2318(.O (g5289), .I (g2808));
INVX1 gate2319(.O (g5292), .I (g2857));
INVX1 gate2320(.O (g5293), .I (g738));
INVX1 gate2321(.O (g5296), .I (g1306));
INVX1 gate2322(.O (I13849), .I (g1486));
INVX1 gate2323(.O (g5297), .I (I13849));
INVX1 gate2324(.O (g5298), .I (g1828));
INVX1 gate2325(.O (g5301), .I (g1964));
INVX1 gate2326(.O (g5304), .I (g1991));
INVX1 gate2327(.O (g5305), .I (g1997));
INVX1 gate2328(.O (g5306), .I (g2102));
INVX1 gate2329(.O (g5309), .I (g2524));
INVX1 gate2330(.O (g5312), .I (g2655));
INVX1 gate2331(.O (g5315), .I (g2660));
INVX1 gate2332(.O (g5318), .I (g2682));
INVX1 gate2333(.O (g5319), .I (g2688));
INVX1 gate2334(.O (g5320), .I (g2793));
INVX1 gate2335(.O (g5323), .I (g2798));
INVX1 gate2336(.O (g5326), .I (g2873));
INVX1 gate2337(.O (g5327), .I (g739));
INVX1 gate2338(.O (g5330), .I (g1424));
INVX1 gate2339(.O (g5333), .I (g2000));
INVX1 gate2340(.O (I13868), .I (g2180));
INVX1 gate2341(.O (g5334), .I (I13868));
INVX1 gate2342(.O (g5335), .I (g2522));
INVX1 gate2343(.O (g5338), .I (g2658));
INVX1 gate2344(.O (g5341), .I (g2685));
INVX1 gate2345(.O (g5342), .I (g2691));
INVX1 gate2346(.O (g5343), .I (g2796));
INVX1 gate2347(.O (g5346), .I (g3106));
INVX1 gate2348(.O (g5349), .I (g2877));
INVX1 gate2349(.O (g5352), .I (g737));
INVX1 gate2350(.O (g5355), .I (g1425));
INVX1 gate2351(.O (g5358), .I (g2118));
INVX1 gate2352(.O (g5361), .I (g2694));
INVX1 gate2353(.O (g5362), .I (g2817));
INVX1 gate2354(.O (g5363), .I (g3107));
INVX1 gate2355(.O (g5366), .I (g2878));
INVX1 gate2356(.O (g5369), .I (g1423));
INVX1 gate2357(.O (g5372), .I (g2119));
INVX1 gate2358(.O (g5375), .I (g2812));
INVX1 gate2359(.O (g5378), .I (g2933));
INVX1 gate2360(.O (g5379), .I (g3108));
INVX1 gate2361(.O (g5382), .I (g2117));
INVX1 gate2362(.O (g5385), .I (g2813));
INVX1 gate2363(.O (I13892), .I (g3040));
INVX1 gate2364(.O (g5388), .I (I13892));
INVX1 gate2365(.O (g5389), .I (g3040));
INVX1 gate2366(.O (I13896), .I (g343));
INVX1 gate2367(.O (g5390), .I (I13896));
INVX1 gate2368(.O (g5391), .I (g2811));
INVX1 gate2369(.O (g5394), .I (g3054));
INVX1 gate2370(.O (I13901), .I (g346));
INVX1 gate2371(.O (g5395), .I (I13901));
INVX1 gate2372(.O (I13904), .I (g358));
INVX1 gate2373(.O (g5396), .I (I13904));
INVX1 gate2374(.O (I13907), .I (g1030));
INVX1 gate2375(.O (g5397), .I (I13907));
INVX1 gate2376(.O (I13910), .I (g361));
INVX1 gate2377(.O (g5398), .I (I13910));
INVX1 gate2378(.O (I13913), .I (g373));
INVX1 gate2379(.O (g5399), .I (I13913));
INVX1 gate2380(.O (I13916), .I (g1033));
INVX1 gate2381(.O (g5400), .I (I13916));
INVX1 gate2382(.O (I13919), .I (g1045));
INVX1 gate2383(.O (g5401), .I (I13919));
INVX1 gate2384(.O (I13922), .I (g1724));
INVX1 gate2385(.O (g5402), .I (I13922));
INVX1 gate2386(.O (I13925), .I (g376));
INVX1 gate2387(.O (g5403), .I (I13925));
INVX1 gate2388(.O (I13928), .I (g388));
INVX1 gate2389(.O (g5404), .I (I13928));
INVX1 gate2390(.O (I13931), .I (g1048));
INVX1 gate2391(.O (g5405), .I (I13931));
INVX1 gate2392(.O (I13934), .I (g1060));
INVX1 gate2393(.O (g5406), .I (I13934));
INVX1 gate2394(.O (I13937), .I (g1727));
INVX1 gate2395(.O (g5407), .I (I13937));
INVX1 gate2396(.O (I13940), .I (g1739));
INVX1 gate2397(.O (g5408), .I (I13940));
INVX1 gate2398(.O (I13943), .I (g2418));
INVX1 gate2399(.O (g5409), .I (I13943));
INVX1 gate2400(.O (g5410), .I (g3079));
INVX1 gate2401(.O (I13947), .I (g391));
INVX1 gate2402(.O (g5411), .I (I13947));
INVX1 gate2403(.O (I13950), .I (g1063));
INVX1 gate2404(.O (g5412), .I (I13950));
INVX1 gate2405(.O (I13953), .I (g1075));
INVX1 gate2406(.O (g5413), .I (I13953));
INVX1 gate2407(.O (I13956), .I (g1742));
INVX1 gate2408(.O (g5414), .I (I13956));
INVX1 gate2409(.O (I13959), .I (g1754));
INVX1 gate2410(.O (g5415), .I (I13959));
INVX1 gate2411(.O (I13962), .I (g2421));
INVX1 gate2412(.O (g5416), .I (I13962));
INVX1 gate2413(.O (I13965), .I (g2433));
INVX1 gate2414(.O (g5417), .I (I13965));
INVX1 gate2415(.O (I13968), .I (g1078));
INVX1 gate2416(.O (g5418), .I (I13968));
INVX1 gate2417(.O (I13971), .I (g1757));
INVX1 gate2418(.O (g5419), .I (I13971));
INVX1 gate2419(.O (I13974), .I (g1769));
INVX1 gate2420(.O (g5420), .I (I13974));
INVX1 gate2421(.O (I13977), .I (g2436));
INVX1 gate2422(.O (g5421), .I (I13977));
INVX1 gate2423(.O (I13980), .I (g2448));
INVX1 gate2424(.O (g5422), .I (I13980));
INVX1 gate2425(.O (g5423), .I (g2879));
INVX1 gate2426(.O (I13984), .I (g1772));
INVX1 gate2427(.O (g5424), .I (I13984));
INVX1 gate2428(.O (I13987), .I (g2451));
INVX1 gate2429(.O (g5425), .I (I13987));
INVX1 gate2430(.O (I13990), .I (g2463));
INVX1 gate2431(.O (g5426), .I (I13990));
INVX1 gate2432(.O (I13993), .I (g2466));
INVX1 gate2433(.O (g5427), .I (I13993));
INVX1 gate2434(.O (g5428), .I (g3210));
INVX1 gate2435(.O (g5431), .I (g3211));
INVX1 gate2436(.O (g5434), .I (g3084));
INVX1 gate2437(.O (I13999), .I (g276));
INVX1 gate2438(.O (g5437), .I (I13999));
INVX1 gate2439(.O (I14002), .I (g276));
INVX1 gate2440(.O (g5438), .I (I14002));
INVX1 gate2441(.O (g5469), .I (g3085));
INVX1 gate2442(.O (I14006), .I (g963));
INVX1 gate2443(.O (g5472), .I (I14006));
INVX1 gate2444(.O (I14009), .I (g963));
INVX1 gate2445(.O (g5473), .I (I14009));
INVX1 gate2446(.O (g5504), .I (g3086));
INVX1 gate2447(.O (g5507), .I (g3155));
INVX1 gate2448(.O (I14014), .I (g499));
INVX1 gate2449(.O (g5508), .I (I14014));
INVX1 gate2450(.O (I14017), .I (g1657));
INVX1 gate2451(.O (g5511), .I (I14017));
INVX1 gate2452(.O (I14020), .I (g1657));
INVX1 gate2453(.O (g5512), .I (I14020));
INVX1 gate2454(.O (g5543), .I (g3087));
INVX1 gate2455(.O (g5546), .I (g3164));
INVX1 gate2456(.O (g5547), .I (g101));
INVX1 gate2457(.O (g5548), .I (g105));
INVX1 gate2458(.O (I14027), .I (g182));
INVX1 gate2459(.O (g5549), .I (I14027));
INVX1 gate2460(.O (I14030), .I (g182));
INVX1 gate2461(.O (g5550), .I (I14030));
INVX1 gate2462(.O (g5551), .I (g514));
INVX1 gate2463(.O (I14034), .I (g1186));
INVX1 gate2464(.O (g5552), .I (I14034));
INVX1 gate2465(.O (I14037), .I (g2351));
INVX1 gate2466(.O (g5555), .I (I14037));
INVX1 gate2467(.O (I14040), .I (g2351));
INVX1 gate2468(.O (g5556), .I (I14040));
INVX1 gate2469(.O (g5587), .I (g3091));
INVX1 gate2470(.O (g5590), .I (g3158));
INVX1 gate2471(.O (g5591), .I (g3173));
INVX1 gate2472(.O (g5592), .I (g515));
INVX1 gate2473(.O (g5593), .I (g789));
INVX1 gate2474(.O (g5594), .I (g793));
INVX1 gate2475(.O (I14049), .I (g870));
INVX1 gate2476(.O (g5595), .I (I14049));
INVX1 gate2477(.O (I14052), .I (g870));
INVX1 gate2478(.O (g5596), .I (I14052));
INVX1 gate2479(.O (g5597), .I (g1200));
INVX1 gate2480(.O (I14056), .I (g1880));
INVX1 gate2481(.O (g5598), .I (I14056));
INVX1 gate2482(.O (g5601), .I (g3092));
INVX1 gate2483(.O (g5604), .I (g3167));
INVX1 gate2484(.O (g5605), .I (g3182));
INVX1 gate2485(.O (g5606), .I (g79));
INVX1 gate2486(.O (g5609), .I (g1201));
INVX1 gate2487(.O (g5610), .I (g1476));
INVX1 gate2488(.O (g5611), .I (g1481));
INVX1 gate2489(.O (I14066), .I (g1564));
INVX1 gate2490(.O (g5612), .I (I14066));
INVX1 gate2491(.O (I14069), .I (g1564));
INVX1 gate2492(.O (g5613), .I (I14069));
INVX1 gate2493(.O (g5614), .I (g1894));
INVX1 gate2494(.O (I14073), .I (g2574));
INVX1 gate2495(.O (g5615), .I (I14073));
INVX1 gate2496(.O (g5618), .I (g3093));
INVX1 gate2497(.O (g5621), .I (g3161));
INVX1 gate2498(.O (g5622), .I (g3176));
INVX1 gate2499(.O (g5623), .I (g70));
INVX1 gate2500(.O (g5626), .I (g121));
INVX1 gate2501(.O (g5627), .I (g125));
INVX1 gate2502(.O (g5628), .I (g300));
INVX1 gate2503(.O (I14083), .I (g325));
INVX1 gate2504(.O (g5629), .I (I14083));
INVX1 gate2505(.O (g5631), .I (g767));
INVX1 gate2506(.O (g5634), .I (g1895));
INVX1 gate2507(.O (g5635), .I (g2170));
INVX1 gate2508(.O (g5636), .I (g2175));
INVX1 gate2509(.O (I14091), .I (g2258));
INVX1 gate2510(.O (g5637), .I (I14091));
INVX1 gate2511(.O (I14094), .I (g2258));
INVX1 gate2512(.O (g5638), .I (I14094));
INVX1 gate2513(.O (g5639), .I (g2588));
INVX1 gate2514(.O (g5640), .I (g3170));
INVX1 gate2515(.O (g5641), .I (g3185));
INVX1 gate2516(.O (g5642), .I (g61));
INVX1 gate2517(.O (g5645), .I (g101));
INVX1 gate2518(.O (g5646), .I (g213));
INVX1 gate2519(.O (g5647), .I (g301));
INVX1 gate2520(.O (I14104), .I (g331));
INVX1 gate2521(.O (g5648), .I (I14104));
INVX1 gate2522(.O (g5651), .I (g758));
INVX1 gate2523(.O (g5654), .I (g809));
INVX1 gate2524(.O (g5655), .I (g813));
INVX1 gate2525(.O (g5656), .I (g987));
INVX1 gate2526(.O (I14113), .I (g1012));
INVX1 gate2527(.O (g5657), .I (I14113));
INVX1 gate2528(.O (g5659), .I (g1453));
INVX1 gate2529(.O (g5662), .I (g2589));
INVX1 gate2530(.O (g5663), .I (g3179));
INVX1 gate2531(.O (g5664), .I (g65));
INVX1 gate2532(.O (g5665), .I (g105));
INVX1 gate2533(.O (g5666), .I (g216));
INVX1 gate2534(.O (g5667), .I (g222));
INVX1 gate2535(.O (g5668), .I (g299));
INVX1 gate2536(.O (g5675), .I (g302));
INVX1 gate2537(.O (g5679), .I (g506));
INVX1 gate2538(.O (g5680), .I (g749));
INVX1 gate2539(.O (g5683), .I (g789));
INVX1 gate2540(.O (g5684), .I (g900));
INVX1 gate2541(.O (g5685), .I (g988));
INVX1 gate2542(.O (I14134), .I (g1018));
INVX1 gate2543(.O (g5686), .I (I14134));
INVX1 gate2544(.O (g5689), .I (g1444));
INVX1 gate2545(.O (g5692), .I (g1501));
INVX1 gate2546(.O (g5693), .I (g1506));
INVX1 gate2547(.O (g5694), .I (g1681));
INVX1 gate2548(.O (I14143), .I (g1706));
INVX1 gate2549(.O (g5695), .I (I14143));
INVX1 gate2550(.O (g5697), .I (g2147));
INVX1 gate2551(.O (g5700), .I (g3088));
INVX1 gate2552(.O (I14149), .I (g3231));
INVX1 gate2553(.O (g5701), .I (I14149));
INVX1 gate2554(.O (g5702), .I (g56));
INVX1 gate2555(.O (g5703), .I (g109));
INVX1 gate2556(.O (g5704), .I (g219));
INVX1 gate2557(.O (g5705), .I (g225));
INVX1 gate2558(.O (g5706), .I (g231));
INVX1 gate2559(.O (g5707), .I (g109));
INVX1 gate2560(.O (g5708), .I (g303));
INVX1 gate2561(.O (g5712), .I (g305));
INVX1 gate2562(.O (I14163), .I (g113));
INVX1 gate2563(.O (g5713), .I (I14163));
INVX1 gate2564(.O (g5714), .I (g507));
INVX1 gate2565(.O (g5715), .I (g541));
INVX1 gate2566(.O (g5716), .I (g753));
INVX1 gate2567(.O (g5717), .I (g793));
INVX1 gate2568(.O (g5718), .I (g903));
INVX1 gate2569(.O (g5719), .I (g909));
INVX1 gate2570(.O (g5720), .I (g986));
INVX1 gate2571(.O (g5727), .I (g989));
INVX1 gate2572(.O (g5731), .I (g1192));
INVX1 gate2573(.O (g5732), .I (g1435));
INVX1 gate2574(.O (g5735), .I (g1476));
INVX1 gate2575(.O (g5736), .I (g1594));
INVX1 gate2576(.O (g5737), .I (g1682));
INVX1 gate2577(.O (I14182), .I (g1712));
INVX1 gate2578(.O (g5738), .I (I14182));
INVX1 gate2579(.O (g5741), .I (g2138));
INVX1 gate2580(.O (g5744), .I (g2195));
INVX1 gate2581(.O (g5745), .I (g2200));
INVX1 gate2582(.O (g5746), .I (g2375));
INVX1 gate2583(.O (I14191), .I (g2400));
INVX1 gate2584(.O (g5747), .I (I14191));
INVX1 gate2585(.O (I14195), .I (g3212));
INVX1 gate2586(.O (g5749), .I (I14195));
INVX1 gate2587(.O (g5750), .I (g92));
INVX1 gate2588(.O (g5751), .I (g52));
INVX1 gate2589(.O (g5752), .I (g113));
INVX1 gate2590(.O (g5753), .I (g228));
INVX1 gate2591(.O (g5754), .I (g234));
INVX1 gate2592(.O (g5755), .I (g240));
INVX1 gate2593(.O (g5756), .I (g304));
INVX1 gate2594(.O (g5759), .I (g508));
INVX1 gate2595(.O (g5760), .I (g744));
INVX1 gate2596(.O (g5761), .I (g797));
INVX1 gate2597(.O (g5762), .I (g906));
INVX1 gate2598(.O (g5763), .I (g912));
INVX1 gate2599(.O (g5764), .I (g918));
INVX1 gate2600(.O (g5765), .I (g797));
INVX1 gate2601(.O (g5766), .I (g990));
INVX1 gate2602(.O (g5770), .I (g992));
INVX1 gate2603(.O (I14219), .I (g801));
INVX1 gate2604(.O (g5771), .I (I14219));
INVX1 gate2605(.O (g5772), .I (g1193));
INVX1 gate2606(.O (g5773), .I (g1227));
INVX1 gate2607(.O (g5774), .I (g1439));
INVX1 gate2608(.O (g5775), .I (g1481));
INVX1 gate2609(.O (g5776), .I (g1597));
INVX1 gate2610(.O (g5777), .I (g1603));
INVX1 gate2611(.O (g5778), .I (g1680));
INVX1 gate2612(.O (g5785), .I (g1683));
INVX1 gate2613(.O (g5789), .I (g1886));
INVX1 gate2614(.O (g5790), .I (g2129));
INVX1 gate2615(.O (g5793), .I (g2170));
INVX1 gate2616(.O (g5794), .I (g2288));
INVX1 gate2617(.O (g5795), .I (g2376));
INVX1 gate2618(.O (I14238), .I (g2406));
INVX1 gate2619(.O (g5796), .I (I14238));
INVX1 gate2620(.O (I14243), .I (g3221));
INVX1 gate2621(.O (g5799), .I (I14243));
INVX1 gate2622(.O (I14246), .I (g3227));
INVX1 gate2623(.O (g5800), .I (I14246));
INVX1 gate2624(.O (I14249), .I (g3216));
INVX1 gate2625(.O (g5801), .I (I14249));
INVX1 gate2626(.O (g5802), .I (g83));
INVX1 gate2627(.O (g5803), .I (g117));
INVX1 gate2628(.O (g5804), .I (g237));
INVX1 gate2629(.O (g5805), .I (g243));
INVX1 gate2630(.O (g5806), .I (g249));
INVX1 gate2631(.O (g5808), .I (g509));
INVX1 gate2632(.O (g5809), .I (g780));
INVX1 gate2633(.O (g5810), .I (g740));
INVX1 gate2634(.O (g5811), .I (g801));
INVX1 gate2635(.O (g5812), .I (g915));
INVX1 gate2636(.O (g5813), .I (g921));
INVX1 gate2637(.O (g5814), .I (g927));
INVX1 gate2638(.O (g5815), .I (g991));
INVX1 gate2639(.O (g5818), .I (g1194));
INVX1 gate2640(.O (g5819), .I (g1430));
INVX1 gate2641(.O (g5820), .I (g1486));
INVX1 gate2642(.O (g5821), .I (g1600));
INVX1 gate2643(.O (g5822), .I (g1606));
INVX1 gate2644(.O (g5823), .I (g1612));
INVX1 gate2645(.O (g5824), .I (g1486));
INVX1 gate2646(.O (g5825), .I (g1684));
INVX1 gate2647(.O (g5829), .I (g1686));
INVX1 gate2648(.O (I14280), .I (g1491));
INVX1 gate2649(.O (g5830), .I (I14280));
INVX1 gate2650(.O (g5831), .I (g1887));
INVX1 gate2651(.O (g5832), .I (g1921));
INVX1 gate2652(.O (g5833), .I (g2133));
INVX1 gate2653(.O (g5834), .I (g2175));
INVX1 gate2654(.O (g5835), .I (g2291));
INVX1 gate2655(.O (g5836), .I (g2297));
INVX1 gate2656(.O (g5837), .I (g2374));
INVX1 gate2657(.O (g5844), .I (g2377));
INVX1 gate2658(.O (g5848), .I (g2580));
INVX1 gate2659(.O (I14295), .I (g3228));
INVX1 gate2660(.O (g5849), .I (I14295));
INVX1 gate2661(.O (I14298), .I (g3217));
INVX1 gate2662(.O (g5850), .I (I14298));
INVX1 gate2663(.O (g5851), .I (g74));
INVX1 gate2664(.O (g5852), .I (g121));
INVX1 gate2665(.O (g5853), .I (g246));
INVX1 gate2666(.O (g5854), .I (g252));
INVX1 gate2667(.O (g5855), .I (g258));
INVX1 gate2668(.O (I14306), .I (g97));
INVX1 gate2669(.O (g5856), .I (I14306));
INVX1 gate2670(.O (g5857), .I (g538));
INVX1 gate2671(.O (g5858), .I (g771));
INVX1 gate2672(.O (g5859), .I (g805));
INVX1 gate2673(.O (g5860), .I (g924));
INVX1 gate2674(.O (g5861), .I (g930));
INVX1 gate2675(.O (g5862), .I (g936));
INVX1 gate2676(.O (g5864), .I (g1195));
INVX1 gate2677(.O (g5865), .I (g1466));
INVX1 gate2678(.O (g5866), .I (g1426));
INVX1 gate2679(.O (g5867), .I (g1491));
INVX1 gate2680(.O (g5868), .I (g1609));
INVX1 gate2681(.O (g5869), .I (g1615));
INVX1 gate2682(.O (g5870), .I (g1621));
INVX1 gate2683(.O (g5871), .I (g1685));
INVX1 gate2684(.O (g5874), .I (g1888));
INVX1 gate2685(.O (g5875), .I (g2124));
INVX1 gate2686(.O (g5876), .I (g2180));
INVX1 gate2687(.O (g5877), .I (g2294));
INVX1 gate2688(.O (g5878), .I (g2300));
INVX1 gate2689(.O (g5879), .I (g2306));
INVX1 gate2690(.O (g5880), .I (g2180));
INVX1 gate2691(.O (g5881), .I (g2378));
INVX1 gate2692(.O (g5885), .I (g2380));
INVX1 gate2693(.O (I14338), .I (g2185));
INVX1 gate2694(.O (g5886), .I (I14338));
INVX1 gate2695(.O (g5887), .I (g2581));
INVX1 gate2696(.O (g5888), .I (g2615));
INVX1 gate2697(.O (I14343), .I (g3219));
INVX1 gate2698(.O (g5889), .I (I14343));
INVX1 gate2699(.O (g5890), .I (g88));
INVX1 gate2700(.O (g5893), .I (g125));
INVX1 gate2701(.O (g5894), .I (g186));
INVX1 gate2702(.O (g5895), .I (g255));
INVX1 gate2703(.O (g5896), .I (g261));
INVX1 gate2704(.O (g5897), .I (g267));
INVX1 gate2705(.O (g5898), .I (g762));
INVX1 gate2706(.O (g5899), .I (g809));
INVX1 gate2707(.O (g5900), .I (g933));
INVX1 gate2708(.O (g5901), .I (g939));
INVX1 gate2709(.O (g5902), .I (g945));
INVX1 gate2710(.O (I14357), .I (g785));
INVX1 gate2711(.O (g5903), .I (I14357));
INVX1 gate2712(.O (g5904), .I (g1224));
INVX1 gate2713(.O (g5905), .I (g1457));
INVX1 gate2714(.O (g5906), .I (g1496));
INVX1 gate2715(.O (g5907), .I (g1618));
INVX1 gate2716(.O (g5908), .I (g1624));
INVX1 gate2717(.O (g5909), .I (g1630));
INVX1 gate2718(.O (g5911), .I (g1889));
INVX1 gate2719(.O (g5912), .I (g2160));
INVX1 gate2720(.O (g5913), .I (g2120));
INVX1 gate2721(.O (g5914), .I (g2185));
INVX1 gate2722(.O (g5915), .I (g2303));
INVX1 gate2723(.O (g5916), .I (g2309));
INVX1 gate2724(.O (g5917), .I (g2315));
INVX1 gate2725(.O (g5918), .I (g2379));
INVX1 gate2726(.O (g5921), .I (g2582));
INVX1 gate2727(.O (I14378), .I (g3234));
INVX1 gate2728(.O (g5922), .I (I14378));
INVX1 gate2729(.O (I14381), .I (g3223));
INVX1 gate2730(.O (g5923), .I (I14381));
INVX1 gate2731(.O (I14384), .I (g3218));
INVX1 gate2732(.O (g5924), .I (I14384));
INVX1 gate2733(.O (g5925), .I (g189));
INVX1 gate2734(.O (g5926), .I (g195));
INVX1 gate2735(.O (g5927), .I (g264));
INVX1 gate2736(.O (g5928), .I (g270));
INVX1 gate2737(.O (g5929), .I (g776));
INVX1 gate2738(.O (g5932), .I (g813));
INVX1 gate2739(.O (g5933), .I (g873));
INVX1 gate2740(.O (g5934), .I (g942));
INVX1 gate2741(.O (g5935), .I (g948));
INVX1 gate2742(.O (g5936), .I (g954));
INVX1 gate2743(.O (g5937), .I (g1448));
INVX1 gate2744(.O (g5938), .I (g1501));
INVX1 gate2745(.O (g5939), .I (g1627));
INVX1 gate2746(.O (g5940), .I (g1633));
INVX1 gate2747(.O (g5941), .I (g1639));
INVX1 gate2748(.O (I14402), .I (g1471));
INVX1 gate2749(.O (g5942), .I (I14402));
INVX1 gate2750(.O (g5943), .I (g1918));
INVX1 gate2751(.O (g5944), .I (g2151));
INVX1 gate2752(.O (g5945), .I (g2190));
INVX1 gate2753(.O (g5946), .I (g2312));
INVX1 gate2754(.O (g5947), .I (g2318));
INVX1 gate2755(.O (g5948), .I (g2324));
INVX1 gate2756(.O (g5950), .I (g2583));
INVX1 gate2757(.O (I14413), .I (g3233));
INVX1 gate2758(.O (g5951), .I (I14413));
INVX1 gate2759(.O (I14416), .I (g3222));
INVX1 gate2760(.O (g5952), .I (I14416));
INVX1 gate2761(.O (g5953), .I (g97));
INVX1 gate2762(.O (g5954), .I (g192));
INVX1 gate2763(.O (g5955), .I (g198));
INVX1 gate2764(.O (g5956), .I (g204));
INVX1 gate2765(.O (g5957), .I (g273));
INVX1 gate2766(.O (I14424), .I (g117));
INVX1 gate2767(.O (g5958), .I (I14424));
INVX1 gate2768(.O (g5959), .I (g876));
INVX1 gate2769(.O (g5960), .I (g882));
INVX1 gate2770(.O (g5961), .I (g951));
INVX1 gate2771(.O (g5962), .I (g957));
INVX1 gate2772(.O (g5963), .I (g1462));
INVX1 gate2773(.O (g5966), .I (g1506));
INVX1 gate2774(.O (g5967), .I (g1567));
INVX1 gate2775(.O (g5968), .I (g1636));
INVX1 gate2776(.O (g5969), .I (g1642));
INVX1 gate2777(.O (g5970), .I (g1648));
INVX1 gate2778(.O (g5971), .I (g2142));
INVX1 gate2779(.O (g5972), .I (g2195));
INVX1 gate2780(.O (g5973), .I (g2321));
INVX1 gate2781(.O (g5974), .I (g2327));
INVX1 gate2782(.O (g5975), .I (g2333));
INVX1 gate2783(.O (I14442), .I (g2165));
INVX1 gate2784(.O (g5976), .I (I14442));
INVX1 gate2785(.O (g5977), .I (g2612));
INVX1 gate2786(.O (I14446), .I (g3230));
INVX1 gate2787(.O (g5978), .I (I14446));
INVX1 gate2788(.O (I14449), .I (g3224));
INVX1 gate2789(.O (g5979), .I (I14449));
INVX1 gate2790(.O (g5980), .I (g201));
INVX1 gate2791(.O (g5981), .I (g207));
INVX1 gate2792(.O (g5982), .I (g785));
INVX1 gate2793(.O (g5983), .I (g879));
INVX1 gate2794(.O (g5984), .I (g885));
INVX1 gate2795(.O (g5985), .I (g891));
INVX1 gate2796(.O (g5986), .I (g960));
INVX1 gate2797(.O (I14459), .I (g805));
INVX1 gate2798(.O (g5987), .I (I14459));
INVX1 gate2799(.O (g5988), .I (g1570));
INVX1 gate2800(.O (g5989), .I (g1576));
INVX1 gate2801(.O (g5990), .I (g1645));
INVX1 gate2802(.O (g5991), .I (g1651));
INVX1 gate2803(.O (g5992), .I (g2156));
INVX1 gate2804(.O (g5995), .I (g2200));
INVX1 gate2805(.O (g5996), .I (g2261));
INVX1 gate2806(.O (g5997), .I (g2330));
INVX1 gate2807(.O (g5998), .I (g2336));
INVX1 gate2808(.O (g5999), .I (g2342));
INVX1 gate2809(.O (I14472), .I (g3080));
INVX1 gate2810(.O (g6000), .I (I14472));
INVX1 gate2811(.O (I14475), .I (g3225));
INVX1 gate2812(.O (g6014), .I (I14475));
INVX1 gate2813(.O (I14478), .I (g3213));
INVX1 gate2814(.O (g6015), .I (I14478));
INVX1 gate2815(.O (g6016), .I (g210));
INVX1 gate2816(.O (g6017), .I (g888));
INVX1 gate2817(.O (g6018), .I (g894));
INVX1 gate2818(.O (g6019), .I (g1471));
INVX1 gate2819(.O (g6020), .I (g1573));
INVX1 gate2820(.O (g6021), .I (g1579));
INVX1 gate2821(.O (g6022), .I (g1585));
INVX1 gate2822(.O (g6023), .I (g1654));
INVX1 gate2823(.O (I14489), .I (g1496));
INVX1 gate2824(.O (g6024), .I (I14489));
INVX1 gate2825(.O (g6025), .I (g2264));
INVX1 gate2826(.O (g6026), .I (g2270));
INVX1 gate2827(.O (g6027), .I (g2339));
INVX1 gate2828(.O (g6028), .I (g2345));
INVX1 gate2829(.O (I14496), .I (g3226));
INVX1 gate2830(.O (g6029), .I (I14496));
INVX1 gate2831(.O (I14499), .I (g3214));
INVX1 gate2832(.O (g6030), .I (I14499));
INVX1 gate2833(.O (I14502), .I (g471));
INVX1 gate2834(.O (g6031), .I (I14502));
INVX1 gate2835(.O (g6032), .I (g897));
INVX1 gate2836(.O (g6033), .I (g1582));
INVX1 gate2837(.O (g6034), .I (g1588));
INVX1 gate2838(.O (g6035), .I (g2165));
INVX1 gate2839(.O (g6036), .I (g2267));
INVX1 gate2840(.O (g6037), .I (g2273));
INVX1 gate2841(.O (g6038), .I (g2279));
INVX1 gate2842(.O (g6039), .I (g2348));
INVX1 gate2843(.O (I14513), .I (g2190));
INVX1 gate2844(.O (g6040), .I (I14513));
INVX1 gate2845(.O (I14516), .I (g3215));
INVX1 gate2846(.O (g6041), .I (I14516));
INVX1 gate2847(.O (I14519), .I (g1158));
INVX1 gate2848(.O (g6042), .I (I14519));
INVX1 gate2849(.O (g6043), .I (g1591));
INVX1 gate2850(.O (g6044), .I (g2276));
INVX1 gate2851(.O (g6045), .I (g2282));
INVX1 gate2852(.O (I14525), .I (g1852));
INVX1 gate2853(.O (g6046), .I (I14525));
INVX1 gate2854(.O (g6047), .I (g2285));
INVX1 gate2855(.O (I14529), .I (g3142));
INVX1 gate2856(.O (g6048), .I (I14529));
INVX1 gate2857(.O (I14532), .I (g354));
INVX1 gate2858(.O (g6051), .I (I14532));
INVX1 gate2859(.O (I14535), .I (g2546));
INVX1 gate2860(.O (g6052), .I (I14535));
INVX1 gate2861(.O (I14538), .I (g369));
INVX1 gate2862(.O (g6053), .I (I14538));
INVX1 gate2863(.O (I14541), .I (g455));
INVX1 gate2864(.O (g6054), .I (I14541));
INVX1 gate2865(.O (I14544), .I (g1041));
INVX1 gate2866(.O (g6055), .I (I14544));
INVX1 gate2867(.O (I14547), .I (g384));
INVX1 gate2868(.O (g6056), .I (I14547));
INVX1 gate2869(.O (I14550), .I (g458));
INVX1 gate2870(.O (g6057), .I (I14550));
INVX1 gate2871(.O (I14553), .I (g1056));
INVX1 gate2872(.O (g6058), .I (I14553));
INVX1 gate2873(.O (I14556), .I (g1142));
INVX1 gate2874(.O (g6059), .I (I14556));
INVX1 gate2875(.O (I14559), .I (g1735));
INVX1 gate2876(.O (g6060), .I (I14559));
INVX1 gate2877(.O (I14562), .I (g398));
INVX1 gate2878(.O (g6061), .I (I14562));
INVX1 gate2879(.O (I14565), .I (g461));
INVX1 gate2880(.O (g6062), .I (I14565));
INVX1 gate2881(.O (I14568), .I (g1071));
INVX1 gate2882(.O (g6063), .I (I14568));
INVX1 gate2883(.O (I14571), .I (g1145));
INVX1 gate2884(.O (g6064), .I (I14571));
INVX1 gate2885(.O (I14574), .I (g1750));
INVX1 gate2886(.O (g6065), .I (I14574));
INVX1 gate2887(.O (I14577), .I (g1836));
INVX1 gate2888(.O (g6066), .I (I14577));
INVX1 gate2889(.O (I14580), .I (g2429));
INVX1 gate2890(.O (g6067), .I (I14580));
INVX1 gate2891(.O (g6068), .I (g499));
INVX1 gate2892(.O (I14584), .I (g465));
INVX1 gate2893(.O (g6079), .I (I14584));
INVX1 gate2894(.O (I14587), .I (g1085));
INVX1 gate2895(.O (g6080), .I (I14587));
INVX1 gate2896(.O (I14590), .I (g1148));
INVX1 gate2897(.O (g6081), .I (I14590));
INVX1 gate2898(.O (I14593), .I (g1765));
INVX1 gate2899(.O (g6082), .I (I14593));
INVX1 gate2900(.O (I14596), .I (g1839));
INVX1 gate2901(.O (g6083), .I (I14596));
INVX1 gate2902(.O (I14599), .I (g2444));
INVX1 gate2903(.O (g6084), .I (I14599));
INVX1 gate2904(.O (I14602), .I (g2530));
INVX1 gate2905(.O (g6085), .I (I14602));
INVX1 gate2906(.O (I14605), .I (g468));
INVX1 gate2907(.O (g6086), .I (I14605));
INVX1 gate2908(.O (g6087), .I (g1186));
INVX1 gate2909(.O (I14609), .I (g1152));
INVX1 gate2910(.O (g6098), .I (I14609));
INVX1 gate2911(.O (I14612), .I (g1779));
INVX1 gate2912(.O (g6099), .I (I14612));
INVX1 gate2913(.O (I14615), .I (g1842));
INVX1 gate2914(.O (g6100), .I (I14615));
INVX1 gate2915(.O (I14618), .I (g2459));
INVX1 gate2916(.O (g6101), .I (I14618));
INVX1 gate2917(.O (I14621), .I (g2533));
INVX1 gate2918(.O (g6102), .I (I14621));
INVX1 gate2919(.O (I14624), .I (g1155));
INVX1 gate2920(.O (g6103), .I (I14624));
INVX1 gate2921(.O (g6104), .I (g1880));
INVX1 gate2922(.O (I14628), .I (g1846));
INVX1 gate2923(.O (g6115), .I (I14628));
INVX1 gate2924(.O (I14631), .I (g2473));
INVX1 gate2925(.O (g6116), .I (I14631));
INVX1 gate2926(.O (I14634), .I (g2536));
INVX1 gate2927(.O (g6117), .I (I14634));
INVX1 gate2928(.O (I14637), .I (g1849));
INVX1 gate2929(.O (g6118), .I (I14637));
INVX1 gate2930(.O (g6119), .I (g2574));
INVX1 gate2931(.O (I14641), .I (g2540));
INVX1 gate2932(.O (g6130), .I (I14641));
INVX1 gate2933(.O (I14644), .I (g3142));
INVX1 gate2934(.O (g6131), .I (I14644));
INVX1 gate2935(.O (I14647), .I (g2543));
INVX1 gate2936(.O (g6134), .I (I14647));
INVX1 gate2937(.O (I14650), .I (g525));
INVX1 gate2938(.O (g6135), .I (I14650));
INVX1 gate2939(.O (g6136), .I (g672));
INVX1 gate2940(.O (I14654), .I (g3220));
INVX1 gate2941(.O (g6139), .I (I14654));
INVX1 gate2942(.O (g6140), .I (g524));
INVX1 gate2943(.O (g6141), .I (g554));
INVX1 gate2944(.O (g6142), .I (g679));
INVX1 gate2945(.O (I14660), .I (g1211));
INVX1 gate2946(.O (g6145), .I (I14660));
INVX1 gate2947(.O (g6146), .I (g1358));
INVX1 gate2948(.O (g6149), .I (g3097));
INVX1 gate2949(.O (I14665), .I (g3147));
INVX1 gate2950(.O (g6153), .I (I14665));
INVX1 gate2951(.O (I14668), .I (g3232));
INVX1 gate2952(.O (g6156), .I (I14668));
INVX1 gate2953(.O (g6157), .I (g686));
INVX1 gate2954(.O (g6161), .I (g1210));
INVX1 gate2955(.O (g6162), .I (g1240));
INVX1 gate2956(.O (g6163), .I (g1365));
INVX1 gate2957(.O (I14675), .I (g1905));
INVX1 gate2958(.O (g6166), .I (I14675));
INVX1 gate2959(.O (g6167), .I (g2052));
INVX1 gate2960(.O (g6170), .I (g3098));
INVX1 gate2961(.O (g6173), .I (g557));
INVX1 gate2962(.O (g6177), .I (g633));
INVX1 gate2963(.O (g6180), .I (g692));
INVX1 gate2964(.O (g6183), .I (g291));
INVX1 gate2965(.O (g6184), .I (g1372));
INVX1 gate2966(.O (g6188), .I (g1904));
INVX1 gate2967(.O (g6189), .I (g1934));
INVX1 gate2968(.O (g6190), .I (g2059));
INVX1 gate2969(.O (I14688), .I (g2599));
INVX1 gate2970(.O (g6193), .I (I14688));
INVX1 gate2971(.O (g6194), .I (g2746));
INVX1 gate2972(.O (g6197), .I (g3099));
INVX1 gate2973(.O (g6200), .I (g542));
INVX1 gate2974(.O (g6201), .I (g646));
INVX1 gate2975(.O (g6204), .I (g289));
INVX1 gate2976(.O (g6205), .I (g1243));
INVX1 gate2977(.O (g6209), .I (g1319));
INVX1 gate2978(.O (g6212), .I (g1378));
INVX1 gate2979(.O (g6215), .I (g978));
INVX1 gate2980(.O (g6216), .I (g2066));
INVX1 gate2981(.O (g6220), .I (g2598));
INVX1 gate2982(.O (g6221), .I (g2628));
INVX1 gate2983(.O (g6222), .I (g2753));
INVX1 gate2984(.O (I14704), .I (g2818));
INVX1 gate2985(.O (g6225), .I (I14704));
INVX1 gate2986(.O (g6226), .I (g2818));
INVX1 gate2987(.O (g6227), .I (g3100));
INVX1 gate2988(.O (I14709), .I (g3229));
INVX1 gate2989(.O (g6230), .I (I14709));
INVX1 gate2990(.O (I14712), .I (g138));
INVX1 gate2991(.O (g6231), .I (I14712));
INVX1 gate2992(.O (I14715), .I (g138));
INVX1 gate2993(.O (g6232), .I (I14715));
INVX1 gate2994(.O (g6281), .I (g510));
INVX1 gate2995(.O (g6284), .I (g640));
INVX1 gate2996(.O (g6288), .I (g287));
INVX1 gate2997(.O (g6289), .I (g1228));
INVX1 gate2998(.O (g6290), .I (g1332));
INVX1 gate2999(.O (g6293), .I (g976));
INVX1 gate3000(.O (g6294), .I (g1937));
INVX1 gate3001(.O (g6298), .I (g2013));
INVX1 gate3002(.O (g6301), .I (g2072));
INVX1 gate3003(.O (g6304), .I (g1672));
INVX1 gate3004(.O (g6305), .I (g2760));
INVX1 gate3005(.O (g6309), .I (g14));
INVX1 gate3006(.O (g6310), .I (g3101));
INVX1 gate3007(.O (I14731), .I (g135));
INVX1 gate3008(.O (g6313), .I (I14731));
INVX1 gate3009(.O (I14734), .I (g135));
INVX1 gate3010(.O (g6314), .I (I14734));
INVX1 gate3011(.O (g6363), .I (g653));
INVX1 gate3012(.O (g6367), .I (g285));
INVX1 gate3013(.O (I14739), .I (g826));
INVX1 gate3014(.O (g6368), .I (I14739));
INVX1 gate3015(.O (I14742), .I (g826));
INVX1 gate3016(.O (g6369), .I (I14742));
INVX1 gate3017(.O (g6418), .I (g1196));
INVX1 gate3018(.O (g6421), .I (g1326));
INVX1 gate3019(.O (g6425), .I (g974));
INVX1 gate3020(.O (g6426), .I (g1922));
INVX1 gate3021(.O (g6427), .I (g2026));
INVX1 gate3022(.O (g6430), .I (g1670));
INVX1 gate3023(.O (g6431), .I (g2631));
INVX1 gate3024(.O (g6435), .I (g2707));
INVX1 gate3025(.O (g6438), .I (g2766));
INVX1 gate3026(.O (g6441), .I (g2366));
INVX1 gate3027(.O (I14755), .I (g2821));
INVX1 gate3028(.O (g6442), .I (I14755));
INVX1 gate3029(.O (g6443), .I (g2821));
INVX1 gate3030(.O (g6444), .I (g3102));
INVX1 gate3031(.O (I14760), .I (g405));
INVX1 gate3032(.O (g6447), .I (I14760));
INVX1 gate3033(.O (I14763), .I (g405));
INVX1 gate3034(.O (g6448), .I (I14763));
INVX1 gate3035(.O (I14766), .I (g545));
INVX1 gate3036(.O (g6485), .I (I14766));
INVX1 gate3037(.O (I14769), .I (g545));
INVX1 gate3038(.O (g6486), .I (I14769));
INVX1 gate3039(.O (g6512), .I (g544));
INVX1 gate3040(.O (g6513), .I (g660));
INVX1 gate3041(.O (g6517), .I (g283));
INVX1 gate3042(.O (I14775), .I (g823));
INVX1 gate3043(.O (g6518), .I (I14775));
INVX1 gate3044(.O (I14778), .I (g823));
INVX1 gate3045(.O (g6519), .I (I14778));
INVX1 gate3046(.O (g6568), .I (g1339));
INVX1 gate3047(.O (g6572), .I (g972));
INVX1 gate3048(.O (I14783), .I (g1520));
INVX1 gate3049(.O (g6573), .I (I14783));
INVX1 gate3050(.O (I14786), .I (g1520));
INVX1 gate3051(.O (g6574), .I (I14786));
INVX1 gate3052(.O (g6623), .I (g1890));
INVX1 gate3053(.O (g6626), .I (g2020));
INVX1 gate3054(.O (g6630), .I (g1668));
INVX1 gate3055(.O (g6631), .I (g2616));
INVX1 gate3056(.O (g6632), .I (g2720));
INVX1 gate3057(.O (g6635), .I (g2364));
INVX1 gate3058(.O (g6636), .I (g1491));
INVX1 gate3059(.O (g6637), .I (g5));
INVX1 gate3060(.O (g6638), .I (g3103));
INVX1 gate3061(.O (g6641), .I (g113));
INVX1 gate3062(.O (I14799), .I (g551));
INVX1 gate3063(.O (g6642), .I (I14799));
INVX1 gate3064(.O (I14802), .I (g551));
INVX1 gate3065(.O (g6643), .I (I14802));
INVX1 gate3066(.O (g6672), .I (g464));
INVX1 gate3067(.O (g6675), .I (g458));
INVX1 gate3068(.O (g6676), .I (g559));
INVX1 gate3069(.O (I14808), .I (g623));
INVX1 gate3070(.O (g6677), .I (I14808));
INVX1 gate3071(.O (I14811), .I (g623));
INVX1 gate3072(.O (g6678), .I (I14811));
INVX1 gate3073(.O (g6707), .I (g666));
INVX1 gate3074(.O (g6711), .I (g281));
INVX1 gate3075(.O (I14816), .I (g1092));
INVX1 gate3076(.O (g6712), .I (I14816));
INVX1 gate3077(.O (I14819), .I (g1092));
INVX1 gate3078(.O (g6713), .I (I14819));
INVX1 gate3079(.O (I14822), .I (g1231));
INVX1 gate3080(.O (g6750), .I (I14822));
INVX1 gate3081(.O (I14825), .I (g1231));
INVX1 gate3082(.O (g6751), .I (I14825));
INVX1 gate3083(.O (g6776), .I (g1230));
INVX1 gate3084(.O (g6777), .I (g1346));
INVX1 gate3085(.O (g6781), .I (g970));
INVX1 gate3086(.O (I14831), .I (g1517));
INVX1 gate3087(.O (g6782), .I (I14831));
INVX1 gate3088(.O (I14834), .I (g1517));
INVX1 gate3089(.O (g6783), .I (I14834));
INVX1 gate3090(.O (g6832), .I (g2033));
INVX1 gate3091(.O (g6836), .I (g1666));
INVX1 gate3092(.O (I14839), .I (g2214));
INVX1 gate3093(.O (g6837), .I (I14839));
INVX1 gate3094(.O (I14842), .I (g2214));
INVX1 gate3095(.O (g6838), .I (I14842));
INVX1 gate3096(.O (g6887), .I (g2584));
INVX1 gate3097(.O (g6890), .I (g2714));
INVX1 gate3098(.O (g6894), .I (g2362));
INVX1 gate3099(.O (I14848), .I (g2824));
INVX1 gate3100(.O (g6895), .I (I14848));
INVX1 gate3101(.O (g6896), .I (g2824));
INVX1 gate3102(.O (g6897), .I (g1486));
INVX1 gate3103(.O (g6898), .I (g2993));
INVX1 gate3104(.O (g6901), .I (g3006));
INVX1 gate3105(.O (g6905), .I (g3104));
INVX1 gate3106(.O (g6908), .I (g484));
INVX1 gate3107(.O (I14857), .I (g626));
INVX1 gate3108(.O (g6911), .I (I14857));
INVX1 gate3109(.O (I14860), .I (g626));
INVX1 gate3110(.O (g6912), .I (I14860));
INVX1 gate3111(.O (g6942), .I (g279));
INVX1 gate3112(.O (g6943), .I (g801));
INVX1 gate3113(.O (I14865), .I (g1237));
INVX1 gate3114(.O (g6944), .I (I14865));
INVX1 gate3115(.O (I14868), .I (g1237));
INVX1 gate3116(.O (g6945), .I (I14868));
INVX1 gate3117(.O (g6974), .I (g1151));
INVX1 gate3118(.O (g6977), .I (g1145));
INVX1 gate3119(.O (g6978), .I (g1245));
INVX1 gate3120(.O (I14874), .I (g1309));
INVX1 gate3121(.O (g6979), .I (I14874));
INVX1 gate3122(.O (I14877), .I (g1309));
INVX1 gate3123(.O (g6980), .I (I14877));
INVX1 gate3124(.O (g7009), .I (g1352));
INVX1 gate3125(.O (g7013), .I (g968));
INVX1 gate3126(.O (I14882), .I (g1786));
INVX1 gate3127(.O (g7014), .I (I14882));
INVX1 gate3128(.O (I14885), .I (g1786));
INVX1 gate3129(.O (g7015), .I (I14885));
INVX1 gate3130(.O (I14888), .I (g1925));
INVX1 gate3131(.O (g7052), .I (I14888));
INVX1 gate3132(.O (I14891), .I (g1925));
INVX1 gate3133(.O (g7053), .I (I14891));
INVX1 gate3134(.O (g7078), .I (g1924));
INVX1 gate3135(.O (g7079), .I (g2040));
INVX1 gate3136(.O (g7083), .I (g1664));
INVX1 gate3137(.O (I14897), .I (g2211));
INVX1 gate3138(.O (g7084), .I (I14897));
INVX1 gate3139(.O (I14900), .I (g2211));
INVX1 gate3140(.O (g7085), .I (I14900));
INVX1 gate3141(.O (g7134), .I (g2727));
INVX1 gate3142(.O (g7138), .I (g2360));
INVX1 gate3143(.O (g7139), .I (g1481));
INVX1 gate3144(.O (g7140), .I (g2170));
INVX1 gate3145(.O (g7141), .I (g2195));
INVX1 gate3146(.O (g7142), .I (g8));
INVX1 gate3147(.O (g7143), .I (g2998));
INVX1 gate3148(.O (g7146), .I (g3013));
INVX1 gate3149(.O (g7149), .I (g3105));
INVX1 gate3150(.O (g7152), .I (g3136));
INVX1 gate3151(.O (g7153), .I (g480));
INVX1 gate3152(.O (g7156), .I (g461));
INVX1 gate3153(.O (g7157), .I (g453));
INVX1 gate3154(.O (g7158), .I (g1171));
INVX1 gate3155(.O (I14917), .I (g1312));
INVX1 gate3156(.O (g7161), .I (I14917));
INVX1 gate3157(.O (I14920), .I (g1312));
INVX1 gate3158(.O (g7162), .I (I14920));
INVX1 gate3159(.O (g7192), .I (g966));
INVX1 gate3160(.O (g7193), .I (g1491));
INVX1 gate3161(.O (I14925), .I (g1931));
INVX1 gate3162(.O (g7194), .I (I14925));
INVX1 gate3163(.O (I14928), .I (g1931));
INVX1 gate3164(.O (g7195), .I (I14928));
INVX1 gate3165(.O (g7224), .I (g1845));
INVX1 gate3166(.O (g7227), .I (g1839));
INVX1 gate3167(.O (g7228), .I (g1939));
INVX1 gate3168(.O (I14934), .I (g2003));
INVX1 gate3169(.O (g7229), .I (I14934));
INVX1 gate3170(.O (I14937), .I (g2003));
INVX1 gate3171(.O (g7230), .I (I14937));
INVX1 gate3172(.O (g7259), .I (g2046));
INVX1 gate3173(.O (g7263), .I (g1662));
INVX1 gate3174(.O (I14942), .I (g2480));
INVX1 gate3175(.O (g7264), .I (I14942));
INVX1 gate3176(.O (I14945), .I (g2480));
INVX1 gate3177(.O (g7265), .I (I14945));
INVX1 gate3178(.O (I14948), .I (g2619));
INVX1 gate3179(.O (g7302), .I (I14948));
INVX1 gate3180(.O (I14951), .I (g2619));
INVX1 gate3181(.O (g7303), .I (I14951));
INVX1 gate3182(.O (g7328), .I (g2618));
INVX1 gate3183(.O (g7329), .I (g2734));
INVX1 gate3184(.O (g7333), .I (g2358));
INVX1 gate3185(.O (I14957), .I (g2827));
INVX1 gate3186(.O (g7334), .I (I14957));
INVX1 gate3187(.O (g7335), .I (g2827));
INVX1 gate3188(.O (g7336), .I (g1476));
INVX1 gate3189(.O (g7337), .I (g2190));
INVX1 gate3190(.O (g7338), .I (g3002));
INVX1 gate3191(.O (g7342), .I (g3024));
INVX1 gate3192(.O (g7345), .I (g3139));
INVX1 gate3193(.O (g7346), .I (g97));
INVX1 gate3194(.O (g7347), .I (g490));
INVX1 gate3195(.O (g7348), .I (g451));
INVX1 gate3196(.O (g7349), .I (g1167));
INVX1 gate3197(.O (g7352), .I (g1148));
INVX1 gate3198(.O (g7353), .I (g1140));
INVX1 gate3199(.O (g7354), .I (g1865));
INVX1 gate3200(.O (I14973), .I (g2006));
INVX1 gate3201(.O (g7357), .I (I14973));
INVX1 gate3202(.O (I14976), .I (g2006));
INVX1 gate3203(.O (g7358), .I (I14976));
INVX1 gate3204(.O (g7388), .I (g1660));
INVX1 gate3205(.O (g7389), .I (g2185));
INVX1 gate3206(.O (I14981), .I (g2625));
INVX1 gate3207(.O (g7390), .I (I14981));
INVX1 gate3208(.O (I14984), .I (g2625));
INVX1 gate3209(.O (g7391), .I (I14984));
INVX1 gate3210(.O (g7420), .I (g2539));
INVX1 gate3211(.O (g7423), .I (g2533));
INVX1 gate3212(.O (g7424), .I (g2633));
INVX1 gate3213(.O (I14990), .I (g2697));
INVX1 gate3214(.O (g7425), .I (I14990));
INVX1 gate3215(.O (I14993), .I (g2697));
INVX1 gate3216(.O (g7426), .I (I14993));
INVX1 gate3217(.O (g7455), .I (g2740));
INVX1 gate3218(.O (g7459), .I (g2356));
INVX1 gate3219(.O (g7460), .I (g1471));
INVX1 gate3220(.O (g7461), .I (g2175));
INVX1 gate3221(.O (g7462), .I (g2912));
INVX1 gate3222(.O (g7465), .I (g2));
INVX1 gate3223(.O (g7466), .I (g3010));
INVX1 gate3224(.O (g7471), .I (g3036));
INVX1 gate3225(.O (g7475), .I (g493));
INVX1 gate3226(.O (g7476), .I (g785));
INVX1 gate3227(.O (g7477), .I (g1177));
INVX1 gate3228(.O (g7478), .I (g1138));
INVX1 gate3229(.O (g7479), .I (g1861));
INVX1 gate3230(.O (g7482), .I (g1842));
INVX1 gate3231(.O (g7483), .I (g1834));
INVX1 gate3232(.O (g7484), .I (g2559));
INVX1 gate3233(.O (I15012), .I (g2700));
INVX1 gate3234(.O (g7487), .I (I15012));
INVX1 gate3235(.O (I15015), .I (g2700));
INVX1 gate3236(.O (g7488), .I (I15015));
INVX1 gate3237(.O (g7518), .I (g2354));
INVX1 gate3238(.O (I15019), .I (g2830));
INVX1 gate3239(.O (g7519), .I (I15019));
INVX1 gate3240(.O (g7520), .I (g2830));
INVX1 gate3241(.O (g7521), .I (g2200));
INVX1 gate3242(.O (g7522), .I (g2917));
INVX1 gate3243(.O (g7527), .I (g3018));
INVX1 gate3244(.O (g7529), .I (g465));
INVX1 gate3245(.O (g7530), .I (g496));
INVX1 gate3246(.O (g7531), .I (g1180));
INVX1 gate3247(.O (g7532), .I (g1471));
INVX1 gate3248(.O (g7533), .I (g1871));
INVX1 gate3249(.O (g7534), .I (g1832));
INVX1 gate3250(.O (g7535), .I (g2555));
INVX1 gate3251(.O (g7538), .I (g2536));
INVX1 gate3252(.O (g7539), .I (g2528));
INVX1 gate3253(.O (g7540), .I (g1506));
INVX1 gate3254(.O (g7541), .I (g2180));
INVX1 gate3255(.O (g7542), .I (g2883));
INVX1 gate3256(.O (g7545), .I (g2920));
INVX1 gate3257(.O (g7548), .I (g2990));
INVX1 gate3258(.O (g7549), .I (g3028));
INVX1 gate3259(.O (g7553), .I (g3114));
INVX1 gate3260(.O (g7554), .I (g117));
INVX1 gate3261(.O (g7555), .I (g1152));
INVX1 gate3262(.O (g7556), .I (g1183));
INVX1 gate3263(.O (g7557), .I (g1874));
INVX1 gate3264(.O (g7558), .I (g2165));
INVX1 gate3265(.O (g7559), .I (g2565));
INVX1 gate3266(.O (g7560), .I (g2526));
INVX1 gate3267(.O (g7561), .I (g1501));
INVX1 gate3268(.O (g7562), .I (g2888));
INVX1 gate3269(.O (g7566), .I (g2896));
INVX1 gate3270(.O (g7570), .I (g3032));
INVX1 gate3271(.O (g7573), .I (g3120));
INVX1 gate3272(.O (g7574), .I (g3128));
INVX1 gate3273(.O (g7576), .I (g468));
INVX1 gate3274(.O (g7577), .I (g805));
INVX1 gate3275(.O (g7578), .I (g1846));
INVX1 gate3276(.O (g7579), .I (g1877));
INVX1 gate3277(.O (g7580), .I (g2568));
INVX1 gate3278(.O (g7581), .I (g1496));
INVX1 gate3279(.O (g7582), .I (g2185));
INVX1 gate3280(.O (g7583), .I (g2892));
INVX1 gate3281(.O (g7587), .I (g2903));
INVX1 gate3282(.O (g7590), .I (g1155));
INVX1 gate3283(.O (g7591), .I (g1496));
INVX1 gate3284(.O (g7592), .I (g2540));
INVX1 gate3285(.O (g7593), .I (g2571));
INVX1 gate3286(.O (g7594), .I (g2165));
INVX1 gate3287(.O (g7595), .I (g2900));
INVX1 gate3288(.O (g7600), .I (g2908));
INVX1 gate3289(.O (g7603), .I (g3133));
INVX1 gate3290(.O (g7604), .I (g471));
INVX1 gate3291(.O (g7605), .I (g1849));
INVX1 gate3292(.O (g7606), .I (g2190));
INVX1 gate3293(.O (g7607), .I (g2924));
INVX1 gate3294(.O (g7610), .I (g312));
INVX1 gate3295(.O (g7613), .I (g1158));
INVX1 gate3296(.O (g7614), .I (g2543));
INVX1 gate3297(.O (g7615), .I (g3123));
INVX1 gate3298(.O (g7616), .I (g313));
INVX1 gate3299(.O (g7619), .I (g999));
INVX1 gate3300(.O (g7622), .I (g1852));
INVX1 gate3301(.O (g7623), .I (g314));
INVX1 gate3302(.O (g7626), .I (g315));
INVX1 gate3303(.O (g7629), .I (g403));
INVX1 gate3304(.O (g7632), .I (g1000));
INVX1 gate3305(.O (g7635), .I (g1693));
INVX1 gate3306(.O (g7638), .I (g2546));
INVX1 gate3307(.O (g7639), .I (g3094));
INVX1 gate3308(.O (g7642), .I (g3125));
INVX1 gate3309(.O (g7643), .I (g316));
INVX1 gate3310(.O (g7646), .I (g318));
INVX1 gate3311(.O (g7649), .I (g404));
INVX1 gate3312(.O (g7652), .I (g1001));
INVX1 gate3313(.O (g7655), .I (g1002));
INVX1 gate3314(.O (g7658), .I (g1090));
INVX1 gate3315(.O (g7661), .I (g1694));
INVX1 gate3316(.O (g7664), .I (g2387));
INVX1 gate3317(.O (g7667), .I (g3095));
INVX1 gate3318(.O (g7670), .I (g317));
INVX1 gate3319(.O (g7673), .I (g319));
INVX1 gate3320(.O (g7676), .I (g402));
INVX1 gate3321(.O (g7679), .I (g1003));
INVX1 gate3322(.O (g7682), .I (g1005));
INVX1 gate3323(.O (g7685), .I (g1091));
INVX1 gate3324(.O (g7688), .I (g1695));
INVX1 gate3325(.O (g7691), .I (g1696));
INVX1 gate3326(.O (g7694), .I (g1784));
INVX1 gate3327(.O (g7697), .I (g2388));
INVX1 gate3328(.O (g7700), .I (g3096));
INVX1 gate3329(.O (g7703), .I (g320));
INVX1 gate3330(.O (g7706), .I (g1004));
INVX1 gate3331(.O (g7709), .I (g1006));
INVX1 gate3332(.O (g7712), .I (g1089));
INVX1 gate3333(.O (g7715), .I (g1697));
INVX1 gate3334(.O (g7718), .I (g1699));
INVX1 gate3335(.O (g7721), .I (g1785));
INVX1 gate3336(.O (g7724), .I (g2389));
INVX1 gate3337(.O (g7727), .I (g2390));
INVX1 gate3338(.O (g7730), .I (g2478));
INVX1 gate3339(.O (g7733), .I (g1007));
INVX1 gate3340(.O (g7736), .I (g1698));
INVX1 gate3341(.O (g7739), .I (g1700));
INVX1 gate3342(.O (g7742), .I (g1783));
INVX1 gate3343(.O (g7745), .I (g2391));
INVX1 gate3344(.O (g7748), .I (g2393));
INVX1 gate3345(.O (g7751), .I (g2479));
INVX1 gate3346(.O (g7754), .I (g322));
INVX1 gate3347(.O (g7757), .I (g1701));
INVX1 gate3348(.O (g7760), .I (g2392));
INVX1 gate3349(.O (g7763), .I (g2394));
INVX1 gate3350(.O (g7766), .I (g2477));
INVX1 gate3351(.O (g7769), .I (g323));
INVX1 gate3352(.O (g7772), .I (g659));
INVX1 gate3353(.O (g7776), .I (g1009));
INVX1 gate3354(.O (g7779), .I (g2395));
INVX1 gate3355(.O (g7782), .I (g321));
INVX1 gate3356(.O (g7785), .I (g1010));
INVX1 gate3357(.O (g7788), .I (g1345));
INVX1 gate3358(.O (g7792), .I (g1703));
INVX1 gate3359(.O (g7796), .I (g1008));
INVX1 gate3360(.O (g7799), .I (g1704));
INVX1 gate3361(.O (g7802), .I (g2039));
INVX1 gate3362(.O (g7806), .I (g2397));
INVX1 gate3363(.O (g7809), .I (g1702));
INVX1 gate3364(.O (g7812), .I (g2398));
INVX1 gate3365(.O (g7815), .I (g2733));
INVX1 gate3366(.O (g7819), .I (g479));
INVX1 gate3367(.O (g7822), .I (g510));
INVX1 gate3368(.O (g7823), .I (g2396));
INVX1 gate3369(.O (g7826), .I (g2987));
INVX1 gate3370(.O (g7827), .I (g478));
INVX1 gate3371(.O (g7830), .I (g1166));
INVX1 gate3372(.O (g7833), .I (g1196));
INVX1 gate3373(.O (g7834), .I (g2953));
INVX1 gate3374(.O (g7837), .I (g3044));
INVX1 gate3375(.O (g7838), .I (g477));
INVX1 gate3376(.O (g7841), .I (g630));
INVX1 gate3377(.O (g7842), .I (g1165));
INVX1 gate3378(.O (g7845), .I (g1860));
INVX1 gate3379(.O (g7848), .I (g1890));
INVX1 gate3380(.O (g7849), .I (g2956));
INVX1 gate3381(.O (g7852), .I (g2981));
INVX1 gate3382(.O (g7856), .I (g3045));
INVX1 gate3383(.O (g7857), .I (g3055));
INVX1 gate3384(.O (g7858), .I (g1164));
INVX1 gate3385(.O (g7861), .I (g1316));
INVX1 gate3386(.O (g7862), .I (g1859));
INVX1 gate3387(.O (g7865), .I (g2554));
INVX1 gate3388(.O (g7868), .I (g2584));
INVX1 gate3389(.O (g7869), .I (g2959));
INVX1 gate3390(.O (g7872), .I (g2874));
INVX1 gate3391(.O (g7877), .I (g3046));
INVX1 gate3392(.O (g7878), .I (g3056));
INVX1 gate3393(.O (g7879), .I (g3065));
INVX1 gate3394(.O (g7880), .I (g3201));
INVX1 gate3395(.O (g7888), .I (g1858));
INVX1 gate3396(.O (g7891), .I (g2010));
INVX1 gate3397(.O (g7892), .I (g2553));
INVX1 gate3398(.O (g7897), .I (g3047));
INVX1 gate3399(.O (g7898), .I (g3057));
INVX1 gate3400(.O (g7899), .I (g3066));
INVX1 gate3401(.O (g7900), .I (g3075));
INVX1 gate3402(.O (I15222), .I (g3151));
INVX1 gate3403(.O (g7901), .I (I15222));
INVX1 gate3404(.O (g7906), .I (g488));
INVX1 gate3405(.O (I15226), .I (g474));
INVX1 gate3406(.O (g7909), .I (I15226));
INVX1 gate3407(.O (g7910), .I (g474));
INVX1 gate3408(.O (I15230), .I (g499));
INVX1 gate3409(.O (g7911), .I (I15230));
INVX1 gate3410(.O (g7912), .I (g2552));
INVX1 gate3411(.O (g7915), .I (g2704));
INVX1 gate3412(.O (g7916), .I (g2935));
INVX1 gate3413(.O (g7919), .I (g2963));
INVX1 gate3414(.O (g7924), .I (g3048));
INVX1 gate3415(.O (g7925), .I (g3058));
INVX1 gate3416(.O (g7926), .I (g3067));
INVX1 gate3417(.O (g7927), .I (g3076));
INVX1 gate3418(.O (g7928), .I (g3204));
INVX1 gate3419(.O (I15256), .I (g2950));
INVX1 gate3420(.O (g7936), .I (I15256));
INVX1 gate3421(.O (g7949), .I (g165));
INVX1 gate3422(.O (g7950), .I (g142));
INVX1 gate3423(.O (g7953), .I (g487));
INVX1 gate3424(.O (I15262), .I (g481));
INVX1 gate3425(.O (g7956), .I (I15262));
INVX1 gate3426(.O (g7957), .I (g481));
INVX1 gate3427(.O (g7958), .I (g1175));
INVX1 gate3428(.O (I15267), .I (g1161));
INVX1 gate3429(.O (g7961), .I (I15267));
INVX1 gate3430(.O (g7962), .I (g1161));
INVX1 gate3431(.O (I15271), .I (g1186));
INVX1 gate3432(.O (g7963), .I (I15271));
INVX1 gate3433(.O (g7964), .I (g2938));
INVX1 gate3434(.O (g7967), .I (g2966));
INVX1 gate3435(.O (g7971), .I (g3049));
INVX1 gate3436(.O (g7972), .I (g3059));
INVX1 gate3437(.O (g7973), .I (g3068));
INVX1 gate3438(.O (g7974), .I (g3077));
INVX1 gate3439(.O (g7975), .I (g39));
INVX1 gate3440(.O (I15288), .I (g3109));
INVX1 gate3441(.O (g7976), .I (I15288));
INVX1 gate3442(.O (g7989), .I (g3191));
INVX1 gate3443(.O (g7990), .I (g143));
INVX1 gate3444(.O (g7993), .I (g145));
INVX1 gate3445(.O (g7996), .I (g486));
INVX1 gate3446(.O (g7999), .I (g485));
INVX1 gate3447(.O (g8000), .I (g853));
INVX1 gate3448(.O (g8001), .I (g830));
INVX1 gate3449(.O (g8004), .I (g1174));
INVX1 gate3450(.O (I15299), .I (g1168));
INVX1 gate3451(.O (g8007), .I (I15299));
INVX1 gate3452(.O (g8008), .I (g1168));
INVX1 gate3453(.O (g8009), .I (g1869));
INVX1 gate3454(.O (I15304), .I (g1855));
INVX1 gate3455(.O (g8012), .I (I15304));
INVX1 gate3456(.O (g8013), .I (g1855));
INVX1 gate3457(.O (I15308), .I (g1880));
INVX1 gate3458(.O (g8014), .I (I15308));
INVX1 gate3459(.O (g8015), .I (g2941));
INVX1 gate3460(.O (g8018), .I (g2969));
INVX1 gate3461(.O (I15313), .I (g2930));
INVX1 gate3462(.O (g8021), .I (I15313));
INVX1 gate3463(.O (g8022), .I (g2930));
INVX1 gate3464(.O (I15317), .I (g2842));
INVX1 gate3465(.O (g8023), .I (I15317));
INVX1 gate3466(.O (g8024), .I (g2842));
INVX1 gate3467(.O (g8025), .I (g3050));
INVX1 gate3468(.O (g8026), .I (g3060));
INVX1 gate3469(.O (g8027), .I (g3069));
INVX1 gate3470(.O (g8028), .I (g3078));
INVX1 gate3471(.O (g8029), .I (g3083));
INVX1 gate3472(.O (I15326), .I (g3117));
INVX1 gate3473(.O (g8030), .I (I15326));
INVX1 gate3474(.O (I15329), .I (g3117));
INVX1 gate3475(.O (g8031), .I (I15329));
INVX1 gate3476(.O (g8044), .I (g3194));
INVX1 gate3477(.O (g8045), .I (g3207));
INVX1 gate3478(.O (g8053), .I (g141));
INVX1 gate3479(.O (g8056), .I (g146));
INVX1 gate3480(.O (g8059), .I (g148));
INVX1 gate3481(.O (g8062), .I (g169));
INVX1 gate3482(.O (g8065), .I (g831));
INVX1 gate3483(.O (g8068), .I (g833));
INVX1 gate3484(.O (g8071), .I (g1173));
INVX1 gate3485(.O (g8074), .I (g1172));
INVX1 gate3486(.O (g8075), .I (g1547));
INVX1 gate3487(.O (g8076), .I (g1524));
INVX1 gate3488(.O (g8079), .I (g1868));
INVX1 gate3489(.O (I15345), .I (g1862));
INVX1 gate3490(.O (g8082), .I (I15345));
INVX1 gate3491(.O (g8083), .I (g1862));
INVX1 gate3492(.O (g8084), .I (g2563));
INVX1 gate3493(.O (I15350), .I (g2549));
INVX1 gate3494(.O (g8087), .I (I15350));
INVX1 gate3495(.O (g8088), .I (g2549));
INVX1 gate3496(.O (I15354), .I (g2574));
INVX1 gate3497(.O (g8089), .I (I15354));
INVX1 gate3498(.O (g8090), .I (g2944));
INVX1 gate3499(.O (g8093), .I (g2972));
INVX1 gate3500(.O (I15359), .I (g2858));
INVX1 gate3501(.O (g8096), .I (I15359));
INVX1 gate3502(.O (g8097), .I (g2858));
INVX1 gate3503(.O (g8098), .I (g3051));
INVX1 gate3504(.O (g8099), .I (g3061));
INVX1 gate3505(.O (g8100), .I (g3070));
INVX1 gate3506(.O (g8101), .I (g2997));
INVX1 gate3507(.O (g8102), .I (g27));
INVX1 gate3508(.O (g8103), .I (g185));
INVX1 gate3509(.O (I15369), .I (g3129));
INVX1 gate3510(.O (g8106), .I (I15369));
INVX1 gate3511(.O (I15372), .I (g3129));
INVX1 gate3512(.O (g8107), .I (I15372));
INVX1 gate3513(.O (g8120), .I (g3197));
INVX1 gate3514(.O (g8123), .I (g144));
INVX1 gate3515(.O (g8126), .I (g149));
INVX1 gate3516(.O (g8129), .I (g151));
INVX1 gate3517(.O (g8132), .I (g170));
INVX1 gate3518(.O (g8135), .I (g172));
INVX1 gate3519(.O (g8138), .I (g829));
INVX1 gate3520(.O (g8141), .I (g834));
INVX1 gate3521(.O (g8144), .I (g836));
INVX1 gate3522(.O (g8147), .I (g857));
INVX1 gate3523(.O (g8150), .I (g1525));
INVX1 gate3524(.O (g8153), .I (g1527));
INVX1 gate3525(.O (g8156), .I (g1867));
INVX1 gate3526(.O (g8159), .I (g1866));
INVX1 gate3527(.O (g8160), .I (g2241));
INVX1 gate3528(.O (g8161), .I (g2218));
INVX1 gate3529(.O (g8164), .I (g2562));
INVX1 gate3530(.O (I15392), .I (g2556));
INVX1 gate3531(.O (g8167), .I (I15392));
INVX1 gate3532(.O (g8168), .I (g2556));
INVX1 gate3533(.O (g8169), .I (g2947));
INVX1 gate3534(.O (g8172), .I (g2975));
INVX1 gate3535(.O (I15398), .I (g2845));
INVX1 gate3536(.O (g8175), .I (I15398));
INVX1 gate3537(.O (g8176), .I (g2845));
INVX1 gate3538(.O (g8177), .I (g3043));
INVX1 gate3539(.O (g8178), .I (g3052));
INVX1 gate3540(.O (g8179), .I (g3062));
INVX1 gate3541(.O (g8180), .I (g3071));
INVX1 gate3542(.O (g8181), .I (g48));
INVX1 gate3543(.O (g8182), .I (g3198));
INVX1 gate3544(.O (g8183), .I (g3188));
INVX1 gate3545(.O (g8191), .I (g147));
INVX1 gate3546(.O (g8194), .I (g152));
INVX1 gate3547(.O (g8197), .I (g154));
INVX1 gate3548(.O (g8200), .I (g168));
INVX1 gate3549(.O (g8203), .I (g173));
INVX1 gate3550(.O (g8206), .I (g175));
INVX1 gate3551(.O (g8209), .I (g832));
INVX1 gate3552(.O (g8212), .I (g837));
INVX1 gate3553(.O (g8215), .I (g839));
INVX1 gate3554(.O (g8218), .I (g858));
INVX1 gate3555(.O (g8221), .I (g860));
INVX1 gate3556(.O (g8224), .I (g1523));
INVX1 gate3557(.O (g8227), .I (g1528));
INVX1 gate3558(.O (g8230), .I (g1530));
INVX1 gate3559(.O (g8233), .I (g1551));
INVX1 gate3560(.O (g8236), .I (g2219));
INVX1 gate3561(.O (g8239), .I (g2221));
INVX1 gate3562(.O (g8242), .I (g2561));
INVX1 gate3563(.O (g8245), .I (g2560));
INVX1 gate3564(.O (g8246), .I (g2978));
INVX1 gate3565(.O (I15429), .I (g2833));
INVX1 gate3566(.O (g8249), .I (I15429));
INVX1 gate3567(.O (g8250), .I (g2833));
INVX1 gate3568(.O (I15433), .I (g2861));
INVX1 gate3569(.O (g8251), .I (I15433));
INVX1 gate3570(.O (g8252), .I (g2861));
INVX1 gate3571(.O (g8253), .I (g3053));
INVX1 gate3572(.O (g8254), .I (g3063));
INVX1 gate3573(.O (g8255), .I (g3072));
INVX1 gate3574(.O (g8256), .I (g30));
INVX1 gate3575(.O (g8257), .I (g3201));
INVX1 gate3576(.O (I15442), .I (g3235));
INVX1 gate3577(.O (g8258), .I (I15442));
INVX1 gate3578(.O (I15445), .I (g3236));
INVX1 gate3579(.O (g8259), .I (I15445));
INVX1 gate3580(.O (I15448), .I (g3237));
INVX1 gate3581(.O (g8260), .I (I15448));
INVX1 gate3582(.O (I15451), .I (g3238));
INVX1 gate3583(.O (g8261), .I (I15451));
INVX1 gate3584(.O (I15454), .I (g3239));
INVX1 gate3585(.O (g8262), .I (I15454));
INVX1 gate3586(.O (I15457), .I (g3240));
INVX1 gate3587(.O (g8263), .I (I15457));
INVX1 gate3588(.O (I15460), .I (g3241));
INVX1 gate3589(.O (g8264), .I (I15460));
INVX1 gate3590(.O (I15463), .I (g3242));
INVX1 gate3591(.O (g8265), .I (I15463));
INVX1 gate3592(.O (I15466), .I (g3243));
INVX1 gate3593(.O (g8266), .I (I15466));
INVX1 gate3594(.O (I15469), .I (g3244));
INVX1 gate3595(.O (g8267), .I (I15469));
INVX1 gate3596(.O (I15472), .I (g3245));
INVX1 gate3597(.O (g8268), .I (I15472));
INVX1 gate3598(.O (I15475), .I (g3246));
INVX1 gate3599(.O (g8269), .I (I15475));
INVX1 gate3600(.O (I15478), .I (g3247));
INVX1 gate3601(.O (g8270), .I (I15478));
INVX1 gate3602(.O (I15481), .I (g3248));
INVX1 gate3603(.O (g8271), .I (I15481));
INVX1 gate3604(.O (I15484), .I (g3249));
INVX1 gate3605(.O (g8272), .I (I15484));
INVX1 gate3606(.O (I15487), .I (g3250));
INVX1 gate3607(.O (g8273), .I (I15487));
INVX1 gate3608(.O (I15490), .I (g3251));
INVX1 gate3609(.O (g8274), .I (I15490));
INVX1 gate3610(.O (I15493), .I (g3252));
INVX1 gate3611(.O (g8275), .I (I15493));
INVX1 gate3612(.O (g8276), .I (g3253));
INVX1 gate3613(.O (g8277), .I (g3305));
INVX1 gate3614(.O (g8278), .I (g3337));
INVX1 gate3615(.O (I15499), .I (g7911));
INVX1 gate3616(.O (g8284), .I (I15499));
INVX1 gate3617(.O (g8285), .I (g3365));
INVX1 gate3618(.O (g8286), .I (g3461));
INVX1 gate3619(.O (g8287), .I (g3493));
INVX1 gate3620(.O (I15505), .I (g7963));
INVX1 gate3621(.O (g8293), .I (I15505));
INVX1 gate3622(.O (g8294), .I (g3521));
INVX1 gate3623(.O (g8295), .I (g3617));
INVX1 gate3624(.O (g8296), .I (g3649));
INVX1 gate3625(.O (I15511), .I (g8014));
INVX1 gate3626(.O (g8302), .I (I15511));
INVX1 gate3627(.O (g8303), .I (g3677));
INVX1 gate3628(.O (g8304), .I (g3773));
INVX1 gate3629(.O (g8305), .I (g3805));
INVX1 gate3630(.O (I15517), .I (g8089));
INVX1 gate3631(.O (g8311), .I (I15517));
INVX1 gate3632(.O (g8312), .I (g3833));
INVX1 gate3633(.O (g8313), .I (g3897));
INVX1 gate3634(.O (g8317), .I (g3919));
INVX1 gate3635(.O (I15523), .I (g3254));
INVX1 gate3636(.O (g8321), .I (I15523));
INVX1 gate3637(.O (I15526), .I (g6314));
INVX1 gate3638(.O (g8324), .I (I15526));
INVX1 gate3639(.O (I15532), .I (g3410));
INVX1 gate3640(.O (g8330), .I (I15532));
INVX1 gate3641(.O (I15535), .I (g6519));
INVX1 gate3642(.O (g8333), .I (I15535));
INVX1 gate3643(.O (I15538), .I (g6369));
INVX1 gate3644(.O (g8336), .I (I15538));
INVX1 gate3645(.O (I15543), .I (g3410));
INVX1 gate3646(.O (g8341), .I (I15543));
INVX1 gate3647(.O (I15546), .I (g6783));
INVX1 gate3648(.O (g8344), .I (I15546));
INVX1 gate3649(.O (I15549), .I (g6574));
INVX1 gate3650(.O (g8347), .I (I15549));
INVX1 gate3651(.O (I15553), .I (g3566));
INVX1 gate3652(.O (g8351), .I (I15553));
INVX1 gate3653(.O (I15556), .I (g6783));
INVX1 gate3654(.O (g8354), .I (I15556));
INVX1 gate3655(.O (I15559), .I (g7015));
INVX1 gate3656(.O (g8357), .I (I15559));
INVX1 gate3657(.O (I15562), .I (g5778));
INVX1 gate3658(.O (g8360), .I (I15562));
INVX1 gate3659(.O (I15565), .I (g6838));
INVX1 gate3660(.O (g8363), .I (I15565));
INVX1 gate3661(.O (I15568), .I (g3722));
INVX1 gate3662(.O (g8366), .I (I15568));
INVX1 gate3663(.O (I15571), .I (g7085));
INVX1 gate3664(.O (g8369), .I (I15571));
INVX1 gate3665(.O (I15574), .I (g6838));
INVX1 gate3666(.O (g8372), .I (I15574));
INVX1 gate3667(.O (I15577), .I (g7265));
INVX1 gate3668(.O (g8375), .I (I15577));
INVX1 gate3669(.O (I15580), .I (g5837));
INVX1 gate3670(.O (g8378), .I (I15580));
INVX1 gate3671(.O (I15584), .I (g3254));
INVX1 gate3672(.O (g8382), .I (I15584));
INVX1 gate3673(.O (I15590), .I (g3410));
INVX1 gate3674(.O (g8388), .I (I15590));
INVX1 gate3675(.O (I15593), .I (g6519));
INVX1 gate3676(.O (g8391), .I (I15593));
INVX1 gate3677(.O (I15599), .I (g3566));
INVX1 gate3678(.O (g8397), .I (I15599));
INVX1 gate3679(.O (I15602), .I (g6783));
INVX1 gate3680(.O (g8400), .I (I15602));
INVX1 gate3681(.O (I15605), .I (g6574));
INVX1 gate3682(.O (g8403), .I (I15605));
INVX1 gate3683(.O (I15610), .I (g3566));
INVX1 gate3684(.O (g8408), .I (I15610));
INVX1 gate3685(.O (I15613), .I (g7085));
INVX1 gate3686(.O (g8411), .I (I15613));
INVX1 gate3687(.O (I15616), .I (g6838));
INVX1 gate3688(.O (g8414), .I (I15616));
INVX1 gate3689(.O (I15620), .I (g3722));
INVX1 gate3690(.O (g8418), .I (I15620));
INVX1 gate3691(.O (I15623), .I (g7085));
INVX1 gate3692(.O (g8421), .I (I15623));
INVX1 gate3693(.O (I15626), .I (g7265));
INVX1 gate3694(.O (g8424), .I (I15626));
INVX1 gate3695(.O (I15629), .I (g5837));
INVX1 gate3696(.O (g8427), .I (I15629));
INVX1 gate3697(.O (I15636), .I (g3410));
INVX1 gate3698(.O (g8434), .I (I15636));
INVX1 gate3699(.O (I15642), .I (g3566));
INVX1 gate3700(.O (g8440), .I (I15642));
INVX1 gate3701(.O (I15645), .I (g6783));
INVX1 gate3702(.O (g8443), .I (I15645));
INVX1 gate3703(.O (I15651), .I (g3722));
INVX1 gate3704(.O (g8449), .I (I15651));
INVX1 gate3705(.O (I15654), .I (g7085));
INVX1 gate3706(.O (g8452), .I (I15654));
INVX1 gate3707(.O (I15657), .I (g6838));
INVX1 gate3708(.O (g8455), .I (I15657));
INVX1 gate3709(.O (I15662), .I (g3722));
INVX1 gate3710(.O (g8460), .I (I15662));
INVX1 gate3711(.O (I15671), .I (g3566));
INVX1 gate3712(.O (g8469), .I (I15671));
INVX1 gate3713(.O (I15677), .I (g3722));
INVX1 gate3714(.O (g8475), .I (I15677));
INVX1 gate3715(.O (I15680), .I (g7085));
INVX1 gate3716(.O (g8478), .I (I15680));
INVX1 gate3717(.O (I15696), .I (g3722));
INVX1 gate3718(.O (g8494), .I (I15696));
INVX1 gate3719(.O (g8514), .I (g6139));
INVX1 gate3720(.O (g8530), .I (g6156));
INVX1 gate3721(.O (g8568), .I (g6230));
INVX1 gate3722(.O (I15771), .I (g6000));
INVX1 gate3723(.O (g8569), .I (I15771));
INVX1 gate3724(.O (I15779), .I (g6000));
INVX1 gate3725(.O (g8575), .I (I15779));
INVX1 gate3726(.O (I15784), .I (g6000));
INVX1 gate3727(.O (g8578), .I (I15784));
INVX1 gate3728(.O (I15787), .I (g6000));
INVX1 gate3729(.O (g8579), .I (I15787));
INVX1 gate3730(.O (g8580), .I (g6281));
INVX1 gate3731(.O (g8587), .I (g6418));
INVX1 gate3732(.O (g8594), .I (g6623));
INVX1 gate3733(.O (I15794), .I (g3338));
INVX1 gate3734(.O (g8602), .I (I15794));
INVX1 gate3735(.O (g8605), .I (g6887));
INVX1 gate3736(.O (I15800), .I (g3494));
INVX1 gate3737(.O (g8614), .I (I15800));
INVX1 gate3738(.O (I15803), .I (g8107));
INVX1 gate3739(.O (g8617), .I (I15803));
INVX1 gate3740(.O (I15806), .I (g5550));
INVX1 gate3741(.O (g8620), .I (I15806));
INVX1 gate3742(.O (I15810), .I (g3338));
INVX1 gate3743(.O (g8622), .I (I15810));
INVX1 gate3744(.O (I15815), .I (g3650));
INVX1 gate3745(.O (g8627), .I (I15815));
INVX1 gate3746(.O (I15818), .I (g5596));
INVX1 gate3747(.O (g8630), .I (I15818));
INVX1 gate3748(.O (I15822), .I (g3494));
INVX1 gate3749(.O (g8632), .I (I15822));
INVX1 gate3750(.O (I15827), .I (g3806));
INVX1 gate3751(.O (g8637), .I (I15827));
INVX1 gate3752(.O (I15830), .I (g8031));
INVX1 gate3753(.O (g8640), .I (I15830));
INVX1 gate3754(.O (I15833), .I (g3338));
INVX1 gate3755(.O (g8643), .I (I15833));
INVX1 gate3756(.O (I15836), .I (g3366));
INVX1 gate3757(.O (g8646), .I (I15836));
INVX1 gate3758(.O (I15839), .I (g5613));
INVX1 gate3759(.O (g8649), .I (I15839));
INVX1 gate3760(.O (I15843), .I (g3650));
INVX1 gate3761(.O (g8651), .I (I15843));
INVX1 gate3762(.O (I15847), .I (g3878));
INVX1 gate3763(.O (g8655), .I (I15847));
INVX1 gate3764(.O (I15850), .I (g5627));
INVX1 gate3765(.O (g8658), .I (I15850));
INVX1 gate3766(.O (I15853), .I (g3494));
INVX1 gate3767(.O (g8659), .I (I15853));
INVX1 gate3768(.O (I15856), .I (g3522));
INVX1 gate3769(.O (g8662), .I (I15856));
INVX1 gate3770(.O (I15859), .I (g5638));
INVX1 gate3771(.O (g8665), .I (I15859));
INVX1 gate3772(.O (I15863), .I (g3806));
INVX1 gate3773(.O (g8667), .I (I15863));
INVX1 gate3774(.O (I15866), .I (g3878));
INVX1 gate3775(.O (g8670), .I (I15866));
INVX1 gate3776(.O (I15869), .I (g7976));
INVX1 gate3777(.O (g8673), .I (I15869));
INVX1 gate3778(.O (I15873), .I (g5655));
INVX1 gate3779(.O (g8677), .I (I15873));
INVX1 gate3780(.O (I15876), .I (g3650));
INVX1 gate3781(.O (g8678), .I (I15876));
INVX1 gate3782(.O (I15879), .I (g3678));
INVX1 gate3783(.O (g8681), .I (I15879));
INVX1 gate3784(.O (I15882), .I (g3878));
INVX1 gate3785(.O (g8684), .I (I15882));
INVX1 gate3786(.O (I15887), .I (g5693));
INVX1 gate3787(.O (g8689), .I (I15887));
INVX1 gate3788(.O (I15890), .I (g3806));
INVX1 gate3789(.O (g8690), .I (I15890));
INVX1 gate3790(.O (I15893), .I (g3834));
INVX1 gate3791(.O (g8693), .I (I15893));
INVX1 gate3792(.O (I15896), .I (g3878));
INVX1 gate3793(.O (g8696), .I (I15896));
INVX1 gate3794(.O (I15899), .I (g5626));
INVX1 gate3795(.O (g8699), .I (I15899));
INVX1 gate3796(.O (I15902), .I (g6486));
INVX1 gate3797(.O (g8700), .I (I15902));
INVX1 gate3798(.O (I15909), .I (g5745));
INVX1 gate3799(.O (g8707), .I (I15909));
INVX1 gate3800(.O (I15912), .I (g3878));
INVX1 gate3801(.O (g8708), .I (I15912));
INVX1 gate3802(.O (I15915), .I (g3878));
INVX1 gate3803(.O (g8711), .I (I15915));
INVX1 gate3804(.O (I15918), .I (g6643));
INVX1 gate3805(.O (g8714), .I (I15918));
INVX1 gate3806(.O (I15922), .I (g5654));
INVX1 gate3807(.O (g8718), .I (I15922));
INVX1 gate3808(.O (I15925), .I (g6751));
INVX1 gate3809(.O (g8719), .I (I15925));
INVX1 gate3810(.O (I15932), .I (g5423));
INVX1 gate3811(.O (g8726), .I (I15932));
INVX1 gate3812(.O (I15935), .I (g3878));
INVX1 gate3813(.O (g8745), .I (I15935));
INVX1 gate3814(.O (I15938), .I (g3338));
INVX1 gate3815(.O (g8748), .I (I15938));
INVX1 gate3816(.O (I15942), .I (g6945));
INVX1 gate3817(.O (g8752), .I (I15942));
INVX1 gate3818(.O (I15946), .I (g5692));
INVX1 gate3819(.O (g8756), .I (I15946));
INVX1 gate3820(.O (I15949), .I (g7053));
INVX1 gate3821(.O (g8757), .I (I15949));
INVX1 gate3822(.O (I15955), .I (g3878));
INVX1 gate3823(.O (g8763), .I (I15955));
INVX1 gate3824(.O (I15958), .I (g3878));
INVX1 gate3825(.O (g8766), .I (I15958));
INVX1 gate3826(.O (I15961), .I (g6051));
INVX1 gate3827(.O (g8769), .I (I15961));
INVX1 gate3828(.O (I15964), .I (g7554));
INVX1 gate3829(.O (g8770), .I (I15964));
INVX1 gate3830(.O (I15967), .I (g3494));
INVX1 gate3831(.O (g8771), .I (I15967));
INVX1 gate3832(.O (I15971), .I (g7195));
INVX1 gate3833(.O (g8775), .I (I15971));
INVX1 gate3834(.O (I15975), .I (g5744));
INVX1 gate3835(.O (g8779), .I (I15975));
INVX1 gate3836(.O (I15978), .I (g7303));
INVX1 gate3837(.O (g8780), .I (I15978));
INVX1 gate3838(.O (I15983), .I (g3878));
INVX1 gate3839(.O (g8785), .I (I15983));
INVX1 gate3840(.O (I15986), .I (g3878));
INVX1 gate3841(.O (g8788), .I (I15986));
INVX1 gate3842(.O (I15989), .I (g6053));
INVX1 gate3843(.O (g8791), .I (I15989));
INVX1 gate3844(.O (I15992), .I (g6055));
INVX1 gate3845(.O (g8792), .I (I15992));
INVX1 gate3846(.O (I15995), .I (g7577));
INVX1 gate3847(.O (g8793), .I (I15995));
INVX1 gate3848(.O (I15998), .I (g3650));
INVX1 gate3849(.O (g8794), .I (I15998));
INVX1 gate3850(.O (I16002), .I (g7391));
INVX1 gate3851(.O (g8798), .I (I16002));
INVX1 gate3852(.O (I16006), .I (g3878));
INVX1 gate3853(.O (g8802), .I (I16006));
INVX1 gate3854(.O (I16009), .I (g3878));
INVX1 gate3855(.O (g8805), .I (I16009));
INVX1 gate3856(.O (I16012), .I (g5390));
INVX1 gate3857(.O (g8808), .I (I16012));
INVX1 gate3858(.O (I16015), .I (g6056));
INVX1 gate3859(.O (g8809), .I (I16015));
INVX1 gate3860(.O (I16018), .I (g6058));
INVX1 gate3861(.O (g8810), .I (I16018));
INVX1 gate3862(.O (I16021), .I (g6060));
INVX1 gate3863(.O (g8811), .I (I16021));
INVX1 gate3864(.O (I16024), .I (g7591));
INVX1 gate3865(.O (g8812), .I (I16024));
INVX1 gate3866(.O (I16027), .I (g3806));
INVX1 gate3867(.O (g8813), .I (I16027));
INVX1 gate3868(.O (I16031), .I (g3878));
INVX1 gate3869(.O (g8817), .I (I16031));
INVX1 gate3870(.O (I16034), .I (g5396));
INVX1 gate3871(.O (g8820), .I (I16034));
INVX1 gate3872(.O (I16037), .I (g6061));
INVX1 gate3873(.O (g8821), .I (I16037));
INVX1 gate3874(.O (g8822), .I (g4602));
INVX1 gate3875(.O (I16041), .I (g6486));
INVX1 gate3876(.O (g8823), .I (I16041));
INVX1 gate3877(.O (I16044), .I (g5397));
INVX1 gate3878(.O (g8824), .I (I16044));
INVX1 gate3879(.O (I16047), .I (g6063));
INVX1 gate3880(.O (g8825), .I (I16047));
INVX1 gate3881(.O (I16050), .I (g6065));
INVX1 gate3882(.O (g8826), .I (I16050));
INVX1 gate3883(.O (I16053), .I (g6067));
INVX1 gate3884(.O (g8827), .I (I16053));
INVX1 gate3885(.O (I16056), .I (g7606));
INVX1 gate3886(.O (g8828), .I (I16056));
INVX1 gate3887(.O (I16059), .I (g3878));
INVX1 gate3888(.O (g8829), .I (I16059));
INVX1 gate3889(.O (I16062), .I (g3900));
INVX1 gate3890(.O (g8832), .I (I16062));
INVX1 gate3891(.O (I16065), .I (g7936));
INVX1 gate3892(.O (g8835), .I (I16065));
INVX1 gate3893(.O (I16068), .I (g5438));
INVX1 gate3894(.O (g8836), .I (I16068));
INVX1 gate3895(.O (I16071), .I (g5395));
INVX1 gate3896(.O (g8839), .I (I16071));
INVX1 gate3897(.O (I16074), .I (g5399));
INVX1 gate3898(.O (g8840), .I (I16074));
INVX1 gate3899(.O (I16079), .I (g6086));
INVX1 gate3900(.O (g8843), .I (I16079));
INVX1 gate3901(.O (I16082), .I (g5401));
INVX1 gate3902(.O (g8844), .I (I16082));
INVX1 gate3903(.O (I16085), .I (g6080));
INVX1 gate3904(.O (g8845), .I (I16085));
INVX1 gate3905(.O (g8846), .I (g4779));
INVX1 gate3906(.O (I16089), .I (g6751));
INVX1 gate3907(.O (g8847), .I (I16089));
INVX1 gate3908(.O (I16092), .I (g5402));
INVX1 gate3909(.O (g8850), .I (I16092));
INVX1 gate3910(.O (I16095), .I (g6082));
INVX1 gate3911(.O (g8851), .I (I16095));
INVX1 gate3912(.O (I16098), .I (g6084));
INVX1 gate3913(.O (g8852), .I (I16098));
INVX1 gate3914(.O (I16101), .I (g3878));
INVX1 gate3915(.O (g8853), .I (I16101));
INVX1 gate3916(.O (I16104), .I (g6448));
INVX1 gate3917(.O (g8856), .I (I16104));
INVX1 gate3918(.O (I16107), .I (g5398));
INVX1 gate3919(.O (g8859), .I (I16107));
INVX1 gate3920(.O (I16110), .I (g5404));
INVX1 gate3921(.O (g8860), .I (I16110));
INVX1 gate3922(.O (I16114), .I (g7936));
INVX1 gate3923(.O (g8862), .I (I16114));
INVX1 gate3924(.O (I16117), .I (g5473));
INVX1 gate3925(.O (g8863), .I (I16117));
INVX1 gate3926(.O (I16120), .I (g5400));
INVX1 gate3927(.O (g8866), .I (I16120));
INVX1 gate3928(.O (I16123), .I (g5406));
INVX1 gate3929(.O (g8867), .I (I16123));
INVX1 gate3930(.O (I16128), .I (g6103));
INVX1 gate3931(.O (g8870), .I (I16128));
INVX1 gate3932(.O (I16131), .I (g5408));
INVX1 gate3933(.O (g8871), .I (I16131));
INVX1 gate3934(.O (I16134), .I (g6099));
INVX1 gate3935(.O (g8872), .I (I16134));
INVX1 gate3936(.O (g8873), .I (g4955));
INVX1 gate3937(.O (I16138), .I (g7053));
INVX1 gate3938(.O (g8874), .I (I16138));
INVX1 gate3939(.O (I16141), .I (g5409));
INVX1 gate3940(.O (g8877), .I (I16141));
INVX1 gate3941(.O (I16144), .I (g6101));
INVX1 gate3942(.O (g8878), .I (I16144));
INVX1 gate3943(.O (I16147), .I (g3878));
INVX1 gate3944(.O (g8879), .I (I16147));
INVX1 gate3945(.O (I16150), .I (g3900));
INVX1 gate3946(.O (g8882), .I (I16150));
INVX1 gate3947(.O (I16153), .I (g3306));
INVX1 gate3948(.O (g8885), .I (I16153));
INVX1 gate3949(.O (I16156), .I (g5438));
INVX1 gate3950(.O (g8888), .I (I16156));
INVX1 gate3951(.O (I16159), .I (g5403));
INVX1 gate3952(.O (g8891), .I (I16159));
INVX1 gate3953(.O (I16163), .I (g6031));
INVX1 gate3954(.O (g8893), .I (I16163));
INVX1 gate3955(.O (I16166), .I (g6713));
INVX1 gate3956(.O (g8894), .I (I16166));
INVX1 gate3957(.O (I16169), .I (g5405));
INVX1 gate3958(.O (g8897), .I (I16169));
INVX1 gate3959(.O (I16172), .I (g5413));
INVX1 gate3960(.O (g8898), .I (I16172));
INVX1 gate3961(.O (I16176), .I (g7936));
INVX1 gate3962(.O (g8900), .I (I16176));
INVX1 gate3963(.O (I16179), .I (g5512));
INVX1 gate3964(.O (g8901), .I (I16179));
INVX1 gate3965(.O (I16182), .I (g5407));
INVX1 gate3966(.O (g8904), .I (I16182));
INVX1 gate3967(.O (I16185), .I (g5415));
INVX1 gate3968(.O (g8905), .I (I16185));
INVX1 gate3969(.O (I16190), .I (g6118));
INVX1 gate3970(.O (g8908), .I (I16190));
INVX1 gate3971(.O (I16193), .I (g5417));
INVX1 gate3972(.O (g8909), .I (I16193));
INVX1 gate3973(.O (I16196), .I (g6116));
INVX1 gate3974(.O (g8910), .I (I16196));
INVX1 gate3975(.O (g8911), .I (g5114));
INVX1 gate3976(.O (I16200), .I (g7303));
INVX1 gate3977(.O (g8912), .I (I16200));
INVX1 gate3978(.O (I16203), .I (g3878));
INVX1 gate3979(.O (g8915), .I (I16203));
INVX1 gate3980(.O (I16206), .I (g6448));
INVX1 gate3981(.O (g8918), .I (I16206));
INVX1 gate3982(.O (I16209), .I (g5438));
INVX1 gate3983(.O (g8921), .I (I16209));
INVX1 gate3984(.O (I16212), .I (g5411));
INVX1 gate3985(.O (g8924), .I (I16212));
INVX1 gate3986(.O (I16215), .I (g3462));
INVX1 gate3987(.O (g8925), .I (I16215));
INVX1 gate3988(.O (I16218), .I (g5473));
INVX1 gate3989(.O (g8928), .I (I16218));
INVX1 gate3990(.O (I16221), .I (g5412));
INVX1 gate3991(.O (g8931), .I (I16221));
INVX1 gate3992(.O (I16225), .I (g6042));
INVX1 gate3993(.O (g8933), .I (I16225));
INVX1 gate3994(.O (I16228), .I (g7015));
INVX1 gate3995(.O (g8934), .I (I16228));
INVX1 gate3996(.O (I16231), .I (g5414));
INVX1 gate3997(.O (g8937), .I (I16231));
INVX1 gate3998(.O (I16234), .I (g5420));
INVX1 gate3999(.O (g8938), .I (I16234));
INVX1 gate4000(.O (I16238), .I (g7936));
INVX1 gate4001(.O (g8940), .I (I16238));
INVX1 gate4002(.O (I16241), .I (g5556));
INVX1 gate4003(.O (g8941), .I (I16241));
INVX1 gate4004(.O (I16244), .I (g5416));
INVX1 gate4005(.O (g8944), .I (I16244));
INVX1 gate4006(.O (I16247), .I (g5422));
INVX1 gate4007(.O (g8945), .I (I16247));
INVX1 gate4008(.O (I16252), .I (g6134));
INVX1 gate4009(.O (g8948), .I (I16252));
INVX1 gate4010(.O (I16255), .I (g3900));
INVX1 gate4011(.O (g8949), .I (I16255));
INVX1 gate4012(.O (I16258), .I (g3306));
INVX1 gate4013(.O (g8952), .I (I16258));
INVX1 gate4014(.O (I16261), .I (g6448));
INVX1 gate4015(.O (g8955), .I (I16261));
INVX1 gate4016(.O (I16264), .I (g6713));
INVX1 gate4017(.O (g8958), .I (I16264));
INVX1 gate4018(.O (I16267), .I (g5473));
INVX1 gate4019(.O (g8961), .I (I16267));
INVX1 gate4020(.O (I16270), .I (g5418));
INVX1 gate4021(.O (g8964), .I (I16270));
INVX1 gate4022(.O (I16273), .I (g3618));
INVX1 gate4023(.O (g8965), .I (I16273));
INVX1 gate4024(.O (I16276), .I (g5512));
INVX1 gate4025(.O (g8968), .I (I16276));
INVX1 gate4026(.O (I16279), .I (g5419));
INVX1 gate4027(.O (g8971), .I (I16279));
INVX1 gate4028(.O (I16283), .I (g6046));
INVX1 gate4029(.O (g8973), .I (I16283));
INVX1 gate4030(.O (I16286), .I (g7265));
INVX1 gate4031(.O (g8974), .I (I16286));
INVX1 gate4032(.O (I16289), .I (g5421));
INVX1 gate4033(.O (g8977), .I (I16289));
INVX1 gate4034(.O (I16292), .I (g5426));
INVX1 gate4035(.O (g8978), .I (I16292));
INVX1 gate4036(.O (I16296), .I (g3306));
INVX1 gate4037(.O (g8980), .I (I16296));
INVX1 gate4038(.O (g8983), .I (g6486));
INVX1 gate4039(.O (I16300), .I (g3462));
INVX1 gate4040(.O (g8984), .I (I16300));
INVX1 gate4041(.O (I16303), .I (g6713));
INVX1 gate4042(.O (g8987), .I (I16303));
INVX1 gate4043(.O (I16306), .I (g7015));
INVX1 gate4044(.O (g8990), .I (I16306));
INVX1 gate4045(.O (I16309), .I (g5512));
INVX1 gate4046(.O (g8993), .I (I16309));
INVX1 gate4047(.O (I16312), .I (g5424));
INVX1 gate4048(.O (g8996), .I (I16312));
INVX1 gate4049(.O (I16315), .I (g3774));
INVX1 gate4050(.O (g8997), .I (I16315));
INVX1 gate4051(.O (I16318), .I (g5556));
INVX1 gate4052(.O (g9000), .I (I16318));
INVX1 gate4053(.O (I16321), .I (g5425));
INVX1 gate4054(.O (g9003), .I (I16321));
INVX1 gate4055(.O (I16325), .I (g6052));
INVX1 gate4056(.O (g9005), .I (I16325));
INVX1 gate4057(.O (I16328), .I (g3900));
INVX1 gate4058(.O (g9006), .I (I16328));
INVX1 gate4059(.O (I16332), .I (g3462));
INVX1 gate4060(.O (g9010), .I (I16332));
INVX1 gate4061(.O (I16335), .I (g3618));
INVX1 gate4062(.O (g9013), .I (I16335));
INVX1 gate4063(.O (I16338), .I (g7015));
INVX1 gate4064(.O (g9016), .I (I16338));
INVX1 gate4065(.O (I16341), .I (g7265));
INVX1 gate4066(.O (g9019), .I (I16341));
INVX1 gate4067(.O (I16344), .I (g5556));
INVX1 gate4068(.O (g9022), .I (I16344));
INVX1 gate4069(.O (I16347), .I (g5427));
INVX1 gate4070(.O (g9025), .I (I16347));
INVX1 gate4071(.O (g9027), .I (g5679));
INVX1 gate4072(.O (I16354), .I (g3618));
INVX1 gate4073(.O (g9035), .I (I16354));
INVX1 gate4074(.O (I16357), .I (g3774));
INVX1 gate4075(.O (g9038), .I (I16357));
INVX1 gate4076(.O (I16360), .I (g7265));
INVX1 gate4077(.O (g9041), .I (I16360));
INVX1 gate4078(.O (I16363), .I (g3900));
INVX1 gate4079(.O (g9044), .I (I16363));
INVX1 gate4080(.O (g9050), .I (g5731));
INVX1 gate4081(.O (I16372), .I (g3774));
INVX1 gate4082(.O (g9058), .I (I16372));
INVX1 gate4083(.O (g9067), .I (g5789));
INVX1 gate4084(.O (g9084), .I (g5848));
INVX1 gate4085(.O (I16432), .I (g3366));
INVX1 gate4086(.O (g9128), .I (I16432));
INVX1 gate4087(.O (I16438), .I (g3522));
INVX1 gate4088(.O (g9134), .I (I16438));
INVX1 gate4089(.O (I16444), .I (g3678));
INVX1 gate4090(.O (g9140), .I (I16444));
INVX1 gate4091(.O (I16450), .I (g3834));
INVX1 gate4092(.O (g9146), .I (I16450));
INVX1 gate4093(.O (I16453), .I (g7936));
INVX1 gate4094(.O (g9149), .I (I16453));
INVX1 gate4095(.O (g9150), .I (g5893));
INVX1 gate4096(.O (I16457), .I (g7936));
INVX1 gate4097(.O (g9159), .I (I16457));
INVX1 gate4098(.O (g9160), .I (g6170));
INVX1 gate4099(.O (g9161), .I (g5852));
INVX1 gate4100(.O (I16462), .I (g5438));
INVX1 gate4101(.O (g9170), .I (I16462));
INVX1 gate4102(.O (I16465), .I (g6000));
INVX1 gate4103(.O (g9173), .I (I16465));
INVX1 gate4104(.O (g9174), .I (g5932));
INVX1 gate4105(.O (I16469), .I (g7936));
INVX1 gate4106(.O (g9183), .I (I16469));
INVX1 gate4107(.O (I16472), .I (g7901));
INVX1 gate4108(.O (g9184), .I (I16472));
INVX1 gate4109(.O (g9187), .I (g5803));
INVX1 gate4110(.O (I16476), .I (g6448));
INVX1 gate4111(.O (g9196), .I (I16476));
INVX1 gate4112(.O (I16479), .I (g5438));
INVX1 gate4113(.O (g9199), .I (I16479));
INVX1 gate4114(.O (I16482), .I (g6000));
INVX1 gate4115(.O (g9202), .I (I16482));
INVX1 gate4116(.O (g9203), .I (g5899));
INVX1 gate4117(.O (I16486), .I (g5473));
INVX1 gate4118(.O (g9212), .I (I16486));
INVX1 gate4119(.O (I16489), .I (g6000));
INVX1 gate4120(.O (g9215), .I (I16489));
INVX1 gate4121(.O (g9216), .I (g5966));
INVX1 gate4122(.O (I16493), .I (g7936));
INVX1 gate4123(.O (g9225), .I (I16493));
INVX1 gate4124(.O (g9226), .I (g5434));
INVX1 gate4125(.O (g9227), .I (g5587));
INVX1 gate4126(.O (g9228), .I (g7667));
INVX1 gate4127(.O (I16499), .I (g7901));
INVX1 gate4128(.O (g9229), .I (I16499));
INVX1 gate4129(.O (g9232), .I (g5752));
INVX1 gate4130(.O (I16504), .I (g3306));
INVX1 gate4131(.O (g9242), .I (I16504));
INVX1 gate4132(.O (I16507), .I (g6448));
INVX1 gate4133(.O (g9245), .I (I16507));
INVX1 gate4134(.O (g9248), .I (g5859));
INVX1 gate4135(.O (I16511), .I (g6713));
INVX1 gate4136(.O (g9257), .I (I16511));
INVX1 gate4137(.O (I16514), .I (g5473));
INVX1 gate4138(.O (g9260), .I (I16514));
INVX1 gate4139(.O (I16517), .I (g6000));
INVX1 gate4140(.O (g9263), .I (I16517));
INVX1 gate4141(.O (g9264), .I (g5938));
INVX1 gate4142(.O (I16521), .I (g5512));
INVX1 gate4143(.O (g9273), .I (I16521));
INVX1 gate4144(.O (I16524), .I (g6000));
INVX1 gate4145(.O (g9276), .I (I16524));
INVX1 gate4146(.O (g9277), .I (g5995));
INVX1 gate4147(.O (g9286), .I (g6197));
INVX1 gate4148(.O (g9287), .I (g6638));
INVX1 gate4149(.O (g9288), .I (g5363));
INVX1 gate4150(.O (g9289), .I (g5379));
INVX1 gate4151(.O (I16532), .I (g7901));
INVX1 gate4152(.O (g9290), .I (I16532));
INVX1 gate4153(.O (g9293), .I (g5703));
INVX1 gate4154(.O (I16538), .I (g3306));
INVX1 gate4155(.O (g9303), .I (I16538));
INVX1 gate4156(.O (I16541), .I (g5438));
INVX1 gate4157(.O (g9306), .I (I16541));
INVX1 gate4158(.O (I16544), .I (g6054));
INVX1 gate4159(.O (g9309), .I (I16544));
INVX1 gate4160(.O (g9310), .I (g5811));
INVX1 gate4161(.O (I16549), .I (g3462));
INVX1 gate4162(.O (g9320), .I (I16549));
INVX1 gate4163(.O (I16552), .I (g6713));
INVX1 gate4164(.O (g9323), .I (I16552));
INVX1 gate4165(.O (g9326), .I (g5906));
INVX1 gate4166(.O (I16556), .I (g7015));
INVX1 gate4167(.O (g9335), .I (I16556));
INVX1 gate4168(.O (I16559), .I (g5512));
INVX1 gate4169(.O (g9338), .I (I16559));
INVX1 gate4170(.O (I16562), .I (g6000));
INVX1 gate4171(.O (g9341), .I (I16562));
INVX1 gate4172(.O (g9342), .I (g5972));
INVX1 gate4173(.O (I16566), .I (g5556));
INVX1 gate4174(.O (g9351), .I (I16566));
INVX1 gate4175(.O (I16569), .I (g6000));
INVX1 gate4176(.O (g9354), .I (I16569));
INVX1 gate4177(.O (g9355), .I (g7639));
INVX1 gate4178(.O (g9356), .I (g5665));
INVX1 gate4179(.O (I16578), .I (g6448));
INVX1 gate4180(.O (g9368), .I (I16578));
INVX1 gate4181(.O (I16581), .I (g5438));
INVX1 gate4182(.O (g9371), .I (I16581));
INVX1 gate4183(.O (g9374), .I (g5761));
INVX1 gate4184(.O (I16587), .I (g3462));
INVX1 gate4185(.O (g9384), .I (I16587));
INVX1 gate4186(.O (I16590), .I (g5473));
INVX1 gate4187(.O (g9387), .I (I16590));
INVX1 gate4188(.O (I16593), .I (g6059));
INVX1 gate4189(.O (g9390), .I (I16593));
INVX1 gate4190(.O (g9391), .I (g5867));
INVX1 gate4191(.O (I16598), .I (g3618));
INVX1 gate4192(.O (g9401), .I (I16598));
INVX1 gate4193(.O (I16601), .I (g7015));
INVX1 gate4194(.O (g9404), .I (I16601));
INVX1 gate4195(.O (g9407), .I (g5945));
INVX1 gate4196(.O (I16605), .I (g7265));
INVX1 gate4197(.O (g9416), .I (I16605));
INVX1 gate4198(.O (I16608), .I (g5556));
INVX1 gate4199(.O (g9419), .I (I16608));
INVX1 gate4200(.O (I16611), .I (g6000));
INVX1 gate4201(.O (g9422), .I (I16611));
INVX1 gate4202(.O (g9423), .I (g5428));
INVX1 gate4203(.O (g9424), .I (g5469));
INVX1 gate4204(.O (g9425), .I (g5346));
INVX1 gate4205(.O (g9426), .I (g5543));
INVX1 gate4206(.O (g9427), .I (g5645));
INVX1 gate4207(.O (I16624), .I (g3306));
INVX1 gate4208(.O (g9443), .I (I16624));
INVX1 gate4209(.O (I16627), .I (g6448));
INVX1 gate4210(.O (g9446), .I (I16627));
INVX1 gate4211(.O (I16630), .I (g6057));
INVX1 gate4212(.O (g9449), .I (I16630));
INVX1 gate4213(.O (I16633), .I (g6486));
INVX1 gate4214(.O (g9450), .I (I16633));
INVX1 gate4215(.O (g9453), .I (g5717));
INVX1 gate4216(.O (I16641), .I (g6713));
INVX1 gate4217(.O (g9465), .I (I16641));
INVX1 gate4218(.O (I16644), .I (g5473));
INVX1 gate4219(.O (g9468), .I (I16644));
INVX1 gate4220(.O (g9471), .I (g5820));
INVX1 gate4221(.O (I16650), .I (g3618));
INVX1 gate4222(.O (g9481), .I (I16650));
INVX1 gate4223(.O (I16653), .I (g5512));
INVX1 gate4224(.O (g9484), .I (I16653));
INVX1 gate4225(.O (I16656), .I (g6066));
INVX1 gate4226(.O (g9487), .I (I16656));
INVX1 gate4227(.O (g9488), .I (g5914));
INVX1 gate4228(.O (I16661), .I (g3774));
INVX1 gate4229(.O (g9498), .I (I16661));
INVX1 gate4230(.O (I16664), .I (g7265));
INVX1 gate4231(.O (g9501), .I (I16664));
INVX1 gate4232(.O (g9504), .I (g6149));
INVX1 gate4233(.O (g9505), .I (g6227));
INVX1 gate4234(.O (g9506), .I (g6444));
INVX1 gate4235(.O (g9507), .I (g5953));
INVX1 gate4236(.O (I16677), .I (g3306));
INVX1 gate4237(.O (g9524), .I (I16677));
INVX1 gate4238(.O (g9527), .I (g5508));
INVX1 gate4239(.O (I16681), .I (g6643));
INVX1 gate4240(.O (g9528), .I (I16681));
INVX1 gate4241(.O (I16684), .I (g6486));
INVX1 gate4242(.O (g9531), .I (I16684));
INVX1 gate4243(.O (g9569), .I (g5683));
INVX1 gate4244(.O (I16694), .I (g3462));
INVX1 gate4245(.O (g9585), .I (I16694));
INVX1 gate4246(.O (I16697), .I (g6713));
INVX1 gate4247(.O (g9588), .I (I16697));
INVX1 gate4248(.O (I16700), .I (g6064));
INVX1 gate4249(.O (g9591), .I (I16700));
INVX1 gate4250(.O (I16703), .I (g6751));
INVX1 gate4251(.O (g9592), .I (I16703));
INVX1 gate4252(.O (g9595), .I (g5775));
INVX1 gate4253(.O (I16711), .I (g7015));
INVX1 gate4254(.O (g9607), .I (I16711));
INVX1 gate4255(.O (I16714), .I (g5512));
INVX1 gate4256(.O (g9610), .I (I16714));
INVX1 gate4257(.O (g9613), .I (g5876));
INVX1 gate4258(.O (I16720), .I (g3774));
INVX1 gate4259(.O (g9623), .I (I16720));
INVX1 gate4260(.O (I16723), .I (g5556));
INVX1 gate4261(.O (g9626), .I (I16723));
INVX1 gate4262(.O (I16726), .I (g6085));
INVX1 gate4263(.O (g9629), .I (I16726));
INVX1 gate4264(.O (I16741), .I (g6062));
INVX1 gate4265(.O (g9640), .I (I16741));
INVX1 gate4266(.O (I16744), .I (g3338));
INVX1 gate4267(.O (g9641), .I (I16744));
INVX1 gate4268(.O (I16747), .I (g6643));
INVX1 gate4269(.O (g9644), .I (I16747));
INVX1 gate4270(.O (g9649), .I (g5982));
INVX1 gate4271(.O (I16759), .I (g3462));
INVX1 gate4272(.O (g9666), .I (I16759));
INVX1 gate4273(.O (g9669), .I (g5552));
INVX1 gate4274(.O (I16763), .I (g6945));
INVX1 gate4275(.O (g9670), .I (I16763));
INVX1 gate4276(.O (I16766), .I (g6751));
INVX1 gate4277(.O (g9673), .I (I16766));
INVX1 gate4278(.O (g9711), .I (g5735));
INVX1 gate4279(.O (I16776), .I (g3618));
INVX1 gate4280(.O (g9727), .I (I16776));
INVX1 gate4281(.O (I16779), .I (g7015));
INVX1 gate4282(.O (g9730), .I (I16779));
INVX1 gate4283(.O (I16782), .I (g6083));
INVX1 gate4284(.O (g9733), .I (I16782));
INVX1 gate4285(.O (I16785), .I (g7053));
INVX1 gate4286(.O (g9734), .I (I16785));
INVX1 gate4287(.O (g9737), .I (g5834));
INVX1 gate4288(.O (I16793), .I (g7265));
INVX1 gate4289(.O (g9749), .I (I16793));
INVX1 gate4290(.O (I16796), .I (g5556));
INVX1 gate4291(.O (g9752), .I (I16796));
INVX1 gate4292(.O (g9755), .I (g5431));
INVX1 gate4293(.O (g9756), .I (g5504));
INVX1 gate4294(.O (g9757), .I (g5601));
INVX1 gate4295(.O (g9758), .I (g5618));
INVX1 gate4296(.O (I16811), .I (g3338));
INVX1 gate4297(.O (g9767), .I (I16811));
INVX1 gate4298(.O (I16814), .I (g6486));
INVX1 gate4299(.O (g9770), .I (I16814));
INVX1 gate4300(.O (I16832), .I (g6081));
INVX1 gate4301(.O (g9786), .I (I16832));
INVX1 gate4302(.O (I16835), .I (g3494));
INVX1 gate4303(.O (g9787), .I (I16835));
INVX1 gate4304(.O (I16838), .I (g6945));
INVX1 gate4305(.O (g9790), .I (I16838));
INVX1 gate4306(.O (g9795), .I (g6019));
INVX1 gate4307(.O (I16850), .I (g3618));
INVX1 gate4308(.O (g9812), .I (I16850));
INVX1 gate4309(.O (g9815), .I (g5598));
INVX1 gate4310(.O (I16854), .I (g7195));
INVX1 gate4311(.O (g9816), .I (I16854));
INVX1 gate4312(.O (I16857), .I (g7053));
INVX1 gate4313(.O (g9819), .I (I16857));
INVX1 gate4314(.O (g9857), .I (g5793));
INVX1 gate4315(.O (I16867), .I (g3774));
INVX1 gate4316(.O (g9873), .I (I16867));
INVX1 gate4317(.O (I16870), .I (g7265));
INVX1 gate4318(.O (g9876), .I (I16870));
INVX1 gate4319(.O (I16873), .I (g6102));
INVX1 gate4320(.O (g9879), .I (I16873));
INVX1 gate4321(.O (I16876), .I (g7303));
INVX1 gate4322(.O (g9880), .I (I16876));
INVX1 gate4323(.O (g9884), .I (g6310));
INVX1 gate4324(.O (g9885), .I (g6905));
INVX1 gate4325(.O (g9886), .I (g7149));
INVX1 gate4326(.O (I16897), .I (g6643));
INVX1 gate4327(.O (g9895), .I (I16897));
INVX1 gate4328(.O (I16900), .I (g6486));
INVX1 gate4329(.O (g9898), .I (I16900));
INVX1 gate4330(.O (I16915), .I (g3494));
INVX1 gate4331(.O (g9913), .I (I16915));
INVX1 gate4332(.O (I16918), .I (g6751));
INVX1 gate4333(.O (g9916), .I (I16918));
INVX1 gate4334(.O (I16936), .I (g6100));
INVX1 gate4335(.O (g9932), .I (I16936));
INVX1 gate4336(.O (I16939), .I (g3650));
INVX1 gate4337(.O (g9933), .I (I16939));
INVX1 gate4338(.O (I16942), .I (g7195));
INVX1 gate4339(.O (g9936), .I (I16942));
INVX1 gate4340(.O (g9941), .I (g6035));
INVX1 gate4341(.O (I16954), .I (g3774));
INVX1 gate4342(.O (g9958), .I (I16954));
INVX1 gate4343(.O (g9961), .I (g5615));
INVX1 gate4344(.O (I16958), .I (g7391));
INVX1 gate4345(.O (g9962), .I (I16958));
INVX1 gate4346(.O (I16961), .I (g7303));
INVX1 gate4347(.O (g9965), .I (I16961));
INVX1 gate4348(.O (I16972), .I (g3900));
INVX1 gate4349(.O (g10004), .I (I16972));
INVX1 gate4350(.O (g10015), .I (g5292));
INVX1 gate4351(.O (I16984), .I (g7936));
INVX1 gate4352(.O (g10016), .I (I16984));
INVX1 gate4353(.O (I16987), .I (g6079));
INVX1 gate4354(.O (g10017), .I (I16987));
INVX1 gate4355(.O (I16990), .I (g3338));
INVX1 gate4356(.O (g10018), .I (I16990));
INVX1 gate4357(.O (I16993), .I (g6643));
INVX1 gate4358(.O (g10021), .I (I16993));
INVX1 gate4359(.O (I17009), .I (g6945));
INVX1 gate4360(.O (g10049), .I (I17009));
INVX1 gate4361(.O (I17012), .I (g6751));
INVX1 gate4362(.O (g10052), .I (I17012));
INVX1 gate4363(.O (I17027), .I (g3650));
INVX1 gate4364(.O (g10067), .I (I17027));
INVX1 gate4365(.O (I17030), .I (g7053));
INVX1 gate4366(.O (g10070), .I (I17030));
INVX1 gate4367(.O (I17048), .I (g6117));
INVX1 gate4368(.O (g10086), .I (I17048));
INVX1 gate4369(.O (I17051), .I (g3806));
INVX1 gate4370(.O (g10087), .I (I17051));
INVX1 gate4371(.O (I17054), .I (g7391));
INVX1 gate4372(.O (g10090), .I (I17054));
INVX1 gate4373(.O (I17066), .I (g3900));
INVX1 gate4374(.O (g10096), .I (I17066));
INVX1 gate4375(.O (g10099), .I (g7700));
INVX1 gate4376(.O (I17070), .I (g7528));
INVX1 gate4377(.O (g10100), .I (I17070));
INVX1 gate4378(.O (I17081), .I (g3338));
INVX1 gate4379(.O (g10109), .I (I17081));
INVX1 gate4380(.O (g10124), .I (g5326));
INVX1 gate4381(.O (I17097), .I (g7936));
INVX1 gate4382(.O (g10125), .I (I17097));
INVX1 gate4383(.O (I17100), .I (g6098));
INVX1 gate4384(.O (g10126), .I (I17100));
INVX1 gate4385(.O (I17103), .I (g3494));
INVX1 gate4386(.O (g10127), .I (I17103));
INVX1 gate4387(.O (I17106), .I (g6945));
INVX1 gate4388(.O (g10130), .I (I17106));
INVX1 gate4389(.O (I17122), .I (g7195));
INVX1 gate4390(.O (g10158), .I (I17122));
INVX1 gate4391(.O (I17125), .I (g7053));
INVX1 gate4392(.O (g10161), .I (I17125));
INVX1 gate4393(.O (I17140), .I (g3806));
INVX1 gate4394(.O (g10176), .I (I17140));
INVX1 gate4395(.O (I17143), .I (g7303));
INVX1 gate4396(.O (g10179), .I (I17143));
INVX1 gate4397(.O (I17159), .I (g3900));
INVX1 gate4398(.O (g10189), .I (I17159));
INVX1 gate4399(.O (I17184), .I (g3494));
INVX1 gate4400(.O (g10214), .I (I17184));
INVX1 gate4401(.O (g10229), .I (g5349));
INVX1 gate4402(.O (I17200), .I (g7936));
INVX1 gate4403(.O (g10230), .I (I17200));
INVX1 gate4404(.O (I17203), .I (g6115));
INVX1 gate4405(.O (g10231), .I (I17203));
INVX1 gate4406(.O (I17206), .I (g3650));
INVX1 gate4407(.O (g10232), .I (I17206));
INVX1 gate4408(.O (I17209), .I (g7195));
INVX1 gate4409(.O (g10235), .I (I17209));
INVX1 gate4410(.O (I17225), .I (g7391));
INVX1 gate4411(.O (g10263), .I (I17225));
INVX1 gate4412(.O (I17228), .I (g7303));
INVX1 gate4413(.O (g10266), .I (I17228));
INVX1 gate4414(.O (I17235), .I (g3900));
INVX1 gate4415(.O (g10273), .I (I17235));
INVX1 gate4416(.O (I17238), .I (g3900));
INVX1 gate4417(.O (g10276), .I (I17238));
INVX1 gate4418(.O (I17278), .I (g3650));
INVX1 gate4419(.O (g10316), .I (I17278));
INVX1 gate4420(.O (g10331), .I (g5366));
INVX1 gate4421(.O (I17294), .I (g7936));
INVX1 gate4422(.O (g10332), .I (I17294));
INVX1 gate4423(.O (I17297), .I (g6130));
INVX1 gate4424(.O (g10333), .I (I17297));
INVX1 gate4425(.O (I17300), .I (g3806));
INVX1 gate4426(.O (g10334), .I (I17300));
INVX1 gate4427(.O (I17303), .I (g7391));
INVX1 gate4428(.O (g10337), .I (I17303));
INVX1 gate4429(.O (I17311), .I (g3900));
INVX1 gate4430(.O (g10357), .I (I17311));
INVX1 gate4431(.O (I17363), .I (g3806));
INVX1 gate4432(.O (g10409), .I (I17363));
INVX1 gate4433(.O (I17370), .I (g3900));
INVX1 gate4434(.O (g10416), .I (I17370));
INVX1 gate4435(.O (I17373), .I (g3900));
INVX1 gate4436(.O (g10419), .I (I17373));
INVX1 gate4437(.O (g10424), .I (g7910));
INVX1 gate4438(.O (g10481), .I (g7826));
INVX1 gate4439(.O (I17433), .I (g3900));
INVX1 gate4440(.O (g10482), .I (I17433));
INVX1 gate4441(.O (g10486), .I (g7957));
INVX1 gate4442(.O (g10500), .I (g7962));
INVX1 gate4443(.O (I17483), .I (g3900));
INVX1 gate4444(.O (g10542), .I (I17483));
INVX1 gate4445(.O (I17486), .I (g3900));
INVX1 gate4446(.O (g10545), .I (I17486));
INVX1 gate4447(.O (g10549), .I (g7999));
INVX1 gate4448(.O (g10560), .I (g8008));
INVX1 gate4449(.O (g10574), .I (g8013));
INVX1 gate4450(.O (I17527), .I (g3900));
INVX1 gate4451(.O (g10601), .I (I17527));
INVX1 gate4452(.O (g10606), .I (g8074));
INVX1 gate4453(.O (g10617), .I (g8083));
INVX1 gate4454(.O (g10631), .I (g8088));
INVX1 gate4455(.O (I17557), .I (g3900));
INVX1 gate4456(.O (g10646), .I (I17557));
INVX1 gate4457(.O (g10653), .I (g8159));
INVX1 gate4458(.O (g10664), .I (g8168));
INVX1 gate4459(.O (g10683), .I (g8245));
INVX1 gate4460(.O (g10694), .I (g4326));
INVX1 gate4461(.O (g10714), .I (g4495));
INVX1 gate4462(.O (g10730), .I (g6173));
INVX1 gate4463(.O (g10735), .I (g4671));
INVX1 gate4464(.O (g10749), .I (g6205));
INVX1 gate4465(.O (g10754), .I (g4848));
INVX1 gate4466(.O (g10765), .I (g6048));
INVX1 gate4467(.O (g10766), .I (g6676));
INVX1 gate4468(.O (g10767), .I (g6294));
INVX1 gate4469(.O (g10772), .I (g6978));
INVX1 gate4470(.O (g10773), .I (g6431));
INVX1 gate4471(.O (I17627), .I (g7575));
INVX1 gate4472(.O (g10779), .I (I17627));
INVX1 gate4473(.O (g10783), .I (g7228));
INVX1 gate4474(.O (I17632), .I (g6183));
INVX1 gate4475(.O (g10787), .I (I17632));
INVX1 gate4476(.O (g10788), .I (g7424));
INVX1 gate4477(.O (I17637), .I (g6204));
INVX1 gate4478(.O (g10792), .I (I17637));
INVX1 gate4479(.O (I17641), .I (g6215));
INVX1 gate4480(.O (g10796), .I (I17641));
INVX1 gate4481(.O (I17645), .I (g6288));
INVX1 gate4482(.O (g10800), .I (I17645));
INVX1 gate4483(.O (I17649), .I (g6293));
INVX1 gate4484(.O (g10804), .I (I17649));
INVX1 gate4485(.O (I17653), .I (g6304));
INVX1 gate4486(.O (g10808), .I (I17653));
INVX1 gate4487(.O (g10809), .I (g5701));
INVX1 gate4488(.O (I17658), .I (g6367));
INVX1 gate4489(.O (g10813), .I (I17658));
INVX1 gate4490(.O (I17662), .I (g6425));
INVX1 gate4491(.O (g10817), .I (I17662));
INVX1 gate4492(.O (I17666), .I (g6430));
INVX1 gate4493(.O (g10821), .I (I17666));
INVX1 gate4494(.O (I17670), .I (g6441));
INVX1 gate4495(.O (g10825), .I (I17670));
INVX1 gate4496(.O (I17673), .I (g8107));
INVX1 gate4497(.O (g10826), .I (I17673));
INVX1 gate4498(.O (g10829), .I (g5749));
INVX1 gate4499(.O (I17677), .I (g6517));
INVX1 gate4500(.O (g10830), .I (I17677));
INVX1 gate4501(.O (I17681), .I (g6572));
INVX1 gate4502(.O (g10834), .I (I17681));
INVX1 gate4503(.O (I17685), .I (g6630));
INVX1 gate4504(.O (g10838), .I (I17685));
INVX1 gate4505(.O (I17689), .I (g6635));
INVX1 gate4506(.O (g10842), .I (I17689));
INVX1 gate4507(.O (I17692), .I (g8107));
INVX1 gate4508(.O (g10843), .I (I17692));
INVX1 gate4509(.O (g10846), .I (g5799));
INVX1 gate4510(.O (g10847), .I (g5800));
INVX1 gate4511(.O (g10848), .I (g5801));
INVX1 gate4512(.O (I17698), .I (g6711));
INVX1 gate4513(.O (g10849), .I (I17698));
INVX1 gate4514(.O (I17701), .I (g6781));
INVX1 gate4515(.O (g10850), .I (I17701));
INVX1 gate4516(.O (I17705), .I (g6836));
INVX1 gate4517(.O (g10854), .I (I17705));
INVX1 gate4518(.O (I17709), .I (g6894));
INVX1 gate4519(.O (g10858), .I (I17709));
INVX1 gate4520(.O (I17712), .I (g8031));
INVX1 gate4521(.O (g10859), .I (I17712));
INVX1 gate4522(.O (I17715), .I (g8107));
INVX1 gate4523(.O (g10862), .I (I17715));
INVX1 gate4524(.O (g10865), .I (g6131));
INVX1 gate4525(.O (g10866), .I (g5849));
INVX1 gate4526(.O (g10867), .I (g5850));
INVX1 gate4527(.O (I17721), .I (g6641));
INVX1 gate4528(.O (g10868), .I (I17721));
INVX1 gate4529(.O (I17724), .I (g6942));
INVX1 gate4530(.O (g10869), .I (I17724));
INVX1 gate4531(.O (I17727), .I (g7013));
INVX1 gate4532(.O (g10870), .I (I17727));
INVX1 gate4533(.O (I17730), .I (g7083));
INVX1 gate4534(.O (g10871), .I (I17730));
INVX1 gate4535(.O (I17734), .I (g7138));
INVX1 gate4536(.O (g10875), .I (I17734));
INVX1 gate4537(.O (I17737), .I (g6000));
INVX1 gate4538(.O (g10876), .I (I17737));
INVX1 gate4539(.O (I17740), .I (g8031));
INVX1 gate4540(.O (g10877), .I (I17740));
INVX1 gate4541(.O (I17743), .I (g8107));
INVX1 gate4542(.O (g10880), .I (I17743));
INVX1 gate4543(.O (I17746), .I (g8107));
INVX1 gate4544(.O (g10883), .I (I17746));
INVX1 gate4545(.O (g10886), .I (g5889));
INVX1 gate4546(.O (I17750), .I (g7157));
INVX1 gate4547(.O (g10887), .I (I17750));
INVX1 gate4548(.O (I17753), .I (g6943));
INVX1 gate4549(.O (g10888), .I (I17753));
INVX1 gate4550(.O (I17756), .I (g7192));
INVX1 gate4551(.O (g10889), .I (I17756));
INVX1 gate4552(.O (I17759), .I (g7263));
INVX1 gate4553(.O (g10890), .I (I17759));
INVX1 gate4554(.O (I17762), .I (g7333));
INVX1 gate4555(.O (g10891), .I (I17762));
INVX1 gate4556(.O (I17765), .I (g7976));
INVX1 gate4557(.O (g10892), .I (I17765));
INVX1 gate4558(.O (I17768), .I (g8031));
INVX1 gate4559(.O (g10895), .I (I17768));
INVX1 gate4560(.O (I17771), .I (g8107));
INVX1 gate4561(.O (g10898), .I (I17771));
INVX1 gate4562(.O (I17774), .I (g8107));
INVX1 gate4563(.O (g10901), .I (I17774));
INVX1 gate4564(.O (g10904), .I (g5922));
INVX1 gate4565(.O (g10905), .I (g5923));
INVX1 gate4566(.O (g10906), .I (g5924));
INVX1 gate4567(.O (I17780), .I (g7348));
INVX1 gate4568(.O (g10907), .I (I17780));
INVX1 gate4569(.O (I17783), .I (g7353));
INVX1 gate4570(.O (g10908), .I (I17783));
INVX1 gate4571(.O (I17786), .I (g7193));
INVX1 gate4572(.O (g10909), .I (I17786));
INVX1 gate4573(.O (I17789), .I (g7388));
INVX1 gate4574(.O (g10910), .I (I17789));
INVX1 gate4575(.O (I17792), .I (g7459));
INVX1 gate4576(.O (g10911), .I (I17792));
INVX1 gate4577(.O (I17795), .I (g7976));
INVX1 gate4578(.O (g10912), .I (I17795));
INVX1 gate4579(.O (I17798), .I (g8031));
INVX1 gate4580(.O (g10915), .I (I17798));
INVX1 gate4581(.O (I17801), .I (g8107));
INVX1 gate4582(.O (g10918), .I (I17801));
INVX1 gate4583(.O (I17804), .I (g8031));
INVX1 gate4584(.O (g10921), .I (I17804));
INVX1 gate4585(.O (I17807), .I (g8107));
INVX1 gate4586(.O (g10924), .I (I17807));
INVX1 gate4587(.O (g10927), .I (g6153));
INVX1 gate4588(.O (g10928), .I (g5951));
INVX1 gate4589(.O (g10929), .I (g5952));
INVX1 gate4590(.O (I17813), .I (g5707));
INVX1 gate4591(.O (g10930), .I (I17813));
INVX1 gate4592(.O (I17816), .I (g7346));
INVX1 gate4593(.O (g10931), .I (I17816));
INVX1 gate4594(.O (I17819), .I (g6448));
INVX1 gate4595(.O (g10932), .I (I17819));
INVX1 gate4596(.O (I17822), .I (g7478));
INVX1 gate4597(.O (g10933), .I (I17822));
INVX1 gate4598(.O (I17825), .I (g7483));
INVX1 gate4599(.O (g10934), .I (I17825));
INVX1 gate4600(.O (I17828), .I (g7389));
INVX1 gate4601(.O (g10935), .I (I17828));
INVX1 gate4602(.O (I17831), .I (g7518));
INVX1 gate4603(.O (g10936), .I (I17831));
INVX1 gate4604(.O (I17834), .I (g7976));
INVX1 gate4605(.O (g10937), .I (I17834));
INVX1 gate4606(.O (I17837), .I (g8031));
INVX1 gate4607(.O (g10940), .I (I17837));
INVX1 gate4608(.O (I17840), .I (g8107));
INVX1 gate4609(.O (g10943), .I (I17840));
INVX1 gate4610(.O (I17843), .I (g8031));
INVX1 gate4611(.O (g10946), .I (I17843));
INVX1 gate4612(.O (I17846), .I (g8107));
INVX1 gate4613(.O (g10949), .I (I17846));
INVX1 gate4614(.O (I17849), .I (g8103));
INVX1 gate4615(.O (g10952), .I (I17849));
INVX1 gate4616(.O (g10961), .I (g5978));
INVX1 gate4617(.O (g10962), .I (g5979));
INVX1 gate4618(.O (I17854), .I (g6232));
INVX1 gate4619(.O (g10963), .I (I17854));
INVX1 gate4620(.O (I17857), .I (g6448));
INVX1 gate4621(.O (g10966), .I (I17857));
INVX1 gate4622(.O (I17860), .I (g5765));
INVX1 gate4623(.O (g10967), .I (I17860));
INVX1 gate4624(.O (I17863), .I (g7476));
INVX1 gate4625(.O (g10968), .I (I17863));
INVX1 gate4626(.O (I17866), .I (g6713));
INVX1 gate4627(.O (g10969), .I (I17866));
INVX1 gate4628(.O (I17869), .I (g7534));
INVX1 gate4629(.O (g10972), .I (I17869));
INVX1 gate4630(.O (I17872), .I (g7539));
INVX1 gate4631(.O (g10973), .I (I17872));
INVX1 gate4632(.O (I17875), .I (g7976));
INVX1 gate4633(.O (g10974), .I (I17875));
INVX1 gate4634(.O (I17878), .I (g8031));
INVX1 gate4635(.O (g10977), .I (I17878));
INVX1 gate4636(.O (I17881), .I (g7976));
INVX1 gate4637(.O (g10980), .I (I17881));
INVX1 gate4638(.O (I17884), .I (g8031));
INVX1 gate4639(.O (g10983), .I (I17884));
INVX1 gate4640(.O (g10986), .I (g6014));
INVX1 gate4641(.O (g10987), .I (g6015));
INVX1 gate4642(.O (I17889), .I (g6314));
INVX1 gate4643(.O (g10988), .I (I17889));
INVX1 gate4644(.O (I17892), .I (g6232));
INVX1 gate4645(.O (g10991), .I (I17892));
INVX1 gate4646(.O (I17895), .I (g6448));
INVX1 gate4647(.O (g10994), .I (I17895));
INVX1 gate4648(.O (I17898), .I (g6643));
INVX1 gate4649(.O (g10995), .I (I17898));
INVX1 gate4650(.O (I17901), .I (g6369));
INVX1 gate4651(.O (g10996), .I (I17901));
INVX1 gate4652(.O (I17904), .I (g6713));
INVX1 gate4653(.O (g10999), .I (I17904));
INVX1 gate4654(.O (I17907), .I (g5824));
INVX1 gate4655(.O (g11002), .I (I17907));
INVX1 gate4656(.O (I17910), .I (g7532));
INVX1 gate4657(.O (g11003), .I (I17910));
INVX1 gate4658(.O (I17913), .I (g7015));
INVX1 gate4659(.O (g11004), .I (I17913));
INVX1 gate4660(.O (I17916), .I (g7560));
INVX1 gate4661(.O (g11007), .I (I17916));
INVX1 gate4662(.O (I17919), .I (g7976));
INVX1 gate4663(.O (g11008), .I (I17919));
INVX1 gate4664(.O (I17922), .I (g8031));
INVX1 gate4665(.O (g11011), .I (I17922));
INVX1 gate4666(.O (I17925), .I (g7976));
INVX1 gate4667(.O (g11014), .I (I17925));
INVX1 gate4668(.O (I17928), .I (g8031));
INVX1 gate4669(.O (g11017), .I (I17928));
INVX1 gate4670(.O (g11020), .I (g6029));
INVX1 gate4671(.O (g11021), .I (g6030));
INVX1 gate4672(.O (I17933), .I (g3254));
INVX1 gate4673(.O (g11022), .I (I17933));
INVX1 gate4674(.O (I17936), .I (g6314));
INVX1 gate4675(.O (g11025), .I (I17936));
INVX1 gate4676(.O (I17939), .I (g6232));
INVX1 gate4677(.O (g11028), .I (I17939));
INVX1 gate4678(.O (I17942), .I (g5548));
INVX1 gate4679(.O (g11031), .I (I17942));
INVX1 gate4680(.O (I17945), .I (g5668));
INVX1 gate4681(.O (g11032), .I (I17945));
INVX1 gate4682(.O (I17948), .I (g6643));
INVX1 gate4683(.O (g11035), .I (I17948));
INVX1 gate4684(.O (I17951), .I (g6519));
INVX1 gate4685(.O (g11036), .I (I17951));
INVX1 gate4686(.O (I17954), .I (g6369));
INVX1 gate4687(.O (g11039), .I (I17954));
INVX1 gate4688(.O (I17957), .I (g6713));
INVX1 gate4689(.O (g11042), .I (I17957));
INVX1 gate4690(.O (I17960), .I (g6945));
INVX1 gate4691(.O (g11045), .I (I17960));
INVX1 gate4692(.O (I17963), .I (g6574));
INVX1 gate4693(.O (g11048), .I (I17963));
INVX1 gate4694(.O (I17966), .I (g7015));
INVX1 gate4695(.O (g11051), .I (I17966));
INVX1 gate4696(.O (I17969), .I (g5880));
INVX1 gate4697(.O (g11054), .I (I17969));
INVX1 gate4698(.O (I17972), .I (g7558));
INVX1 gate4699(.O (g11055), .I (I17972));
INVX1 gate4700(.O (I17975), .I (g7265));
INVX1 gate4701(.O (g11056), .I (I17975));
INVX1 gate4702(.O (I17978), .I (g7795));
INVX1 gate4703(.O (g11059), .I (I17978));
INVX1 gate4704(.O (I17981), .I (g7976));
INVX1 gate4705(.O (g11063), .I (I17981));
INVX1 gate4706(.O (I17984), .I (g7976));
INVX1 gate4707(.O (g11066), .I (I17984));
INVX1 gate4708(.O (g11069), .I (g8257));
INVX1 gate4709(.O (g11078), .I (g6041));
INVX1 gate4710(.O (I17989), .I (g3254));
INVX1 gate4711(.O (g11079), .I (I17989));
INVX1 gate4712(.O (I17992), .I (g6314));
INVX1 gate4713(.O (g11082), .I (I17992));
INVX1 gate4714(.O (I17995), .I (g6232));
INVX1 gate4715(.O (g11085), .I (I17995));
INVX1 gate4716(.O (I17998), .I (g5668));
INVX1 gate4717(.O (g11088), .I (I17998));
INVX1 gate4718(.O (I18001), .I (g6643));
INVX1 gate4719(.O (g11091), .I (I18001));
INVX1 gate4720(.O (I18004), .I (g3410));
INVX1 gate4721(.O (g11092), .I (I18004));
INVX1 gate4722(.O (I18007), .I (g6519));
INVX1 gate4723(.O (g11095), .I (I18007));
INVX1 gate4724(.O (I18010), .I (g6369));
INVX1 gate4725(.O (g11098), .I (I18010));
INVX1 gate4726(.O (I18013), .I (g5594));
INVX1 gate4727(.O (g11101), .I (I18013));
INVX1 gate4728(.O (I18016), .I (g5720));
INVX1 gate4729(.O (g11102), .I (I18016));
INVX1 gate4730(.O (I18019), .I (g6945));
INVX1 gate4731(.O (g11105), .I (I18019));
INVX1 gate4732(.O (I18022), .I (g6783));
INVX1 gate4733(.O (g11108), .I (I18022));
INVX1 gate4734(.O (I18025), .I (g6574));
INVX1 gate4735(.O (g11111), .I (I18025));
INVX1 gate4736(.O (I18028), .I (g7015));
INVX1 gate4737(.O (g11114), .I (I18028));
INVX1 gate4738(.O (I18031), .I (g7195));
INVX1 gate4739(.O (g11117), .I (I18031));
INVX1 gate4740(.O (I18034), .I (g6838));
INVX1 gate4741(.O (g11120), .I (I18034));
INVX1 gate4742(.O (I18037), .I (g7265));
INVX1 gate4743(.O (g11123), .I (I18037));
INVX1 gate4744(.O (I18040), .I (g7976));
INVX1 gate4745(.O (g11126), .I (I18040));
INVX1 gate4746(.O (I18043), .I (g7976));
INVX1 gate4747(.O (g11129), .I (I18043));
INVX1 gate4748(.O (I18046), .I (g3254));
INVX1 gate4749(.O (g11132), .I (I18046));
INVX1 gate4750(.O (I18049), .I (g6314));
INVX1 gate4751(.O (g11135), .I (I18049));
INVX1 gate4752(.O (I18052), .I (g6232));
INVX1 gate4753(.O (g11138), .I (I18052));
INVX1 gate4754(.O (I18055), .I (g5668));
INVX1 gate4755(.O (g11141), .I (I18055));
INVX1 gate4756(.O (I18058), .I (g6643));
INVX1 gate4757(.O (g11144), .I (I18058));
INVX1 gate4758(.O (I18061), .I (g3410));
INVX1 gate4759(.O (g11145), .I (I18061));
INVX1 gate4760(.O (I18064), .I (g6519));
INVX1 gate4761(.O (g11148), .I (I18064));
INVX1 gate4762(.O (I18067), .I (g6369));
INVX1 gate4763(.O (g11151), .I (I18067));
INVX1 gate4764(.O (I18070), .I (g5720));
INVX1 gate4765(.O (g11154), .I (I18070));
INVX1 gate4766(.O (I18073), .I (g6945));
INVX1 gate4767(.O (g11157), .I (I18073));
INVX1 gate4768(.O (I18076), .I (g3566));
INVX1 gate4769(.O (g11160), .I (I18076));
INVX1 gate4770(.O (I18079), .I (g6783));
INVX1 gate4771(.O (g11163), .I (I18079));
INVX1 gate4772(.O (I18082), .I (g6574));
INVX1 gate4773(.O (g11166), .I (I18082));
INVX1 gate4774(.O (I18085), .I (g5611));
INVX1 gate4775(.O (g11169), .I (I18085));
INVX1 gate4776(.O (I18088), .I (g5778));
INVX1 gate4777(.O (g11170), .I (I18088));
INVX1 gate4778(.O (I18091), .I (g7195));
INVX1 gate4779(.O (g11173), .I (I18091));
INVX1 gate4780(.O (I18094), .I (g7085));
INVX1 gate4781(.O (g11176), .I (I18094));
INVX1 gate4782(.O (I18097), .I (g6838));
INVX1 gate4783(.O (g11179), .I (I18097));
INVX1 gate4784(.O (I18100), .I (g7265));
INVX1 gate4785(.O (g11182), .I (I18100));
INVX1 gate4786(.O (I18103), .I (g7391));
INVX1 gate4787(.O (g11185), .I (I18103));
INVX1 gate4788(.O (g11190), .I (g3999));
INVX1 gate4789(.O (I18121), .I (g3254));
INVX1 gate4790(.O (g11199), .I (I18121));
INVX1 gate4791(.O (I18124), .I (g6314));
INVX1 gate4792(.O (g11202), .I (I18124));
INVX1 gate4793(.O (I18127), .I (g6232));
INVX1 gate4794(.O (g11205), .I (I18127));
INVX1 gate4795(.O (I18130), .I (g5547));
INVX1 gate4796(.O (g11208), .I (I18130));
INVX1 gate4797(.O (I18133), .I (g6448));
INVX1 gate4798(.O (g11209), .I (I18133));
INVX1 gate4799(.O (I18136), .I (g5668));
INVX1 gate4800(.O (g11210), .I (I18136));
INVX1 gate4801(.O (I18139), .I (g6643));
INVX1 gate4802(.O (g11213), .I (I18139));
INVX1 gate4803(.O (I18142), .I (g3410));
INVX1 gate4804(.O (g11216), .I (I18142));
INVX1 gate4805(.O (I18145), .I (g6519));
INVX1 gate4806(.O (g11219), .I (I18145));
INVX1 gate4807(.O (I18148), .I (g6369));
INVX1 gate4808(.O (g11222), .I (I18148));
INVX1 gate4809(.O (I18151), .I (g5720));
INVX1 gate4810(.O (g11225), .I (I18151));
INVX1 gate4811(.O (I18154), .I (g6945));
INVX1 gate4812(.O (g11228), .I (I18154));
INVX1 gate4813(.O (I18157), .I (g3566));
INVX1 gate4814(.O (g11231), .I (I18157));
INVX1 gate4815(.O (I18160), .I (g6783));
INVX1 gate4816(.O (g11234), .I (I18160));
INVX1 gate4817(.O (I18163), .I (g6574));
INVX1 gate4818(.O (g11237), .I (I18163));
INVX1 gate4819(.O (I18166), .I (g5778));
INVX1 gate4820(.O (g11240), .I (I18166));
INVX1 gate4821(.O (I18169), .I (g7195));
INVX1 gate4822(.O (g11243), .I (I18169));
INVX1 gate4823(.O (I18172), .I (g3722));
INVX1 gate4824(.O (g11246), .I (I18172));
INVX1 gate4825(.O (I18175), .I (g7085));
INVX1 gate4826(.O (g11249), .I (I18175));
INVX1 gate4827(.O (I18178), .I (g6838));
INVX1 gate4828(.O (g11252), .I (I18178));
INVX1 gate4829(.O (I18181), .I (g5636));
INVX1 gate4830(.O (g11255), .I (I18181));
INVX1 gate4831(.O (I18184), .I (g5837));
INVX1 gate4832(.O (g11256), .I (I18184));
INVX1 gate4833(.O (I18187), .I (g7391));
INVX1 gate4834(.O (g11259), .I (I18187));
INVX1 gate4835(.O (I18211), .I (g6232));
INVX1 gate4836(.O (g11265), .I (I18211));
INVX1 gate4837(.O (I18214), .I (g3254));
INVX1 gate4838(.O (g11268), .I (I18214));
INVX1 gate4839(.O (I18217), .I (g6314));
INVX1 gate4840(.O (g11271), .I (I18217));
INVX1 gate4841(.O (I18220), .I (g6232));
INVX1 gate4842(.O (g11274), .I (I18220));
INVX1 gate4843(.O (I18223), .I (g6448));
INVX1 gate4844(.O (g11277), .I (I18223));
INVX1 gate4845(.O (I18226), .I (g5668));
INVX1 gate4846(.O (g11278), .I (I18226));
INVX1 gate4847(.O (I18229), .I (g3410));
INVX1 gate4848(.O (g11281), .I (I18229));
INVX1 gate4849(.O (I18232), .I (g6519));
INVX1 gate4850(.O (g11284), .I (I18232));
INVX1 gate4851(.O (I18235), .I (g6369));
INVX1 gate4852(.O (g11287), .I (I18235));
INVX1 gate4853(.O (I18238), .I (g5593));
INVX1 gate4854(.O (g11290), .I (I18238));
INVX1 gate4855(.O (I18241), .I (g6713));
INVX1 gate4856(.O (g11291), .I (I18241));
INVX1 gate4857(.O (I18244), .I (g5720));
INVX1 gate4858(.O (g11294), .I (I18244));
INVX1 gate4859(.O (I18247), .I (g6945));
INVX1 gate4860(.O (g11297), .I (I18247));
INVX1 gate4861(.O (I18250), .I (g3566));
INVX1 gate4862(.O (g11300), .I (I18250));
INVX1 gate4863(.O (I18253), .I (g6783));
INVX1 gate4864(.O (g11303), .I (I18253));
INVX1 gate4865(.O (I18256), .I (g6574));
INVX1 gate4866(.O (g11306), .I (I18256));
INVX1 gate4867(.O (I18259), .I (g5778));
INVX1 gate4868(.O (g11309), .I (I18259));
INVX1 gate4869(.O (I18262), .I (g7195));
INVX1 gate4870(.O (g11312), .I (I18262));
INVX1 gate4871(.O (I18265), .I (g3722));
INVX1 gate4872(.O (g11315), .I (I18265));
INVX1 gate4873(.O (I18268), .I (g7085));
INVX1 gate4874(.O (g11318), .I (I18268));
INVX1 gate4875(.O (I18271), .I (g6838));
INVX1 gate4876(.O (g11321), .I (I18271));
INVX1 gate4877(.O (I18274), .I (g5837));
INVX1 gate4878(.O (g11324), .I (I18274));
INVX1 gate4879(.O (I18277), .I (g7391));
INVX1 gate4880(.O (g11327), .I (I18277));
INVX1 gate4881(.O (g11332), .I (g4094));
INVX1 gate4882(.O (I18295), .I (g6314));
INVX1 gate4883(.O (g11341), .I (I18295));
INVX1 gate4884(.O (I18298), .I (g6232));
INVX1 gate4885(.O (g11344), .I (I18298));
INVX1 gate4886(.O (I18302), .I (g3254));
INVX1 gate4887(.O (g11348), .I (I18302));
INVX1 gate4888(.O (I18305), .I (g6314));
INVX1 gate4889(.O (g11351), .I (I18305));
INVX1 gate4890(.O (I18308), .I (g6448));
INVX1 gate4891(.O (g11354), .I (I18308));
INVX1 gate4892(.O (I18311), .I (g5668));
INVX1 gate4893(.O (g11355), .I (I18311));
INVX1 gate4894(.O (I18314), .I (g6369));
INVX1 gate4895(.O (g11358), .I (I18314));
INVX1 gate4896(.O (I18317), .I (g3410));
INVX1 gate4897(.O (g11361), .I (I18317));
INVX1 gate4898(.O (I18320), .I (g6519));
INVX1 gate4899(.O (g11364), .I (I18320));
INVX1 gate4900(.O (I18323), .I (g6369));
INVX1 gate4901(.O (g11367), .I (I18323));
INVX1 gate4902(.O (I18326), .I (g6713));
INVX1 gate4903(.O (g11370), .I (I18326));
INVX1 gate4904(.O (I18329), .I (g5720));
INVX1 gate4905(.O (g11373), .I (I18329));
INVX1 gate4906(.O (I18332), .I (g3566));
INVX1 gate4907(.O (g11376), .I (I18332));
INVX1 gate4908(.O (I18335), .I (g6783));
INVX1 gate4909(.O (g11379), .I (I18335));
INVX1 gate4910(.O (I18338), .I (g6574));
INVX1 gate4911(.O (g11382), .I (I18338));
INVX1 gate4912(.O (I18341), .I (g5610));
INVX1 gate4913(.O (g11385), .I (I18341));
INVX1 gate4914(.O (I18344), .I (g7015));
INVX1 gate4915(.O (g11386), .I (I18344));
INVX1 gate4916(.O (I18347), .I (g5778));
INVX1 gate4917(.O (g11389), .I (I18347));
INVX1 gate4918(.O (I18350), .I (g7195));
INVX1 gate4919(.O (g11392), .I (I18350));
INVX1 gate4920(.O (I18353), .I (g3722));
INVX1 gate4921(.O (g11395), .I (I18353));
INVX1 gate4922(.O (I18356), .I (g7085));
INVX1 gate4923(.O (g11398), .I (I18356));
INVX1 gate4924(.O (I18359), .I (g6838));
INVX1 gate4925(.O (g11401), .I (I18359));
INVX1 gate4926(.O (I18362), .I (g5837));
INVX1 gate4927(.O (g11404), .I (I18362));
INVX1 gate4928(.O (I18365), .I (g7391));
INVX1 gate4929(.O (g11407), .I (I18365));
INVX1 gate4930(.O (I18375), .I (g3254));
INVX1 gate4931(.O (g11411), .I (I18375));
INVX1 gate4932(.O (I18378), .I (g6314));
INVX1 gate4933(.O (g11414), .I (I18378));
INVX1 gate4934(.O (I18381), .I (g6232));
INVX1 gate4935(.O (g11417), .I (I18381));
INVX1 gate4936(.O (I18386), .I (g3254));
INVX1 gate4937(.O (g11422), .I (I18386));
INVX1 gate4938(.O (I18389), .I (g6519));
INVX1 gate4939(.O (g11425), .I (I18389));
INVX1 gate4940(.O (I18392), .I (g6369));
INVX1 gate4941(.O (g11428), .I (I18392));
INVX1 gate4942(.O (I18396), .I (g3410));
INVX1 gate4943(.O (g11432), .I (I18396));
INVX1 gate4944(.O (I18399), .I (g6519));
INVX1 gate4945(.O (g11435), .I (I18399));
INVX1 gate4946(.O (I18402), .I (g6713));
INVX1 gate4947(.O (g11438), .I (I18402));
INVX1 gate4948(.O (I18405), .I (g5720));
INVX1 gate4949(.O (g11441), .I (I18405));
INVX1 gate4950(.O (I18408), .I (g6574));
INVX1 gate4951(.O (g11444), .I (I18408));
INVX1 gate4952(.O (I18411), .I (g3566));
INVX1 gate4953(.O (g11447), .I (I18411));
INVX1 gate4954(.O (I18414), .I (g6783));
INVX1 gate4955(.O (g11450), .I (I18414));
INVX1 gate4956(.O (I18417), .I (g6574));
INVX1 gate4957(.O (g11453), .I (I18417));
INVX1 gate4958(.O (I18420), .I (g7015));
INVX1 gate4959(.O (g11456), .I (I18420));
INVX1 gate4960(.O (I18423), .I (g5778));
INVX1 gate4961(.O (g11459), .I (I18423));
INVX1 gate4962(.O (I18426), .I (g3722));
INVX1 gate4963(.O (g11462), .I (I18426));
INVX1 gate4964(.O (I18429), .I (g7085));
INVX1 gate4965(.O (g11465), .I (I18429));
INVX1 gate4966(.O (I18432), .I (g6838));
INVX1 gate4967(.O (g11468), .I (I18432));
INVX1 gate4968(.O (I18435), .I (g5635));
INVX1 gate4969(.O (g11471), .I (I18435));
INVX1 gate4970(.O (I18438), .I (g7265));
INVX1 gate4971(.O (g11472), .I (I18438));
INVX1 gate4972(.O (I18441), .I (g5837));
INVX1 gate4973(.O (g11475), .I (I18441));
INVX1 gate4974(.O (I18444), .I (g7391));
INVX1 gate4975(.O (g11478), .I (I18444));
INVX1 gate4976(.O (g11481), .I (g4204));
INVX1 gate4977(.O (g11490), .I (g8276));
INVX1 gate4978(.O (I18449), .I (g10868));
INVX1 gate4979(.O (g11491), .I (I18449));
INVX1 gate4980(.O (I18452), .I (g10930));
INVX1 gate4981(.O (g11492), .I (I18452));
INVX1 gate4982(.O (I18455), .I (g11031));
INVX1 gate4983(.O (g11493), .I (I18455));
INVX1 gate4984(.O (I18458), .I (g11208));
INVX1 gate4985(.O (g11494), .I (I18458));
INVX1 gate4986(.O (I18461), .I (g10931));
INVX1 gate4987(.O (g11495), .I (I18461));
INVX1 gate4988(.O (I18464), .I (g8620));
INVX1 gate4989(.O (g11496), .I (I18464));
INVX1 gate4990(.O (I18467), .I (g8769));
INVX1 gate4991(.O (g11497), .I (I18467));
INVX1 gate4992(.O (I18470), .I (g8808));
INVX1 gate4993(.O (g11498), .I (I18470));
INVX1 gate4994(.O (I18473), .I (g8839));
INVX1 gate4995(.O (g11499), .I (I18473));
INVX1 gate4996(.O (I18476), .I (g8791));
INVX1 gate4997(.O (g11500), .I (I18476));
INVX1 gate4998(.O (I18479), .I (g8820));
INVX1 gate4999(.O (g11501), .I (I18479));
INVX1 gate5000(.O (I18482), .I (g8859));
INVX1 gate5001(.O (g11502), .I (I18482));
INVX1 gate5002(.O (I18485), .I (g8809));
INVX1 gate5003(.O (g11503), .I (I18485));
INVX1 gate5004(.O (I18488), .I (g8840));
INVX1 gate5005(.O (g11504), .I (I18488));
INVX1 gate5006(.O (I18491), .I (g8891));
INVX1 gate5007(.O (g11505), .I (I18491));
INVX1 gate5008(.O (I18494), .I (g8821));
INVX1 gate5009(.O (g11506), .I (I18494));
INVX1 gate5010(.O (I18497), .I (g8860));
INVX1 gate5011(.O (g11507), .I (I18497));
INVX1 gate5012(.O (I18500), .I (g8924));
INVX1 gate5013(.O (g11508), .I (I18500));
INVX1 gate5014(.O (I18503), .I (g8658));
INVX1 gate5015(.O (g11509), .I (I18503));
INVX1 gate5016(.O (I18506), .I (g8699));
INVX1 gate5017(.O (g11510), .I (I18506));
INVX1 gate5018(.O (I18509), .I (g8770));
INVX1 gate5019(.O (g11511), .I (I18509));
INVX1 gate5020(.O (I18512), .I (g9309));
INVX1 gate5021(.O (g11512), .I (I18512));
INVX1 gate5022(.O (I18515), .I (g8843));
INVX1 gate5023(.O (g11513), .I (I18515));
INVX1 gate5024(.O (I18518), .I (g8893));
INVX1 gate5025(.O (g11514), .I (I18518));
INVX1 gate5026(.O (I18521), .I (g9449));
INVX1 gate5027(.O (g11515), .I (I18521));
INVX1 gate5028(.O (I18524), .I (g9640));
INVX1 gate5029(.O (g11516), .I (I18524));
INVX1 gate5030(.O (I18527), .I (g10017));
INVX1 gate5031(.O (g11517), .I (I18527));
INVX1 gate5032(.O (I18530), .I (g10888));
INVX1 gate5033(.O (g11518), .I (I18530));
INVX1 gate5034(.O (I18533), .I (g10967));
INVX1 gate5035(.O (g11519), .I (I18533));
INVX1 gate5036(.O (I18536), .I (g11101));
INVX1 gate5037(.O (g11520), .I (I18536));
INVX1 gate5038(.O (I18539), .I (g11290));
INVX1 gate5039(.O (g11521), .I (I18539));
INVX1 gate5040(.O (I18542), .I (g10968));
INVX1 gate5041(.O (g11522), .I (I18542));
INVX1 gate5042(.O (I18545), .I (g8630));
INVX1 gate5043(.O (g11523), .I (I18545));
INVX1 gate5044(.O (I18548), .I (g8792));
INVX1 gate5045(.O (g11524), .I (I18548));
INVX1 gate5046(.O (I18551), .I (g8824));
INVX1 gate5047(.O (g11525), .I (I18551));
INVX1 gate5048(.O (I18554), .I (g8866));
INVX1 gate5049(.O (g11526), .I (I18554));
INVX1 gate5050(.O (I18557), .I (g8810));
INVX1 gate5051(.O (g11527), .I (I18557));
INVX1 gate5052(.O (I18560), .I (g8844));
INVX1 gate5053(.O (g11528), .I (I18560));
INVX1 gate5054(.O (I18563), .I (g8897));
INVX1 gate5055(.O (g11529), .I (I18563));
INVX1 gate5056(.O (I18566), .I (g8825));
INVX1 gate5057(.O (g11530), .I (I18566));
INVX1 gate5058(.O (I18569), .I (g8867));
INVX1 gate5059(.O (g11531), .I (I18569));
INVX1 gate5060(.O (I18572), .I (g8931));
INVX1 gate5061(.O (g11532), .I (I18572));
INVX1 gate5062(.O (I18575), .I (g8845));
INVX1 gate5063(.O (g11533), .I (I18575));
INVX1 gate5064(.O (I18578), .I (g8898));
INVX1 gate5065(.O (g11534), .I (I18578));
INVX1 gate5066(.O (I18581), .I (g8964));
INVX1 gate5067(.O (g11535), .I (I18581));
INVX1 gate5068(.O (I18584), .I (g8677));
INVX1 gate5069(.O (g11536), .I (I18584));
INVX1 gate5070(.O (I18587), .I (g8718));
INVX1 gate5071(.O (g11537), .I (I18587));
INVX1 gate5072(.O (I18590), .I (g8793));
INVX1 gate5073(.O (g11538), .I (I18590));
INVX1 gate5074(.O (I18593), .I (g9390));
INVX1 gate5075(.O (g11539), .I (I18593));
INVX1 gate5076(.O (I18596), .I (g8870));
INVX1 gate5077(.O (g11540), .I (I18596));
INVX1 gate5078(.O (I18599), .I (g8933));
INVX1 gate5079(.O (g11541), .I (I18599));
INVX1 gate5080(.O (I18602), .I (g9591));
INVX1 gate5081(.O (g11542), .I (I18602));
INVX1 gate5082(.O (I18605), .I (g9786));
INVX1 gate5083(.O (g11543), .I (I18605));
INVX1 gate5084(.O (I18608), .I (g10126));
INVX1 gate5085(.O (g11544), .I (I18608));
INVX1 gate5086(.O (I18611), .I (g10909));
INVX1 gate5087(.O (g11545), .I (I18611));
INVX1 gate5088(.O (I18614), .I (g11002));
INVX1 gate5089(.O (g11546), .I (I18614));
INVX1 gate5090(.O (I18617), .I (g11169));
INVX1 gate5091(.O (g11547), .I (I18617));
INVX1 gate5092(.O (I18620), .I (g11385));
INVX1 gate5093(.O (g11548), .I (I18620));
INVX1 gate5094(.O (I18623), .I (g11003));
INVX1 gate5095(.O (g11549), .I (I18623));
INVX1 gate5096(.O (I18626), .I (g8649));
INVX1 gate5097(.O (g11550), .I (I18626));
INVX1 gate5098(.O (I18629), .I (g8811));
INVX1 gate5099(.O (g11551), .I (I18629));
INVX1 gate5100(.O (I18632), .I (g8850));
INVX1 gate5101(.O (g11552), .I (I18632));
INVX1 gate5102(.O (I18635), .I (g8904));
INVX1 gate5103(.O (g11553), .I (I18635));
INVX1 gate5104(.O (I18638), .I (g8826));
INVX1 gate5105(.O (g11554), .I (I18638));
INVX1 gate5106(.O (I18641), .I (g8871));
INVX1 gate5107(.O (g11555), .I (I18641));
INVX1 gate5108(.O (I18644), .I (g8937));
INVX1 gate5109(.O (g11556), .I (I18644));
INVX1 gate5110(.O (I18647), .I (g8851));
INVX1 gate5111(.O (g11557), .I (I18647));
INVX1 gate5112(.O (I18650), .I (g8905));
INVX1 gate5113(.O (g11558), .I (I18650));
INVX1 gate5114(.O (I18653), .I (g8971));
INVX1 gate5115(.O (g11559), .I (I18653));
INVX1 gate5116(.O (I18656), .I (g8872));
INVX1 gate5117(.O (g11560), .I (I18656));
INVX1 gate5118(.O (I18659), .I (g8938));
INVX1 gate5119(.O (g11561), .I (I18659));
INVX1 gate5120(.O (I18662), .I (g8996));
INVX1 gate5121(.O (g11562), .I (I18662));
INVX1 gate5122(.O (I18665), .I (g8689));
INVX1 gate5123(.O (g11563), .I (I18665));
INVX1 gate5124(.O (I18668), .I (g8756));
INVX1 gate5125(.O (g11564), .I (I18668));
INVX1 gate5126(.O (I18671), .I (g8812));
INVX1 gate5127(.O (g11565), .I (I18671));
INVX1 gate5128(.O (I18674), .I (g9487));
INVX1 gate5129(.O (g11566), .I (I18674));
INVX1 gate5130(.O (I18677), .I (g8908));
INVX1 gate5131(.O (g11567), .I (I18677));
INVX1 gate5132(.O (I18680), .I (g8973));
INVX1 gate5133(.O (g11568), .I (I18680));
INVX1 gate5134(.O (I18683), .I (g9733));
INVX1 gate5135(.O (g11569), .I (I18683));
INVX1 gate5136(.O (I18686), .I (g9932));
INVX1 gate5137(.O (g11570), .I (I18686));
INVX1 gate5138(.O (I18689), .I (g10231));
INVX1 gate5139(.O (g11571), .I (I18689));
INVX1 gate5140(.O (I18692), .I (g10935));
INVX1 gate5141(.O (g11572), .I (I18692));
INVX1 gate5142(.O (I18695), .I (g11054));
INVX1 gate5143(.O (g11573), .I (I18695));
INVX1 gate5144(.O (I18698), .I (g11255));
INVX1 gate5145(.O (g11574), .I (I18698));
INVX1 gate5146(.O (I18701), .I (g11471));
INVX1 gate5147(.O (g11575), .I (I18701));
INVX1 gate5148(.O (I18704), .I (g11055));
INVX1 gate5149(.O (g11576), .I (I18704));
INVX1 gate5150(.O (I18707), .I (g8665));
INVX1 gate5151(.O (g11577), .I (I18707));
INVX1 gate5152(.O (I18710), .I (g8827));
INVX1 gate5153(.O (g11578), .I (I18710));
INVX1 gate5154(.O (I18713), .I (g8877));
INVX1 gate5155(.O (g11579), .I (I18713));
INVX1 gate5156(.O (I18716), .I (g8944));
INVX1 gate5157(.O (g11580), .I (I18716));
INVX1 gate5158(.O (I18719), .I (g8852));
INVX1 gate5159(.O (g11581), .I (I18719));
INVX1 gate5160(.O (I18722), .I (g8909));
INVX1 gate5161(.O (g11582), .I (I18722));
INVX1 gate5162(.O (I18725), .I (g8977));
INVX1 gate5163(.O (g11583), .I (I18725));
INVX1 gate5164(.O (I18728), .I (g8878));
INVX1 gate5165(.O (g11584), .I (I18728));
INVX1 gate5166(.O (I18731), .I (g8945));
INVX1 gate5167(.O (g11585), .I (I18731));
INVX1 gate5168(.O (I18734), .I (g9003));
INVX1 gate5169(.O (g11586), .I (I18734));
INVX1 gate5170(.O (I18737), .I (g8910));
INVX1 gate5171(.O (g11587), .I (I18737));
INVX1 gate5172(.O (I18740), .I (g8978));
INVX1 gate5173(.O (g11588), .I (I18740));
INVX1 gate5174(.O (I18743), .I (g9025));
INVX1 gate5175(.O (g11589), .I (I18743));
INVX1 gate5176(.O (I18746), .I (g8707));
INVX1 gate5177(.O (g11590), .I (I18746));
INVX1 gate5178(.O (I18749), .I (g8779));
INVX1 gate5179(.O (g11591), .I (I18749));
INVX1 gate5180(.O (I18752), .I (g8828));
INVX1 gate5181(.O (g11592), .I (I18752));
INVX1 gate5182(.O (I18755), .I (g9629));
INVX1 gate5183(.O (g11593), .I (I18755));
INVX1 gate5184(.O (I18758), .I (g8948));
INVX1 gate5185(.O (g11594), .I (I18758));
INVX1 gate5186(.O (I18761), .I (g9005));
INVX1 gate5187(.O (g11595), .I (I18761));
INVX1 gate5188(.O (I18764), .I (g9879));
INVX1 gate5189(.O (g11596), .I (I18764));
INVX1 gate5190(.O (I18767), .I (g10086));
INVX1 gate5191(.O (g11597), .I (I18767));
INVX1 gate5192(.O (I18770), .I (g10333));
INVX1 gate5193(.O (g11598), .I (I18770));
INVX1 gate5194(.O (I18773), .I (g10830));
INVX1 gate5195(.O (g11599), .I (I18773));
INVX1 gate5196(.O (I18777), .I (g9050));
INVX1 gate5197(.O (g11603), .I (I18777));
INVX1 gate5198(.O (I18780), .I (g10870));
INVX1 gate5199(.O (g11606), .I (I18780));
INVX1 gate5200(.O (I18784), .I (g9067));
INVX1 gate5201(.O (g11608), .I (I18784));
INVX1 gate5202(.O (I18787), .I (g10910));
INVX1 gate5203(.O (g11611), .I (I18787));
INVX1 gate5204(.O (I18791), .I (g9084));
INVX1 gate5205(.O (g11613), .I (I18791));
INVX1 gate5206(.O (I18794), .I (g10973));
INVX1 gate5207(.O (g11616), .I (I18794));
INVX1 gate5208(.O (g11620), .I (g10601));
INVX1 gate5209(.O (g11623), .I (g10961));
INVX1 gate5210(.O (I18810), .I (g10813));
INVX1 gate5211(.O (g11628), .I (I18810));
INVX1 gate5212(.O (I18813), .I (g10850));
INVX1 gate5213(.O (g11629), .I (I18813));
INVX1 gate5214(.O (I18817), .I (g9067));
INVX1 gate5215(.O (g11633), .I (I18817));
INVX1 gate5216(.O (I18820), .I (g10890));
INVX1 gate5217(.O (g11636), .I (I18820));
INVX1 gate5218(.O (I18824), .I (g9084));
INVX1 gate5219(.O (g11638), .I (I18824));
INVX1 gate5220(.O (I18827), .I (g10936));
INVX1 gate5221(.O (g11641), .I (I18827));
INVX1 gate5222(.O (g11642), .I (g10646));
INVX1 gate5223(.O (I18835), .I (g10834));
INVX1 gate5224(.O (g11651), .I (I18835));
INVX1 gate5225(.O (I18838), .I (g10871));
INVX1 gate5226(.O (g11652), .I (I18838));
INVX1 gate5227(.O (I18842), .I (g9084));
INVX1 gate5228(.O (g11656), .I (I18842));
INVX1 gate5229(.O (I18845), .I (g10911));
INVX1 gate5230(.O (g11659), .I (I18845));
INVX1 gate5231(.O (I18854), .I (g10854));
INVX1 gate5232(.O (g11670), .I (I18854));
INVX1 gate5233(.O (I18857), .I (g10891));
INVX1 gate5234(.O (g11671), .I (I18857));
INVX1 gate5235(.O (I18866), .I (g10875));
INVX1 gate5236(.O (g11682), .I (I18866));
INVX1 gate5237(.O (g11706), .I (g10928));
INVX1 gate5238(.O (g11732), .I (g10826));
INVX1 gate5239(.O (g11734), .I (g10843));
INVX1 gate5240(.O (g11735), .I (g10859));
INVX1 gate5241(.O (g11736), .I (g10862));
INVX1 gate5242(.O (g11737), .I (g10809));
INVX1 gate5243(.O (g11740), .I (g10877));
INVX1 gate5244(.O (g11741), .I (g10880));
INVX1 gate5245(.O (g11742), .I (g10883));
INVX1 gate5246(.O (g11743), .I (g8530));
INVX1 gate5247(.O (g11745), .I (g10892));
INVX1 gate5248(.O (g11746), .I (g10895));
INVX1 gate5249(.O (g11747), .I (g10898));
INVX1 gate5250(.O (g11748), .I (g10901));
INVX1 gate5251(.O (I18929), .I (g10711));
INVX1 gate5252(.O (g11749), .I (I18929));
INVX1 gate5253(.O (g11758), .I (g8514));
INVX1 gate5254(.O (g11761), .I (g10912));
INVX1 gate5255(.O (g11762), .I (g10915));
INVX1 gate5256(.O (g11763), .I (g10918));
INVX1 gate5257(.O (g11764), .I (g10921));
INVX1 gate5258(.O (g11765), .I (g10924));
INVX1 gate5259(.O (g11766), .I (g10886));
INVX1 gate5260(.O (I18943), .I (g9149));
INVX1 gate5261(.O (g11769), .I (I18943));
INVX1 gate5262(.O (g11770), .I (g10932));
INVX1 gate5263(.O (g11774), .I (g10937));
INVX1 gate5264(.O (g11775), .I (g10940));
INVX1 gate5265(.O (g11776), .I (g10943));
INVX1 gate5266(.O (g11777), .I (g10946));
INVX1 gate5267(.O (g11778), .I (g10949));
INVX1 gate5268(.O (g11779), .I (g10906));
INVX1 gate5269(.O (g11782), .I (g10963));
INVX1 gate5270(.O (g11783), .I (g10966));
INVX1 gate5271(.O (I18962), .I (g9159));
INVX1 gate5272(.O (g11786), .I (I18962));
INVX1 gate5273(.O (g11787), .I (g10969));
INVX1 gate5274(.O (I18969), .I (g8726));
INVX1 gate5275(.O (g11791), .I (I18969));
INVX1 gate5276(.O (g11794), .I (g10974));
INVX1 gate5277(.O (g11795), .I (g10977));
INVX1 gate5278(.O (g11796), .I (g10980));
INVX1 gate5279(.O (g11797), .I (g10983));
INVX1 gate5280(.O (g11798), .I (g10867));
INVX1 gate5281(.O (g11801), .I (g10988));
INVX1 gate5282(.O (g11802), .I (g10991));
INVX1 gate5283(.O (g11803), .I (g10994));
INVX1 gate5284(.O (g11804), .I (g10995));
INVX1 gate5285(.O (g11808), .I (g10996));
INVX1 gate5286(.O (g11809), .I (g10999));
INVX1 gate5287(.O (I18990), .I (g9183));
INVX1 gate5288(.O (g11812), .I (I18990));
INVX1 gate5289(.O (g11813), .I (g11004));
INVX1 gate5290(.O (g11817), .I (g11008));
INVX1 gate5291(.O (g11818), .I (g11011));
INVX1 gate5292(.O (g11819), .I (g11014));
INVX1 gate5293(.O (g11820), .I (g11017));
INVX1 gate5294(.O (g11821), .I (g10848));
INVX1 gate5295(.O (g11824), .I (g11022));
INVX1 gate5296(.O (g11825), .I (g11025));
INVX1 gate5297(.O (g11826), .I (g11028));
INVX1 gate5298(.O (g11827), .I (g11032));
INVX1 gate5299(.O (g11829), .I (g11035));
INVX1 gate5300(.O (g11834), .I (g11036));
INVX1 gate5301(.O (g11835), .I (g11039));
INVX1 gate5302(.O (g11836), .I (g11042));
INVX1 gate5303(.O (g11837), .I (g11045));
INVX1 gate5304(.O (g11841), .I (g11048));
INVX1 gate5305(.O (g11842), .I (g11051));
INVX1 gate5306(.O (I19025), .I (g9225));
INVX1 gate5307(.O (g11845), .I (I19025));
INVX1 gate5308(.O (g11846), .I (g11056));
INVX1 gate5309(.O (I19030), .I (g8726));
INVX1 gate5310(.O (g11848), .I (I19030));
INVX1 gate5311(.O (g11852), .I (g11063));
INVX1 gate5312(.O (g11853), .I (g11066));
INVX1 gate5313(.O (g11854), .I (g11078));
INVX1 gate5314(.O (g11856), .I (g11079));
INVX1 gate5315(.O (g11857), .I (g11082));
INVX1 gate5316(.O (g11858), .I (g11085));
INVX1 gate5317(.O (g11859), .I (g11088));
INVX1 gate5318(.O (g11862), .I (g11091));
INVX1 gate5319(.O (g11866), .I (g11092));
INVX1 gate5320(.O (g11867), .I (g11095));
INVX1 gate5321(.O (g11868), .I (g11098));
INVX1 gate5322(.O (g11869), .I (g11102));
INVX1 gate5323(.O (g11871), .I (g11105));
INVX1 gate5324(.O (g11876), .I (g11108));
INVX1 gate5325(.O (g11877), .I (g11111));
INVX1 gate5326(.O (g11878), .I (g11114));
INVX1 gate5327(.O (g11879), .I (g11117));
INVX1 gate5328(.O (g11883), .I (g11120));
INVX1 gate5329(.O (g11884), .I (g11123));
INVX1 gate5330(.O (g11886), .I (g11126));
INVX1 gate5331(.O (g11887), .I (g11129));
INVX1 gate5332(.O (g11888), .I (g11021));
INVX1 gate5333(.O (g11891), .I (g11132));
INVX1 gate5334(.O (g11892), .I (g11135));
INVX1 gate5335(.O (g11893), .I (g11138));
INVX1 gate5336(.O (g11894), .I (g11141));
INVX1 gate5337(.O (g11895), .I (g11144));
INVX1 gate5338(.O (g11898), .I (g11145));
INVX1 gate5339(.O (g11899), .I (g11148));
INVX1 gate5340(.O (g11900), .I (g11151));
INVX1 gate5341(.O (g11901), .I (g11154));
INVX1 gate5342(.O (g11904), .I (g11157));
INVX1 gate5343(.O (g11908), .I (g11160));
INVX1 gate5344(.O (g11909), .I (g11163));
INVX1 gate5345(.O (g11910), .I (g11166));
INVX1 gate5346(.O (g11911), .I (g11170));
INVX1 gate5347(.O (g11913), .I (g11173));
INVX1 gate5348(.O (g11918), .I (g11176));
INVX1 gate5349(.O (g11919), .I (g11179));
INVX1 gate5350(.O (g11920), .I (g11182));
INVX1 gate5351(.O (g11921), .I (g11185));
INVX1 gate5352(.O (I19105), .I (g8726));
INVX1 gate5353(.O (g11923), .I (I19105));
INVX1 gate5354(.O (g11927), .I (g10987));
INVX1 gate5355(.O (g11929), .I (g11199));
INVX1 gate5356(.O (g11930), .I (g11202));
INVX1 gate5357(.O (g11931), .I (g11205));
INVX1 gate5358(.O (g11932), .I (g11209));
INVX1 gate5359(.O (g11933), .I (g11210));
INVX1 gate5360(.O (g11936), .I (g11213));
INVX1 gate5361(.O (I19119), .I (g9202));
INVX1 gate5362(.O (g11937), .I (I19119));
INVX1 gate5363(.O (g11941), .I (g11216));
INVX1 gate5364(.O (g11942), .I (g11219));
INVX1 gate5365(.O (g11943), .I (g11222));
INVX1 gate5366(.O (g11944), .I (g11225));
INVX1 gate5367(.O (g11945), .I (g11228));
INVX1 gate5368(.O (g11948), .I (g11231));
INVX1 gate5369(.O (g11949), .I (g11234));
INVX1 gate5370(.O (g11950), .I (g11237));
INVX1 gate5371(.O (g11951), .I (g11240));
INVX1 gate5372(.O (g11954), .I (g11243));
INVX1 gate5373(.O (g11958), .I (g11246));
INVX1 gate5374(.O (g11959), .I (g11249));
INVX1 gate5375(.O (g11960), .I (g11252));
INVX1 gate5376(.O (g11961), .I (g11256));
INVX1 gate5377(.O (g11963), .I (g11259));
INVX1 gate5378(.O (g11968), .I (g11265));
INVX1 gate5379(.O (g11969), .I (g11268));
INVX1 gate5380(.O (g11970), .I (g11271));
INVX1 gate5381(.O (g11971), .I (g11274));
INVX1 gate5382(.O (g11972), .I (g11277));
INVX1 gate5383(.O (g11973), .I (g11278));
INVX1 gate5384(.O (I19160), .I (g10549));
INVX1 gate5385(.O (g11976), .I (I19160));
INVX1 gate5386(.O (g11982), .I (g11281));
INVX1 gate5387(.O (g11983), .I (g11284));
INVX1 gate5388(.O (g11984), .I (g11287));
INVX1 gate5389(.O (g11985), .I (g11291));
INVX1 gate5390(.O (g11986), .I (g11294));
INVX1 gate5391(.O (g11989), .I (g11297));
INVX1 gate5392(.O (I19174), .I (g9263));
INVX1 gate5393(.O (g11990), .I (I19174));
INVX1 gate5394(.O (g11994), .I (g11300));
INVX1 gate5395(.O (g11995), .I (g11303));
INVX1 gate5396(.O (g11996), .I (g11306));
INVX1 gate5397(.O (g11997), .I (g11309));
INVX1 gate5398(.O (g11998), .I (g11312));
INVX1 gate5399(.O (g12001), .I (g11315));
INVX1 gate5400(.O (g12002), .I (g11318));
INVX1 gate5401(.O (g12003), .I (g11321));
INVX1 gate5402(.O (g12004), .I (g11324));
INVX1 gate5403(.O (g12007), .I (g11327));
INVX1 gate5404(.O (I19195), .I (g8726));
INVX1 gate5405(.O (g12009), .I (I19195));
INVX1 gate5406(.O (g12013), .I (g10772));
INVX1 gate5407(.O (g12017), .I (g10100));
INVX1 gate5408(.O (g12020), .I (g11341));
INVX1 gate5409(.O (g12021), .I (g11344));
INVX1 gate5410(.O (g12022), .I (g11348));
INVX1 gate5411(.O (g12023), .I (g11351));
INVX1 gate5412(.O (g12024), .I (g11354));
INVX1 gate5413(.O (g12025), .I (g11355));
INVX1 gate5414(.O (I19208), .I (g10424));
INVX1 gate5415(.O (g12027), .I (I19208));
INVX1 gate5416(.O (I19211), .I (g10486));
INVX1 gate5417(.O (g12030), .I (I19211));
INVX1 gate5418(.O (g12037), .I (g11358));
INVX1 gate5419(.O (g12038), .I (g11361));
INVX1 gate5420(.O (g12039), .I (g11364));
INVX1 gate5421(.O (g12040), .I (g11367));
INVX1 gate5422(.O (g12041), .I (g11370));
INVX1 gate5423(.O (g12042), .I (g11373));
INVX1 gate5424(.O (I19226), .I (g10606));
INVX1 gate5425(.O (g12045), .I (I19226));
INVX1 gate5426(.O (g12051), .I (g11376));
INVX1 gate5427(.O (g12052), .I (g11379));
INVX1 gate5428(.O (g12053), .I (g11382));
INVX1 gate5429(.O (g12054), .I (g11386));
INVX1 gate5430(.O (g12055), .I (g11389));
INVX1 gate5431(.O (g12058), .I (g11392));
INVX1 gate5432(.O (I19240), .I (g9341));
INVX1 gate5433(.O (g12059), .I (I19240));
INVX1 gate5434(.O (g12063), .I (g11395));
INVX1 gate5435(.O (g12064), .I (g11398));
INVX1 gate5436(.O (g12065), .I (g11401));
INVX1 gate5437(.O (g12066), .I (g11404));
INVX1 gate5438(.O (g12067), .I (g11407));
INVX1 gate5439(.O (g12071), .I (g10783));
INVX1 gate5440(.O (g12075), .I (g11411));
INVX1 gate5441(.O (g12076), .I (g11414));
INVX1 gate5442(.O (g12077), .I (g11417));
INVX1 gate5443(.O (g12078), .I (g11422));
INVX1 gate5444(.O (g12084), .I (g11425));
INVX1 gate5445(.O (g12085), .I (g11428));
INVX1 gate5446(.O (g12086), .I (g11432));
INVX1 gate5447(.O (g12087), .I (g11435));
INVX1 gate5448(.O (g12088), .I (g11438));
INVX1 gate5449(.O (g12089), .I (g11441));
INVX1 gate5450(.O (I19271), .I (g10500));
INVX1 gate5451(.O (g12091), .I (I19271));
INVX1 gate5452(.O (I19274), .I (g10560));
INVX1 gate5453(.O (g12094), .I (I19274));
INVX1 gate5454(.O (g12101), .I (g11444));
INVX1 gate5455(.O (g12102), .I (g11447));
INVX1 gate5456(.O (g12103), .I (g11450));
INVX1 gate5457(.O (g12104), .I (g11453));
INVX1 gate5458(.O (g12105), .I (g11456));
INVX1 gate5459(.O (g12106), .I (g11459));
INVX1 gate5460(.O (I19289), .I (g10653));
INVX1 gate5461(.O (g12109), .I (I19289));
INVX1 gate5462(.O (g12115), .I (g11462));
INVX1 gate5463(.O (g12116), .I (g11465));
INVX1 gate5464(.O (g12117), .I (g11468));
INVX1 gate5465(.O (g12118), .I (g11472));
INVX1 gate5466(.O (g12119), .I (g11475));
INVX1 gate5467(.O (g12122), .I (g11478));
INVX1 gate5468(.O (I19303), .I (g9422));
INVX1 gate5469(.O (g12123), .I (I19303));
INVX1 gate5470(.O (I19307), .I (g8726));
INVX1 gate5471(.O (g12125), .I (I19307));
INVX1 gate5472(.O (g12130), .I (g10788));
INVX1 gate5473(.O (g12134), .I (g8321));
INVX1 gate5474(.O (g12135), .I (g8324));
INVX1 gate5475(.O (I19315), .I (g10424));
INVX1 gate5476(.O (g12136), .I (I19315));
INVX1 gate5477(.O (I19318), .I (g10486));
INVX1 gate5478(.O (g12139), .I (I19318));
INVX1 gate5479(.O (I19321), .I (g10549));
INVX1 gate5480(.O (g12142), .I (I19321));
INVX1 gate5481(.O (g12147), .I (g8330));
INVX1 gate5482(.O (g12148), .I (g8333));
INVX1 gate5483(.O (g12149), .I (g8336));
INVX1 gate5484(.O (g12150), .I (g8341));
INVX1 gate5485(.O (g12156), .I (g8344));
INVX1 gate5486(.O (g12157), .I (g8347));
INVX1 gate5487(.O (g12158), .I (g8351));
INVX1 gate5488(.O (g12159), .I (g8354));
INVX1 gate5489(.O (g12160), .I (g8357));
INVX1 gate5490(.O (g12161), .I (g8360));
INVX1 gate5491(.O (I19342), .I (g10574));
INVX1 gate5492(.O (g12163), .I (I19342));
INVX1 gate5493(.O (I19345), .I (g10617));
INVX1 gate5494(.O (g12166), .I (I19345));
INVX1 gate5495(.O (g12173), .I (g8363));
INVX1 gate5496(.O (g12174), .I (g8366));
INVX1 gate5497(.O (g12175), .I (g8369));
INVX1 gate5498(.O (g12176), .I (g8372));
INVX1 gate5499(.O (g12177), .I (g8375));
INVX1 gate5500(.O (g12178), .I (g8378));
INVX1 gate5501(.O (I19360), .I (g10683));
INVX1 gate5502(.O (g12181), .I (I19360));
INVX1 gate5503(.O (g12187), .I (g8285));
INVX1 gate5504(.O (g12191), .I (g8382));
INVX1 gate5505(.O (g12196), .I (g8388));
INVX1 gate5506(.O (g12197), .I (g8391));
INVX1 gate5507(.O (I19374), .I (g10500));
INVX1 gate5508(.O (g12198), .I (I19374));
INVX1 gate5509(.O (I19377), .I (g10560));
INVX1 gate5510(.O (g12201), .I (I19377));
INVX1 gate5511(.O (I19380), .I (g10606));
INVX1 gate5512(.O (g12204), .I (I19380));
INVX1 gate5513(.O (g12209), .I (g8397));
INVX1 gate5514(.O (g12210), .I (g8400));
INVX1 gate5515(.O (g12211), .I (g8403));
INVX1 gate5516(.O (g12212), .I (g8408));
INVX1 gate5517(.O (g12218), .I (g8411));
INVX1 gate5518(.O (g12219), .I (g8414));
INVX1 gate5519(.O (g12220), .I (g8418));
INVX1 gate5520(.O (g12221), .I (g8421));
INVX1 gate5521(.O (g12222), .I (g8424));
INVX1 gate5522(.O (g12223), .I (g8427));
INVX1 gate5523(.O (I19401), .I (g10631));
INVX1 gate5524(.O (g12225), .I (I19401));
INVX1 gate5525(.O (I19404), .I (g10664));
INVX1 gate5526(.O (g12228), .I (I19404));
INVX1 gate5527(.O (g12235), .I (g8294));
INVX1 gate5528(.O (I19412), .I (g10486));
INVX1 gate5529(.O (g12239), .I (I19412));
INVX1 gate5530(.O (I19415), .I (g10549));
INVX1 gate5531(.O (g12242), .I (I19415));
INVX1 gate5532(.O (g12246), .I (g8434));
INVX1 gate5533(.O (g12251), .I (g8440));
INVX1 gate5534(.O (g12252), .I (g8443));
INVX1 gate5535(.O (I19426), .I (g10574));
INVX1 gate5536(.O (g12253), .I (I19426));
INVX1 gate5537(.O (I19429), .I (g10617));
INVX1 gate5538(.O (g12256), .I (I19429));
INVX1 gate5539(.O (I19432), .I (g10653));
INVX1 gate5540(.O (g12259), .I (I19432));
INVX1 gate5541(.O (g12264), .I (g8449));
INVX1 gate5542(.O (g12265), .I (g8452));
INVX1 gate5543(.O (g12266), .I (g8455));
INVX1 gate5544(.O (g12267), .I (g8460));
INVX1 gate5545(.O (g12275), .I (g8303));
INVX1 gate5546(.O (I19449), .I (g10424));
INVX1 gate5547(.O (g12279), .I (I19449));
INVX1 gate5548(.O (I19452), .I (g10560));
INVX1 gate5549(.O (g12282), .I (I19452));
INVX1 gate5550(.O (I19455), .I (g10606));
INVX1 gate5551(.O (g12285), .I (I19455));
INVX1 gate5552(.O (g12289), .I (g8469));
INVX1 gate5553(.O (g12294), .I (g8475));
INVX1 gate5554(.O (g12295), .I (g8478));
INVX1 gate5555(.O (I19466), .I (g10631));
INVX1 gate5556(.O (g12296), .I (I19466));
INVX1 gate5557(.O (I19469), .I (g10664));
INVX1 gate5558(.O (g12299), .I (I19469));
INVX1 gate5559(.O (I19472), .I (g10683));
INVX1 gate5560(.O (g12302), .I (I19472));
INVX1 gate5561(.O (g12308), .I (g8312));
INVX1 gate5562(.O (I19479), .I (g10549));
INVX1 gate5563(.O (g12312), .I (I19479));
INVX1 gate5564(.O (I19482), .I (g10500));
INVX1 gate5565(.O (g12315), .I (I19482));
INVX1 gate5566(.O (I19485), .I (g10617));
INVX1 gate5567(.O (g12318), .I (I19485));
INVX1 gate5568(.O (I19488), .I (g10653));
INVX1 gate5569(.O (g12321), .I (I19488));
INVX1 gate5570(.O (g12325), .I (g8494));
INVX1 gate5571(.O (g12332), .I (g10829));
INVX1 gate5572(.O (I19500), .I (g10424));
INVX1 gate5573(.O (g12333), .I (I19500));
INVX1 gate5574(.O (I19503), .I (g10486));
INVX1 gate5575(.O (g12336), .I (I19503));
INVX1 gate5576(.O (I19507), .I (g10606));
INVX1 gate5577(.O (g12340), .I (I19507));
INVX1 gate5578(.O (I19510), .I (g10574));
INVX1 gate5579(.O (g12343), .I (I19510));
INVX1 gate5580(.O (I19513), .I (g10664));
INVX1 gate5581(.O (g12346), .I (I19513));
INVX1 gate5582(.O (I19516), .I (g10683));
INVX1 gate5583(.O (g12349), .I (I19516));
INVX1 gate5584(.O (g12354), .I (g8381));
INVX1 gate5585(.O (g12362), .I (g10866));
INVX1 gate5586(.O (I19523), .I (g10500));
INVX1 gate5587(.O (g12363), .I (I19523));
INVX1 gate5588(.O (I19526), .I (g10560));
INVX1 gate5589(.O (g12366), .I (I19526));
INVX1 gate5590(.O (I19530), .I (g10653));
INVX1 gate5591(.O (g12370), .I (I19530));
INVX1 gate5592(.O (I19533), .I (g10631));
INVX1 gate5593(.O (g12373), .I (I19533));
INVX1 gate5594(.O (g12378), .I (g10847));
INVX1 gate5595(.O (I19539), .I (g10549));
INVX1 gate5596(.O (g12379), .I (I19539));
INVX1 gate5597(.O (I19542), .I (g10574));
INVX1 gate5598(.O (g12382), .I (I19542));
INVX1 gate5599(.O (I19545), .I (g10617));
INVX1 gate5600(.O (g12385), .I (I19545));
INVX1 gate5601(.O (I19549), .I (g10683));
INVX1 gate5602(.O (g12389), .I (I19549));
INVX1 gate5603(.O (I19552), .I (g8430));
INVX1 gate5604(.O (g12392), .I (I19552));
INVX1 gate5605(.O (g12408), .I (g11020));
INVX1 gate5606(.O (I19557), .I (g10606));
INVX1 gate5607(.O (g12409), .I (I19557));
INVX1 gate5608(.O (I19560), .I (g10631));
INVX1 gate5609(.O (g12412), .I (I19560));
INVX1 gate5610(.O (I19563), .I (g10664));
INVX1 gate5611(.O (g12415), .I (I19563));
INVX1 gate5612(.O (g12420), .I (g10986));
INVX1 gate5613(.O (I19569), .I (g10653));
INVX1 gate5614(.O (g12421), .I (I19569));
INVX1 gate5615(.O (g12424), .I (g10962));
INVX1 gate5616(.O (I19573), .I (g8835));
INVX1 gate5617(.O (g12425), .I (I19573));
INVX1 gate5618(.O (I19576), .I (g10683));
INVX1 gate5619(.O (g12426), .I (I19576));
INVX1 gate5620(.O (g12430), .I (g10905));
INVX1 gate5621(.O (I19582), .I (g8862));
INVX1 gate5622(.O (g12432), .I (I19582));
INVX1 gate5623(.O (g12434), .I (g10929));
INVX1 gate5624(.O (I19587), .I (g9173));
INVX1 gate5625(.O (g12435), .I (I19587));
INVX1 gate5626(.O (I19591), .I (g8900));
INVX1 gate5627(.O (g12437), .I (I19591));
INVX1 gate5628(.O (g12438), .I (g10846));
INVX1 gate5629(.O (I19595), .I (g10810));
INVX1 gate5630(.O (g12439), .I (I19595));
INVX1 gate5631(.O (I19598), .I (g9215));
INVX1 gate5632(.O (g12440), .I (I19598));
INVX1 gate5633(.O (I19602), .I (g8940));
INVX1 gate5634(.O (g12442), .I (I19602));
INVX1 gate5635(.O (I19605), .I (g10797));
INVX1 gate5636(.O (g12443), .I (I19605));
INVX1 gate5637(.O (I19608), .I (g10831));
INVX1 gate5638(.O (g12444), .I (I19608));
INVX1 gate5639(.O (I19611), .I (g9276));
INVX1 gate5640(.O (g12445), .I (I19611));
INVX1 gate5641(.O (I19615), .I (g10789));
INVX1 gate5642(.O (g12447), .I (I19615));
INVX1 gate5643(.O (I19618), .I (g10814));
INVX1 gate5644(.O (g12448), .I (I19618));
INVX1 gate5645(.O (I19621), .I (g10851));
INVX1 gate5646(.O (g12449), .I (I19621));
INVX1 gate5647(.O (I19624), .I (g9354));
INVX1 gate5648(.O (g12450), .I (I19624));
INVX1 gate5649(.O (I19628), .I (g10784));
INVX1 gate5650(.O (g12452), .I (I19628));
INVX1 gate5651(.O (I19631), .I (g10801));
INVX1 gate5652(.O (g12453), .I (I19631));
INVX1 gate5653(.O (I19634), .I (g10835));
INVX1 gate5654(.O (g12454), .I (I19634));
INVX1 gate5655(.O (I19637), .I (g10872));
INVX1 gate5656(.O (g12455), .I (I19637));
INVX1 gate5657(.O (g12456), .I (g8602));
INVX1 gate5658(.O (I19642), .I (g10793));
INVX1 gate5659(.O (g12460), .I (I19642));
INVX1 gate5660(.O (I19645), .I (g10818));
INVX1 gate5661(.O (g12461), .I (I19645));
INVX1 gate5662(.O (I19648), .I (g10855));
INVX1 gate5663(.O (g12462), .I (I19648));
INVX1 gate5664(.O (g12463), .I (g10730));
INVX1 gate5665(.O (g12466), .I (g8614));
INVX1 gate5666(.O (I19654), .I (g10805));
INVX1 gate5667(.O (g12470), .I (I19654));
INVX1 gate5668(.O (I19657), .I (g10839));
INVX1 gate5669(.O (g12471), .I (I19657));
INVX1 gate5670(.O (g12472), .I (g8617));
INVX1 gate5671(.O (g12473), .I (g8580));
INVX1 gate5672(.O (g12476), .I (g8622));
INVX1 gate5673(.O (g12478), .I (g10749));
INVX1 gate5674(.O (g12481), .I (g8627));
INVX1 gate5675(.O (I19667), .I (g10822));
INVX1 gate5676(.O (g12485), .I (I19667));
INVX1 gate5677(.O (g12490), .I (g8587));
INVX1 gate5678(.O (g12493), .I (g8632));
INVX1 gate5679(.O (g12495), .I (g10767));
INVX1 gate5680(.O (g12498), .I (g8637));
INVX1 gate5681(.O (g12502), .I (g8640));
INVX1 gate5682(.O (g12504), .I (g8643));
INVX1 gate5683(.O (g12505), .I (g8646));
INVX1 gate5684(.O (g12510), .I (g8594));
INVX1 gate5685(.O (g12513), .I (g8651));
INVX1 gate5686(.O (g12515), .I (g10773));
INVX1 gate5687(.O (g12518), .I (g8655));
INVX1 gate5688(.O (I19689), .I (g10016));
INVX1 gate5689(.O (g12519), .I (I19689));
INVX1 gate5690(.O (g12521), .I (g8659));
INVX1 gate5691(.O (g12522), .I (g8662));
INVX1 gate5692(.O (g12527), .I (g8605));
INVX1 gate5693(.O (g12530), .I (g8667));
INVX1 gate5694(.O (g12532), .I (g8670));
INVX1 gate5695(.O (g12533), .I (g8673));
INVX1 gate5696(.O (I19702), .I (g10125));
INVX1 gate5697(.O (g12534), .I (I19702));
INVX1 gate5698(.O (g12536), .I (g8678));
INVX1 gate5699(.O (g12537), .I (g8681));
INVX1 gate5700(.O (g12542), .I (g8684));
INVX1 gate5701(.O (I19711), .I (g10230));
INVX1 gate5702(.O (g12543), .I (I19711));
INVX1 gate5703(.O (g12545), .I (g8690));
INVX1 gate5704(.O (g12546), .I (g8693));
INVX1 gate5705(.O (g12547), .I (g8696));
INVX1 gate5706(.O (I19718), .I (g8726));
INVX1 gate5707(.O (g12548), .I (I19718));
INVX1 gate5708(.O (g12551), .I (g8700));
INVX1 gate5709(.O (I19722), .I (g10332));
INVX1 gate5710(.O (g12552), .I (I19722));
INVX1 gate5711(.O (g12553), .I (g8708));
INVX1 gate5712(.O (g12554), .I (g8711));
INVX1 gate5713(.O (I19727), .I (g8726));
INVX1 gate5714(.O (g12555), .I (I19727));
INVX1 gate5715(.O (g12558), .I (g8714));
INVX1 gate5716(.O (g12559), .I (g8719));
INVX1 gate5717(.O (g12560), .I (g8745));
INVX1 gate5718(.O (I19733), .I (g8726));
INVX1 gate5719(.O (g12561), .I (I19733));
INVX1 gate5720(.O (I19736), .I (g9184));
INVX1 gate5721(.O (g12564), .I (I19736));
INVX1 gate5722(.O (I19739), .I (g10694));
INVX1 gate5723(.O (g12565), .I (I19739));
INVX1 gate5724(.O (g12596), .I (g8748));
INVX1 gate5725(.O (g12597), .I (g8752));
INVX1 gate5726(.O (g12598), .I (g8757));
INVX1 gate5727(.O (g12599), .I (g8763));
INVX1 gate5728(.O (g12600), .I (g8766));
INVX1 gate5729(.O (I19747), .I (g8726));
INVX1 gate5730(.O (g12601), .I (I19747));
INVX1 gate5731(.O (I19750), .I (g8726));
INVX1 gate5732(.O (g12604), .I (I19750));
INVX1 gate5733(.O (I19753), .I (g9229));
INVX1 gate5734(.O (g12607), .I (I19753));
INVX1 gate5735(.O (I19756), .I (g10424));
INVX1 gate5736(.O (g12608), .I (I19756));
INVX1 gate5737(.O (I19759), .I (g10714));
INVX1 gate5738(.O (g12611), .I (I19759));
INVX1 gate5739(.O (g12642), .I (g8771));
INVX1 gate5740(.O (g12643), .I (g8775));
INVX1 gate5741(.O (g12644), .I (g8780));
INVX1 gate5742(.O (g12645), .I (g8785));
INVX1 gate5743(.O (g12646), .I (g8788));
INVX1 gate5744(.O (I19767), .I (g8726));
INVX1 gate5745(.O (g12647), .I (I19767));
INVX1 gate5746(.O (I19771), .I (g10038));
INVX1 gate5747(.O (g12651), .I (I19771));
INVX1 gate5748(.O (I19774), .I (g10500));
INVX1 gate5749(.O (g12654), .I (I19774));
INVX1 gate5750(.O (I19777), .I (g10735));
INVX1 gate5751(.O (g12657), .I (I19777));
INVX1 gate5752(.O (g12688), .I (g8794));
INVX1 gate5753(.O (g12689), .I (g8798));
INVX1 gate5754(.O (g12690), .I (g8802));
INVX1 gate5755(.O (g12691), .I (g8805));
INVX1 gate5756(.O (I19784), .I (g8726));
INVX1 gate5757(.O (g12692), .I (I19784));
INVX1 gate5758(.O (I19787), .I (g8726));
INVX1 gate5759(.O (g12695), .I (I19787));
INVX1 gate5760(.O (I19791), .I (g10486));
INVX1 gate5761(.O (g12699), .I (I19791));
INVX1 gate5762(.O (I19794), .I (g10676));
INVX1 gate5763(.O (g12702), .I (I19794));
INVX1 gate5764(.O (I19797), .I (g10147));
INVX1 gate5765(.O (g12705), .I (I19797));
INVX1 gate5766(.O (I19800), .I (g10574));
INVX1 gate5767(.O (g12708), .I (I19800));
INVX1 gate5768(.O (I19803), .I (g10754));
INVX1 gate5769(.O (g12711), .I (I19803));
INVX1 gate5770(.O (g12742), .I (g8813));
INVX1 gate5771(.O (g12743), .I (g8817));
INVX1 gate5772(.O (I19808), .I (g8726));
INVX1 gate5773(.O (g12744), .I (I19808));
INVX1 gate5774(.O (g12748), .I (g8823));
INVX1 gate5775(.O (I19813), .I (g10649));
INVX1 gate5776(.O (g12749), .I (I19813));
INVX1 gate5777(.O (I19816), .I (g10703));
INVX1 gate5778(.O (g12752), .I (I19816));
INVX1 gate5779(.O (I19820), .I (g10560));
INVX1 gate5780(.O (g12756), .I (I19820));
INVX1 gate5781(.O (I19823), .I (g10705));
INVX1 gate5782(.O (g12759), .I (I19823));
INVX1 gate5783(.O (I19826), .I (g10252));
INVX1 gate5784(.O (g12762), .I (I19826));
INVX1 gate5785(.O (I19829), .I (g10631));
INVX1 gate5786(.O (g12765), .I (I19829));
INVX1 gate5787(.O (g12768), .I (g8829));
INVX1 gate5788(.O (I19833), .I (g8726));
INVX1 gate5789(.O (g12769), .I (I19833));
INVX1 gate5790(.O (I19836), .I (g8726));
INVX1 gate5791(.O (g12772), .I (I19836));
INVX1 gate5792(.O (g12775), .I (g8832));
INVX1 gate5793(.O (g12776), .I (g10766));
INVX1 gate5794(.O (g12782), .I (g8836));
INVX1 gate5795(.O (I19844), .I (g8533));
INVX1 gate5796(.O (g12783), .I (I19844));
INVX1 gate5797(.O (I19847), .I (g10677));
INVX1 gate5798(.O (g12786), .I (I19847));
INVX1 gate5799(.O (g12790), .I (g8847));
INVX1 gate5800(.O (I19852), .I (g10679));
INVX1 gate5801(.O (g12791), .I (I19852));
INVX1 gate5802(.O (I19855), .I (g10723));
INVX1 gate5803(.O (g12794), .I (I19855));
INVX1 gate5804(.O (I19859), .I (g10617));
INVX1 gate5805(.O (g12798), .I (I19859));
INVX1 gate5806(.O (I19862), .I (g10725));
INVX1 gate5807(.O (g12801), .I (I19862));
INVX1 gate5808(.O (I19865), .I (g10354));
INVX1 gate5809(.O (g12804), .I (I19865));
INVX1 gate5810(.O (g12807), .I (g8853));
INVX1 gate5811(.O (I19869), .I (g8726));
INVX1 gate5812(.O (g12808), .I (I19869));
INVX1 gate5813(.O (I19872), .I (g8317));
INVX1 gate5814(.O (g12811), .I (I19872));
INVX1 gate5815(.O (g12815), .I (g8856));
INVX1 gate5816(.O (I19877), .I (g8547));
INVX1 gate5817(.O (g12816), .I (I19877));
INVX1 gate5818(.O (g12821), .I (g8863));
INVX1 gate5819(.O (I19883), .I (g8550));
INVX1 gate5820(.O (g12822), .I (I19883));
INVX1 gate5821(.O (I19886), .I (g10706));
INVX1 gate5822(.O (g12825), .I (I19886));
INVX1 gate5823(.O (g12829), .I (g8874));
INVX1 gate5824(.O (I19891), .I (g10708));
INVX1 gate5825(.O (g12830), .I (I19891));
INVX1 gate5826(.O (I19894), .I (g10744));
INVX1 gate5827(.O (g12833), .I (I19894));
INVX1 gate5828(.O (I19898), .I (g10664));
INVX1 gate5829(.O (g12837), .I (I19898));
INVX1 gate5830(.O (I19901), .I (g10746));
INVX1 gate5831(.O (g12840), .I (I19901));
INVX1 gate5832(.O (g12843), .I (g8879));
INVX1 gate5833(.O (I19905), .I (g8726));
INVX1 gate5834(.O (g12844), .I (I19905));
INVX1 gate5835(.O (g12847), .I (g8882));
INVX1 gate5836(.O (g12848), .I (g11059));
INVX1 gate5837(.O (g12850), .I (g8885));
INVX1 gate5838(.O (g12851), .I (g8888));
INVX1 gate5839(.O (g12853), .I (g8894));
INVX1 gate5840(.O (I19915), .I (g8560));
INVX1 gate5841(.O (g12854), .I (I19915));
INVX1 gate5842(.O (g12859), .I (g8901));
INVX1 gate5843(.O (I19921), .I (g8563));
INVX1 gate5844(.O (g12860), .I (I19921));
INVX1 gate5845(.O (I19924), .I (g10726));
INVX1 gate5846(.O (g12863), .I (I19924));
INVX1 gate5847(.O (g12867), .I (g8912));
INVX1 gate5848(.O (I19929), .I (g10728));
INVX1 gate5849(.O (g12868), .I (I19929));
INVX1 gate5850(.O (I19932), .I (g10763));
INVX1 gate5851(.O (g12871), .I (I19932));
INVX1 gate5852(.O (g12874), .I (g8915));
INVX1 gate5853(.O (g12875), .I (g10779));
INVX1 gate5854(.O (g12881), .I (g8918));
INVX1 gate5855(.O (g12882), .I (g8921));
INVX1 gate5856(.O (g12891), .I (g8925));
INVX1 gate5857(.O (g12892), .I (g8928));
INVX1 gate5858(.O (g12894), .I (g8934));
INVX1 gate5859(.O (I19952), .I (g8571));
INVX1 gate5860(.O (g12895), .I (I19952));
INVX1 gate5861(.O (g12900), .I (g8941));
INVX1 gate5862(.O (I19958), .I (g8574));
INVX1 gate5863(.O (g12901), .I (I19958));
INVX1 gate5864(.O (I19961), .I (g10747));
INVX1 gate5865(.O (g12904), .I (I19961));
INVX1 gate5866(.O (g12907), .I (g8949));
INVX1 gate5867(.O (g12909), .I (g10904));
INVX1 gate5868(.O (g12914), .I (g8952));
INVX1 gate5869(.O (g12915), .I (g8955));
INVX1 gate5870(.O (g12921), .I (g8958));
INVX1 gate5871(.O (g12922), .I (g8961));
INVX1 gate5872(.O (g12931), .I (g8965));
INVX1 gate5873(.O (g12932), .I (g8968));
INVX1 gate5874(.O (g12934), .I (g8974));
INVX1 gate5875(.O (I19986), .I (g8577));
INVX1 gate5876(.O (g12935), .I (I19986));
INVX1 gate5877(.O (g12940), .I (g8980));
INVX1 gate5878(.O (g12943), .I (g8984));
INVX1 gate5879(.O (g12944), .I (g8987));
INVX1 gate5880(.O (g12950), .I (g8990));
INVX1 gate5881(.O (g12951), .I (g8993));
INVX1 gate5882(.O (g12960), .I (g8997));
INVX1 gate5883(.O (g12961), .I (g9000));
INVX1 gate5884(.O (I20009), .I (g8313));
INVX1 gate5885(.O (g12962), .I (I20009));
INVX1 gate5886(.O (g12965), .I (g9006));
INVX1 gate5887(.O (g12969), .I (g9010));
INVX1 gate5888(.O (g12972), .I (g9013));
INVX1 gate5889(.O (g12973), .I (g9016));
INVX1 gate5890(.O (g12979), .I (g9019));
INVX1 gate5891(.O (g12980), .I (g9022));
INVX1 gate5892(.O (g12993), .I (g9035));
INVX1 gate5893(.O (g12996), .I (g9038));
INVX1 gate5894(.O (g12997), .I (g9041));
INVX1 gate5895(.O (g12998), .I (g9044));
INVX1 gate5896(.O (g13003), .I (g9058));
INVX1 gate5897(.O (I20062), .I (g10480));
INVX1 gate5898(.O (g13011), .I (I20062));
INVX1 gate5899(.O (g13025), .I (g10810));
INVX1 gate5900(.O (g13033), .I (g10797));
INVX1 gate5901(.O (g13036), .I (g10831));
INVX1 gate5902(.O (g13043), .I (g10789));
INVX1 gate5903(.O (g13046), .I (g10814));
INVX1 gate5904(.O (g13049), .I (g10851));
INVX1 gate5905(.O (g13057), .I (g10784));
INVX1 gate5906(.O (g13060), .I (g10801));
INVX1 gate5907(.O (g13063), .I (g10835));
INVX1 gate5908(.O (g13066), .I (g10872));
INVX1 gate5909(.O (I20117), .I (g10876));
INVX1 gate5910(.O (g13070), .I (I20117));
INVX1 gate5911(.O (g13073), .I (g10793));
INVX1 gate5912(.O (g13076), .I (g10818));
INVX1 gate5913(.O (g13079), .I (g10855));
INVX1 gate5914(.O (g13092), .I (g10805));
INVX1 gate5915(.O (g13095), .I (g10839));
INVX1 gate5916(.O (g13101), .I (g9128));
INVX1 gate5917(.O (g13107), .I (g10822));
INVX1 gate5918(.O (g13117), .I (g9134));
INVX1 gate5919(.O (g13130), .I (g9140));
INVX1 gate5920(.O (g13141), .I (g9146));
INVX1 gate5921(.O (g13148), .I (g9170));
INVX1 gate5922(.O (g13151), .I (g9184));
INVX1 gate5923(.O (g13152), .I (g9196));
INVX1 gate5924(.O (g13153), .I (g9199));
INVX1 gate5925(.O (g13154), .I (g9212));
INVX1 gate5926(.O (g13157), .I (g9229));
INVX1 gate5927(.O (g13158), .I (g9242));
INVX1 gate5928(.O (g13159), .I (g9245));
INVX1 gate5929(.O (g13161), .I (g9257));
INVX1 gate5930(.O (g13162), .I (g9260));
INVX1 gate5931(.O (g13163), .I (g9273));
INVX1 gate5932(.O (g13166), .I (g9290));
INVX1 gate5933(.O (g13167), .I (g9303));
INVX1 gate5934(.O (g13168), .I (g9306));
INVX1 gate5935(.O (g13169), .I (g9320));
INVX1 gate5936(.O (g13170), .I (g9323));
INVX1 gate5937(.O (g13172), .I (g9335));
INVX1 gate5938(.O (g13173), .I (g9338));
INVX1 gate5939(.O (g13174), .I (g9351));
INVX1 gate5940(.O (g13176), .I (g9368));
INVX1 gate5941(.O (g13177), .I (g9371));
INVX1 gate5942(.O (g13178), .I (g9384));
INVX1 gate5943(.O (g13179), .I (g9387));
INVX1 gate5944(.O (g13180), .I (g9401));
INVX1 gate5945(.O (g13181), .I (g9404));
INVX1 gate5946(.O (g13183), .I (g9416));
INVX1 gate5947(.O (g13184), .I (g9419));
INVX1 gate5948(.O (g13185), .I (g9443));
INVX1 gate5949(.O (g13186), .I (g9446));
INVX1 gate5950(.O (g13187), .I (g9450));
INVX1 gate5951(.O (g13188), .I (g9465));
INVX1 gate5952(.O (g13189), .I (g9468));
INVX1 gate5953(.O (g13190), .I (g9481));
INVX1 gate5954(.O (g13191), .I (g9484));
INVX1 gate5955(.O (g13192), .I (g9498));
INVX1 gate5956(.O (g13193), .I (g9501));
INVX1 gate5957(.O (g13195), .I (g9524));
INVX1 gate5958(.O (g13196), .I (g9528));
INVX1 gate5959(.O (g13197), .I (g9531));
INVX1 gate5960(.O (g13198), .I (g9585));
INVX1 gate5961(.O (g13199), .I (g9588));
INVX1 gate5962(.O (g13200), .I (g9592));
INVX1 gate5963(.O (g13201), .I (g9607));
INVX1 gate5964(.O (g13202), .I (g9610));
INVX1 gate5965(.O (g13203), .I (g9623));
INVX1 gate5966(.O (g13204), .I (g9626));
INVX1 gate5967(.O (g13205), .I (g9641));
INVX1 gate5968(.O (g13206), .I (g9644));
INVX1 gate5969(.O (g13207), .I (g9666));
INVX1 gate5970(.O (g13208), .I (g9670));
INVX1 gate5971(.O (g13209), .I (g9673));
INVX1 gate5972(.O (g13210), .I (g9727));
INVX1 gate5973(.O (g13211), .I (g9730));
INVX1 gate5974(.O (g13212), .I (g9734));
INVX1 gate5975(.O (g13213), .I (g9749));
INVX1 gate5976(.O (g13214), .I (g9752));
INVX1 gate5977(.O (I20264), .I (g9027));
INVX1 gate5978(.O (g13215), .I (I20264));
INVX1 gate5979(.O (g13218), .I (g9767));
INVX1 gate5980(.O (g13219), .I (g9770));
INVX1 gate5981(.O (g13220), .I (g9787));
INVX1 gate5982(.O (g13221), .I (g9790));
INVX1 gate5983(.O (g13222), .I (g9812));
INVX1 gate5984(.O (g13223), .I (g9816));
INVX1 gate5985(.O (g13224), .I (g9819));
INVX1 gate5986(.O (g13225), .I (g9873));
INVX1 gate5987(.O (g13226), .I (g9876));
INVX1 gate5988(.O (g13227), .I (g9880));
INVX1 gate5989(.O (I20278), .I (g9027));
INVX1 gate5990(.O (g13229), .I (I20278));
INVX1 gate5991(.O (g13232), .I (g9895));
INVX1 gate5992(.O (g13233), .I (g9898));
INVX1 gate5993(.O (I20283), .I (g9050));
INVX1 gate5994(.O (g13234), .I (I20283));
INVX1 gate5995(.O (g13237), .I (g9913));
INVX1 gate5996(.O (g13238), .I (g9916));
INVX1 gate5997(.O (g13239), .I (g9933));
INVX1 gate5998(.O (g13240), .I (g9936));
INVX1 gate5999(.O (g13241), .I (g9958));
INVX1 gate6000(.O (g13242), .I (g9962));
INVX1 gate6001(.O (g13243), .I (g9965));
INVX1 gate6002(.O (g13244), .I (g10004));
INVX1 gate6003(.O (I20295), .I (g10015));
INVX1 gate6004(.O (g13246), .I (I20295));
INVX1 gate6005(.O (I20299), .I (g10800));
INVX1 gate6006(.O (g13248), .I (I20299));
INVX1 gate6007(.O (g13249), .I (g10018));
INVX1 gate6008(.O (g13250), .I (g10021));
INVX1 gate6009(.O (I20305), .I (g9050));
INVX1 gate6010(.O (g13252), .I (I20305));
INVX1 gate6011(.O (g13255), .I (g10049));
INVX1 gate6012(.O (g13256), .I (g10052));
INVX1 gate6013(.O (I20310), .I (g9067));
INVX1 gate6014(.O (g13257), .I (I20310));
INVX1 gate6015(.O (g13260), .I (g10067));
INVX1 gate6016(.O (g13261), .I (g10070));
INVX1 gate6017(.O (g13262), .I (g10087));
INVX1 gate6018(.O (g13263), .I (g10090));
INVX1 gate6019(.O (g13264), .I (g10096));
INVX1 gate6020(.O (g13265), .I (g8568));
INVX1 gate6021(.O (I20320), .I (g10792));
INVX1 gate6022(.O (g13267), .I (I20320));
INVX1 gate6023(.O (g13268), .I (g10109));
INVX1 gate6024(.O (I20324), .I (g10124));
INVX1 gate6025(.O (g13269), .I (I20324));
INVX1 gate6026(.O (I20328), .I (g10817));
INVX1 gate6027(.O (g13271), .I (I20328));
INVX1 gate6028(.O (g13272), .I (g10127));
INVX1 gate6029(.O (g13273), .I (g10130));
INVX1 gate6030(.O (I20334), .I (g9067));
INVX1 gate6031(.O (g13275), .I (I20334));
INVX1 gate6032(.O (g13278), .I (g10158));
INVX1 gate6033(.O (g13279), .I (g10161));
INVX1 gate6034(.O (I20339), .I (g9084));
INVX1 gate6035(.O (g13280), .I (I20339));
INVX1 gate6036(.O (g13283), .I (g10176));
INVX1 gate6037(.O (g13284), .I (g10179));
INVX1 gate6038(.O (g13285), .I (g10189));
INVX1 gate6039(.O (I20347), .I (g10787));
INVX1 gate6040(.O (g13290), .I (I20347));
INVX1 gate6041(.O (I20351), .I (g10804));
INVX1 gate6042(.O (g13292), .I (I20351));
INVX1 gate6043(.O (g13293), .I (g10214));
INVX1 gate6044(.O (I20355), .I (g10229));
INVX1 gate6045(.O (g13294), .I (I20355));
INVX1 gate6046(.O (I20359), .I (g10838));
INVX1 gate6047(.O (g13296), .I (I20359));
INVX1 gate6048(.O (g13297), .I (g10232));
INVX1 gate6049(.O (g13298), .I (g10235));
INVX1 gate6050(.O (I20365), .I (g9084));
INVX1 gate6051(.O (g13300), .I (I20365));
INVX1 gate6052(.O (g13303), .I (g10263));
INVX1 gate6053(.O (g13304), .I (g10266));
INVX1 gate6054(.O (g13308), .I (g10273));
INVX1 gate6055(.O (g13309), .I (g10276));
INVX1 gate6056(.O (I20376), .I (g8569));
INVX1 gate6057(.O (g13317), .I (I20376));
INVX1 gate6058(.O (I20379), .I (g11213));
INVX1 gate6059(.O (g13318), .I (I20379));
INVX1 gate6060(.O (I20382), .I (g10907));
INVX1 gate6061(.O (g13319), .I (I20382));
INVX1 gate6062(.O (I20386), .I (g10796));
INVX1 gate6063(.O (g13321), .I (I20386));
INVX1 gate6064(.O (I20390), .I (g10821));
INVX1 gate6065(.O (g13323), .I (I20390));
INVX1 gate6066(.O (g13324), .I (g10316));
INVX1 gate6067(.O (I20394), .I (g10331));
INVX1 gate6068(.O (g13325), .I (I20394));
INVX1 gate6069(.O (I20398), .I (g10858));
INVX1 gate6070(.O (g13327), .I (I20398));
INVX1 gate6071(.O (g13328), .I (g10334));
INVX1 gate6072(.O (g13329), .I (g10337));
INVX1 gate6073(.O (g13330), .I (g10357));
INVX1 gate6074(.O (I20407), .I (g9027));
INVX1 gate6075(.O (g13336), .I (I20407));
INVX1 gate6076(.O (I20410), .I (g10887));
INVX1 gate6077(.O (g13339), .I (I20410));
INVX1 gate6078(.O (I20414), .I (g8575));
INVX1 gate6079(.O (g13341), .I (I20414));
INVX1 gate6080(.O (I20417), .I (g10933));
INVX1 gate6081(.O (g13342), .I (I20417));
INVX1 gate6082(.O (I20421), .I (g10808));
INVX1 gate6083(.O (g13344), .I (I20421));
INVX1 gate6084(.O (I20425), .I (g10842));
INVX1 gate6085(.O (g13346), .I (I20425));
INVX1 gate6086(.O (g13347), .I (g10409));
INVX1 gate6087(.O (g13351), .I (g10416));
INVX1 gate6088(.O (g13352), .I (g10419));
INVX1 gate6089(.O (I20441), .I (g9027));
INVX1 gate6090(.O (g13356), .I (I20441));
INVX1 gate6091(.O (I20444), .I (g10869));
INVX1 gate6092(.O (g13359), .I (I20444));
INVX1 gate6093(.O (I20448), .I (g9050));
INVX1 gate6094(.O (g13361), .I (I20448));
INVX1 gate6095(.O (I20451), .I (g10908));
INVX1 gate6096(.O (g13364), .I (I20451));
INVX1 gate6097(.O (I20455), .I (g8578));
INVX1 gate6098(.O (g13366), .I (I20455));
INVX1 gate6099(.O (I20458), .I (g10972));
INVX1 gate6100(.O (g13367), .I (I20458));
INVX1 gate6101(.O (I20462), .I (g10825));
INVX1 gate6102(.O (g13369), .I (I20462));
INVX1 gate6103(.O (g13373), .I (g10482));
INVX1 gate6104(.O (I20476), .I (g9027));
INVX1 gate6105(.O (g13381), .I (I20476));
INVX1 gate6106(.O (I20479), .I (g10849));
INVX1 gate6107(.O (g13384), .I (I20479));
INVX1 gate6108(.O (I20483), .I (g9050));
INVX1 gate6109(.O (g13386), .I (I20483));
INVX1 gate6110(.O (I20486), .I (g10889));
INVX1 gate6111(.O (g13389), .I (I20486));
INVX1 gate6112(.O (I20490), .I (g9067));
INVX1 gate6113(.O (g13391), .I (I20490));
INVX1 gate6114(.O (I20493), .I (g10934));
INVX1 gate6115(.O (g13394), .I (I20493));
INVX1 gate6116(.O (I20497), .I (g8579));
INVX1 gate6117(.O (g13396), .I (I20497));
INVX1 gate6118(.O (I20500), .I (g11007));
INVX1 gate6119(.O (g13397), .I (I20500));
INVX1 gate6120(.O (g13398), .I (g10542));
INVX1 gate6121(.O (g13400), .I (g10545));
INVX1 gate6122(.O (I20514), .I (g11769));
INVX1 gate6123(.O (g13405), .I (I20514));
INVX1 gate6124(.O (I20517), .I (g12425));
INVX1 gate6125(.O (g13406), .I (I20517));
INVX1 gate6126(.O (I20520), .I (g13246));
INVX1 gate6127(.O (g13407), .I (I20520));
INVX1 gate6128(.O (I20523), .I (g13317));
INVX1 gate6129(.O (g13408), .I (I20523));
INVX1 gate6130(.O (I20526), .I (g12519));
INVX1 gate6131(.O (g13409), .I (I20526));
INVX1 gate6132(.O (I20529), .I (g13319));
INVX1 gate6133(.O (g13410), .I (I20529));
INVX1 gate6134(.O (I20532), .I (g13339));
INVX1 gate6135(.O (g13411), .I (I20532));
INVX1 gate6136(.O (I20535), .I (g13359));
INVX1 gate6137(.O (g13412), .I (I20535));
INVX1 gate6138(.O (I20538), .I (g13384));
INVX1 gate6139(.O (g13413), .I (I20538));
INVX1 gate6140(.O (I20541), .I (g11599));
INVX1 gate6141(.O (g13414), .I (I20541));
INVX1 gate6142(.O (I20544), .I (g11628));
INVX1 gate6143(.O (g13415), .I (I20544));
INVX1 gate6144(.O (I20547), .I (g13248));
INVX1 gate6145(.O (g13416), .I (I20547));
INVX1 gate6146(.O (I20550), .I (g13267));
INVX1 gate6147(.O (g13417), .I (I20550));
INVX1 gate6148(.O (I20553), .I (g13290));
INVX1 gate6149(.O (g13418), .I (I20553));
INVX1 gate6150(.O (I20556), .I (g12435));
INVX1 gate6151(.O (g13419), .I (I20556));
INVX1 gate6152(.O (I20559), .I (g11937));
INVX1 gate6153(.O (g13420), .I (I20559));
INVX1 gate6154(.O (I20562), .I (g11786));
INVX1 gate6155(.O (g13421), .I (I20562));
INVX1 gate6156(.O (I20565), .I (g12432));
INVX1 gate6157(.O (g13422), .I (I20565));
INVX1 gate6158(.O (I20568), .I (g13269));
INVX1 gate6159(.O (g13423), .I (I20568));
INVX1 gate6160(.O (I20571), .I (g13341));
INVX1 gate6161(.O (g13424), .I (I20571));
INVX1 gate6162(.O (I20574), .I (g12534));
INVX1 gate6163(.O (g13425), .I (I20574));
INVX1 gate6164(.O (I20577), .I (g13342));
INVX1 gate6165(.O (g13426), .I (I20577));
INVX1 gate6166(.O (I20580), .I (g13364));
INVX1 gate6167(.O (g13427), .I (I20580));
INVX1 gate6168(.O (I20583), .I (g13389));
INVX1 gate6169(.O (g13428), .I (I20583));
INVX1 gate6170(.O (I20586), .I (g11606));
INVX1 gate6171(.O (g13429), .I (I20586));
INVX1 gate6172(.O (I20589), .I (g11629));
INVX1 gate6173(.O (g13430), .I (I20589));
INVX1 gate6174(.O (I20592), .I (g11651));
INVX1 gate6175(.O (g13431), .I (I20592));
INVX1 gate6176(.O (I20595), .I (g13271));
INVX1 gate6177(.O (g13432), .I (I20595));
INVX1 gate6178(.O (I20598), .I (g13292));
INVX1 gate6179(.O (g13433), .I (I20598));
INVX1 gate6180(.O (I20601), .I (g13321));
INVX1 gate6181(.O (g13434), .I (I20601));
INVX1 gate6182(.O (I20604), .I (g12440));
INVX1 gate6183(.O (g13435), .I (I20604));
INVX1 gate6184(.O (I20607), .I (g11990));
INVX1 gate6185(.O (g13436), .I (I20607));
INVX1 gate6186(.O (I20610), .I (g11812));
INVX1 gate6187(.O (g13437), .I (I20610));
INVX1 gate6188(.O (I20613), .I (g12437));
INVX1 gate6189(.O (g13438), .I (I20613));
INVX1 gate6190(.O (I20616), .I (g13294));
INVX1 gate6191(.O (g13439), .I (I20616));
INVX1 gate6192(.O (I20619), .I (g13366));
INVX1 gate6193(.O (g13440), .I (I20619));
INVX1 gate6194(.O (I20622), .I (g12543));
INVX1 gate6195(.O (g13441), .I (I20622));
INVX1 gate6196(.O (I20625), .I (g13367));
INVX1 gate6197(.O (g13442), .I (I20625));
INVX1 gate6198(.O (I20628), .I (g13394));
INVX1 gate6199(.O (g13443), .I (I20628));
INVX1 gate6200(.O (I20631), .I (g11611));
INVX1 gate6201(.O (g13444), .I (I20631));
INVX1 gate6202(.O (I20634), .I (g11636));
INVX1 gate6203(.O (g13445), .I (I20634));
INVX1 gate6204(.O (I20637), .I (g11652));
INVX1 gate6205(.O (g13446), .I (I20637));
INVX1 gate6206(.O (I20640), .I (g11670));
INVX1 gate6207(.O (g13447), .I (I20640));
INVX1 gate6208(.O (I20643), .I (g13296));
INVX1 gate6209(.O (g13448), .I (I20643));
INVX1 gate6210(.O (I20646), .I (g13323));
INVX1 gate6211(.O (g13449), .I (I20646));
INVX1 gate6212(.O (I20649), .I (g13344));
INVX1 gate6213(.O (g13450), .I (I20649));
INVX1 gate6214(.O (I20652), .I (g12445));
INVX1 gate6215(.O (g13451), .I (I20652));
INVX1 gate6216(.O (I20655), .I (g12059));
INVX1 gate6217(.O (g13452), .I (I20655));
INVX1 gate6218(.O (I20658), .I (g11845));
INVX1 gate6219(.O (g13453), .I (I20658));
INVX1 gate6220(.O (I20661), .I (g12442));
INVX1 gate6221(.O (g13454), .I (I20661));
INVX1 gate6222(.O (I20664), .I (g13325));
INVX1 gate6223(.O (g13455), .I (I20664));
INVX1 gate6224(.O (I20667), .I (g13396));
INVX1 gate6225(.O (g13456), .I (I20667));
INVX1 gate6226(.O (I20670), .I (g12552));
INVX1 gate6227(.O (g13457), .I (I20670));
INVX1 gate6228(.O (I20673), .I (g13397));
INVX1 gate6229(.O (g13458), .I (I20673));
INVX1 gate6230(.O (I20676), .I (g11616));
INVX1 gate6231(.O (g13459), .I (I20676));
INVX1 gate6232(.O (I20679), .I (g11641));
INVX1 gate6233(.O (g13460), .I (I20679));
INVX1 gate6234(.O (I20682), .I (g11659));
INVX1 gate6235(.O (g13461), .I (I20682));
INVX1 gate6236(.O (I20685), .I (g11671));
INVX1 gate6237(.O (g13462), .I (I20685));
INVX1 gate6238(.O (I20688), .I (g11682));
INVX1 gate6239(.O (g13463), .I (I20688));
INVX1 gate6240(.O (I20691), .I (g13327));
INVX1 gate6241(.O (g13464), .I (I20691));
INVX1 gate6242(.O (I20694), .I (g13346));
INVX1 gate6243(.O (g13465), .I (I20694));
INVX1 gate6244(.O (I20697), .I (g13369));
INVX1 gate6245(.O (g13466), .I (I20697));
INVX1 gate6246(.O (I20700), .I (g12450));
INVX1 gate6247(.O (g13467), .I (I20700));
INVX1 gate6248(.O (I20703), .I (g12123));
INVX1 gate6249(.O (g13468), .I (I20703));
INVX1 gate6250(.O (I20706), .I (g11490));
INVX1 gate6251(.O (g13469), .I (I20706));
INVX1 gate6252(.O (I20709), .I (g13070));
INVX1 gate6253(.O (g13475), .I (I20709));
INVX1 gate6254(.O (g13519), .I (g13228));
INVX1 gate6255(.O (g13530), .I (g13251));
INVX1 gate6256(.O (g13541), .I (g13274));
INVX1 gate6257(.O (g13552), .I (g13299));
INVX1 gate6258(.O (g13565), .I (g12192));
INVX1 gate6259(.O (g13568), .I (g11627));
INVX1 gate6260(.O (I20791), .I (g13149));
INVX1 gate6261(.O (g13571), .I (I20791));
INVX1 gate6262(.O (I20794), .I (g13111));
INVX1 gate6263(.O (g13572), .I (I20794));
INVX1 gate6264(.O (g13573), .I (g12247));
INVX1 gate6265(.O (g13576), .I (g11650));
INVX1 gate6266(.O (I20799), .I (g13155));
INVX1 gate6267(.O (g13579), .I (I20799));
INVX1 gate6268(.O (I20802), .I (g13160));
INVX1 gate6269(.O (g13580), .I (I20802));
INVX1 gate6270(.O (I20805), .I (g13124));
INVX1 gate6271(.O (g13581), .I (I20805));
INVX1 gate6272(.O (g13582), .I (g12290));
INVX1 gate6273(.O (g13585), .I (g11669));
INVX1 gate6274(.O (I20810), .I (g13164));
INVX1 gate6275(.O (g13588), .I (I20810));
INVX1 gate6276(.O (I20813), .I (g13265));
INVX1 gate6277(.O (g13589), .I (I20813));
INVX1 gate6278(.O (I20816), .I (g12487));
INVX1 gate6279(.O (g13598), .I (I20816));
INVX1 gate6280(.O (I20820), .I (g13171));
INVX1 gate6281(.O (g13600), .I (I20820));
INVX1 gate6282(.O (I20823), .I (g13135));
INVX1 gate6283(.O (g13601), .I (I20823));
INVX1 gate6284(.O (g13602), .I (g12326));
INVX1 gate6285(.O (g13605), .I (g11681));
INVX1 gate6286(.O (I20828), .I (g13175));
INVX1 gate6287(.O (g13608), .I (I20828));
INVX1 gate6288(.O (I20832), .I (g12507));
INVX1 gate6289(.O (g13610), .I (I20832));
INVX1 gate6290(.O (I20836), .I (g13182));
INVX1 gate6291(.O (g13612), .I (I20836));
INVX1 gate6292(.O (I20839), .I (g13143));
INVX1 gate6293(.O (g13613), .I (I20839));
INVX1 gate6294(.O (g13614), .I (g11690));
INVX1 gate6295(.O (I20844), .I (g12524));
INVX1 gate6296(.O (g13620), .I (I20844));
INVX1 gate6297(.O (I20848), .I (g13194));
INVX1 gate6298(.O (g13622), .I (I20848));
INVX1 gate6299(.O (I20852), .I (g12457));
INVX1 gate6300(.O (g13624), .I (I20852));
INVX1 gate6301(.O (g13626), .I (g11697));
INVX1 gate6302(.O (I20858), .I (g12539));
INVX1 gate6303(.O (g13632), .I (I20858));
INVX1 gate6304(.O (I20863), .I (g12467));
INVX1 gate6305(.O (g13635), .I (I20863));
INVX1 gate6306(.O (g13637), .I (g11703));
INVX1 gate6307(.O (g13644), .I (g13215));
INVX1 gate6308(.O (I20873), .I (g12482));
INVX1 gate6309(.O (g13647), .I (I20873));
INVX1 gate6310(.O (g13649), .I (g11711));
INVX1 gate6311(.O (g13657), .I (g12452));
INVX1 gate6312(.O (g13669), .I (g13229));
INVX1 gate6313(.O (g13670), .I (g13234));
INVX1 gate6314(.O (I20886), .I (g12499));
INVX1 gate6315(.O (g13673), .I (I20886));
INVX1 gate6316(.O (g13677), .I (g12447));
INVX1 gate6317(.O (g13687), .I (g12460));
INVX1 gate6318(.O (g13699), .I (g13252));
INVX1 gate6319(.O (g13700), .I (g13257));
INVX1 gate6320(.O (g13706), .I (g12443));
INVX1 gate6321(.O (g13714), .I (g12453));
INVX1 gate6322(.O (g13724), .I (g12470));
INVX1 gate6323(.O (g13736), .I (g13275));
INVX1 gate6324(.O (g13737), .I (g13280));
INVX1 gate6325(.O (I20909), .I (g13055));
INVX1 gate6326(.O (g13741), .I (I20909));
INVX1 gate6327(.O (g13750), .I (g12439));
INVX1 gate6328(.O (g13756), .I (g12448));
INVX1 gate6329(.O (g13764), .I (g12461));
INVX1 gate6330(.O (g13774), .I (g12485));
INVX1 gate6331(.O (g13786), .I (g13300));
INVX1 gate6332(.O (g13791), .I (g12444));
INVX1 gate6333(.O (g13797), .I (g12454));
INVX1 gate6334(.O (g13805), .I (g12471));
INVX1 gate6335(.O (g13817), .I (g13336));
INVX1 gate6336(.O (g13819), .I (g12449));
INVX1 gate6337(.O (g13825), .I (g12462));
INVX1 gate6338(.O (g13836), .I (g13356));
INVX1 gate6339(.O (g13838), .I (g13361));
INVX1 gate6340(.O (g13840), .I (g12455));
INVX1 gate6341(.O (g13848), .I (g11744));
INVX1 gate6342(.O (g13849), .I (g13381));
INVX1 gate6343(.O (g13850), .I (g13386));
INVX1 gate6344(.O (g13852), .I (g13391));
INVX1 gate6345(.O (g13856), .I (g11759));
INVX1 gate6346(.O (g13857), .I (g11760));
INVX1 gate6347(.O (g13858), .I (g11603));
INVX1 gate6348(.O (g13859), .I (g11608));
INVX1 gate6349(.O (g13861), .I (g11613));
INVX1 gate6350(.O (I20959), .I (g11713));
INVX1 gate6351(.O (g13863), .I (I20959));
INVX1 gate6352(.O (g13864), .I (g11767));
INVX1 gate6353(.O (g13866), .I (g11772));
INVX1 gate6354(.O (g13867), .I (g11773));
INVX1 gate6355(.O (g13868), .I (g11633));
INVX1 gate6356(.O (g13869), .I (g11638));
INVX1 gate6357(.O (g13872), .I (g11780));
INVX1 gate6358(.O (g13873), .I (g12698));
INVX1 gate6359(.O (g13879), .I (g11784));
INVX1 gate6360(.O (g13881), .I (g11789));
INVX1 gate6361(.O (g13882), .I (g11790));
INVX1 gate6362(.O (g13883), .I (g11656));
INVX1 gate6363(.O (g13885), .I (g11799));
INVX1 gate6364(.O (g13886), .I (g12747));
INVX1 gate6365(.O (g13894), .I (g11806));
INVX1 gate6366(.O (g13895), .I (g12755));
INVX1 gate6367(.O (g13901), .I (g11810));
INVX1 gate6368(.O (g13903), .I (g11815));
INVX1 gate6369(.O (g13906), .I (g11822));
INVX1 gate6370(.O (g13907), .I (g12781));
INVX1 gate6371(.O (g13918), .I (g11830));
INVX1 gate6372(.O (g13922), .I (g11831));
INVX1 gate6373(.O (g13926), .I (g11832));
INVX1 gate6374(.O (g13927), .I (g12789));
INVX1 gate6375(.O (g13935), .I (g11839));
INVX1 gate6376(.O (g13936), .I (g12797));
INVX1 gate6377(.O (g13942), .I (g11843));
INVX1 gate6378(.O (g13945), .I (g11855));
INVX1 gate6379(.O (g13946), .I (g12814));
INVX1 gate6380(.O (I21012), .I (g12503));
INVX1 gate6381(.O (g13954), .I (I21012));
INVX1 gate6382(.O (g13958), .I (g11863));
INVX1 gate6383(.O (g13962), .I (g11864));
INVX1 gate6384(.O (g13963), .I (g12820));
INVX1 gate6385(.O (g13974), .I (g11872));
INVX1 gate6386(.O (g13978), .I (g11873));
INVX1 gate6387(.O (g13982), .I (g11874));
INVX1 gate6388(.O (g13983), .I (g12828));
INVX1 gate6389(.O (g13991), .I (g11881));
INVX1 gate6390(.O (g13992), .I (g12836));
INVX1 gate6391(.O (g13999), .I (g11889));
INVX1 gate6392(.O (g14000), .I (g11890));
INVX1 gate6393(.O (g14001), .I (g12849));
INVX1 gate6394(.O (I21037), .I (g12486));
INVX1 gate6395(.O (g14008), .I (I21037));
INVX1 gate6396(.O (g14011), .I (g11896));
INVX1 gate6397(.O (g14015), .I (g11897));
INVX1 gate6398(.O (g14016), .I (g12852));
INVX1 gate6399(.O (I21045), .I (g12520));
INVX1 gate6400(.O (g14024), .I (I21045));
INVX1 gate6401(.O (g14028), .I (g11905));
INVX1 gate6402(.O (g14032), .I (g11906));
INVX1 gate6403(.O (g14033), .I (g12858));
INVX1 gate6404(.O (g14044), .I (g11914));
INVX1 gate6405(.O (g14048), .I (g11915));
INVX1 gate6406(.O (g14052), .I (g11916));
INVX1 gate6407(.O (g14053), .I (g12866));
INVX1 gate6408(.O (g14061), .I (g11928));
INVX1 gate6409(.O (g14062), .I (g12880));
INVX1 gate6410(.O (I21064), .I (g13147));
INVX1 gate6411(.O (g14068), .I (I21064));
INVX1 gate6412(.O (g14071), .I (g11934));
INVX1 gate6413(.O (g14079), .I (g11935));
INVX1 gate6414(.O (g14086), .I (g11938));
INVX1 gate6415(.O (g14090), .I (g11939));
INVX1 gate6416(.O (g14091), .I (g11940));
INVX1 gate6417(.O (g14092), .I (g12890));
INVX1 gate6418(.O (I21075), .I (g12506));
INVX1 gate6419(.O (g14099), .I (I21075));
INVX1 gate6420(.O (g14102), .I (g11946));
INVX1 gate6421(.O (g14106), .I (g11947));
INVX1 gate6422(.O (g14107), .I (g12893));
INVX1 gate6423(.O (I21083), .I (g12535));
INVX1 gate6424(.O (g14115), .I (I21083));
INVX1 gate6425(.O (g14119), .I (g11955));
INVX1 gate6426(.O (g14123), .I (g11956));
INVX1 gate6427(.O (g14124), .I (g12899));
INVX1 gate6428(.O (g14135), .I (g11964));
INVX1 gate6429(.O (g14139), .I (g11965));
INVX1 gate6430(.O (I21096), .I (g11749));
INVX1 gate6431(.O (g14144), .I (I21096));
INVX1 gate6432(.O (g14148), .I (g12912));
INVX1 gate6433(.O (g14153), .I (g12913));
INVX1 gate6434(.O (g14158), .I (g11974));
INVX1 gate6435(.O (g14165), .I (g11975));
INVX1 gate6436(.O (g14171), .I (g11979));
INVX1 gate6437(.O (g14175), .I (g11980));
INVX1 gate6438(.O (g14176), .I (g11981));
INVX1 gate6439(.O (g14177), .I (g12920));
INVX1 gate6440(.O (I21108), .I (g13150));
INVX1 gate6441(.O (g14183), .I (I21108));
INVX1 gate6442(.O (g14186), .I (g11987));
INVX1 gate6443(.O (g14194), .I (g11988));
INVX1 gate6444(.O (g14201), .I (g11991));
INVX1 gate6445(.O (g14205), .I (g11992));
INVX1 gate6446(.O (g14206), .I (g11993));
INVX1 gate6447(.O (g14207), .I (g12930));
INVX1 gate6448(.O (I21119), .I (g12523));
INVX1 gate6449(.O (g14214), .I (I21119));
INVX1 gate6450(.O (g14217), .I (g11999));
INVX1 gate6451(.O (g14221), .I (g12000));
INVX1 gate6452(.O (g14222), .I (g12933));
INVX1 gate6453(.O (I21127), .I (g12544));
INVX1 gate6454(.O (g14230), .I (I21127));
INVX1 gate6455(.O (g14234), .I (g12008));
INVX1 gate6456(.O (g14238), .I (g12939));
INVX1 gate6457(.O (g14244), .I (g12026));
INVX1 gate6458(.O (g14249), .I (g12034));
INVX1 gate6459(.O (g14252), .I (g12035));
INVX1 gate6460(.O (g14256), .I (g12036));
INVX1 gate6461(.O (I21137), .I (g11749));
INVX1 gate6462(.O (g14259), .I (I21137));
INVX1 gate6463(.O (g14263), .I (g12941));
INVX1 gate6464(.O (g14268), .I (g12942));
INVX1 gate6465(.O (g14273), .I (g12043));
INVX1 gate6466(.O (g14280), .I (g12044));
INVX1 gate6467(.O (g14286), .I (g12048));
INVX1 gate6468(.O (g14290), .I (g12049));
INVX1 gate6469(.O (g14291), .I (g12050));
INVX1 gate6470(.O (g14292), .I (g12949));
INVX1 gate6471(.O (I21149), .I (g13156));
INVX1 gate6472(.O (g14298), .I (I21149));
INVX1 gate6473(.O (g14301), .I (g12056));
INVX1 gate6474(.O (g14309), .I (g12057));
INVX1 gate6475(.O (g14316), .I (g12060));
INVX1 gate6476(.O (g14320), .I (g12061));
INVX1 gate6477(.O (g14321), .I (g12062));
INVX1 gate6478(.O (g14322), .I (g12959));
INVX1 gate6479(.O (I21160), .I (g12538));
INVX1 gate6480(.O (g14329), .I (I21160));
INVX1 gate6481(.O (g14332), .I (g12068));
INVX1 gate6482(.O (I21165), .I (g13110));
INVX1 gate6483(.O (g14337), .I (I21165));
INVX1 gate6484(.O (g14342), .I (g12967));
INVX1 gate6485(.O (g14347), .I (g12079));
INVX1 gate6486(.O (g14352), .I (g12081));
INVX1 gate6487(.O (g14355), .I (g12082));
INVX1 gate6488(.O (g14359), .I (g12083));
INVX1 gate6489(.O (g14360), .I (g12968));
INVX1 gate6490(.O (g14366), .I (g12090));
INVX1 gate6491(.O (g14371), .I (g12098));
INVX1 gate6492(.O (g14374), .I (g12099));
INVX1 gate6493(.O (g14378), .I (g12100));
INVX1 gate6494(.O (I21178), .I (g11749));
INVX1 gate6495(.O (g14381), .I (I21178));
INVX1 gate6496(.O (g14385), .I (g12970));
INVX1 gate6497(.O (g14390), .I (g12971));
INVX1 gate6498(.O (g14395), .I (g12107));
INVX1 gate6499(.O (g14402), .I (g12108));
INVX1 gate6500(.O (g14408), .I (g12112));
INVX1 gate6501(.O (g14412), .I (g12113));
INVX1 gate6502(.O (g14413), .I (g12114));
INVX1 gate6503(.O (g14414), .I (g12978));
INVX1 gate6504(.O (I21190), .I (g13165));
INVX1 gate6505(.O (g14420), .I (I21190));
INVX1 gate6506(.O (g14423), .I (g12120));
INVX1 gate6507(.O (g14431), .I (g12121));
INVX1 gate6508(.O (g14438), .I (g12124));
INVX1 gate6509(.O (g14442), .I (g11768));
INVX1 gate6510(.O (g14450), .I (g12146));
INVX1 gate6511(.O (g14454), .I (g12991));
INVX1 gate6512(.O (g14459), .I (g12151));
INVX1 gate6513(.O (g14464), .I (g12153));
INVX1 gate6514(.O (g14467), .I (g12154));
INVX1 gate6515(.O (g14471), .I (g12155));
INVX1 gate6516(.O (g14472), .I (g12992));
INVX1 gate6517(.O (g14478), .I (g12162));
INVX1 gate6518(.O (g14483), .I (g12170));
INVX1 gate6519(.O (g14486), .I (g12171));
INVX1 gate6520(.O (g14490), .I (g12172));
INVX1 gate6521(.O (I21208), .I (g11749));
INVX1 gate6522(.O (g14493), .I (I21208));
INVX1 gate6523(.O (g14497), .I (g12994));
INVX1 gate6524(.O (g14502), .I (g12995));
INVX1 gate6525(.O (g14507), .I (g12179));
INVX1 gate6526(.O (g14514), .I (g12180));
INVX1 gate6527(.O (g14520), .I (g12184));
INVX1 gate6528(.O (g14524), .I (g12185));
INVX1 gate6529(.O (g14525), .I (g12195));
INVX1 gate6530(.O (g14529), .I (g11785));
INVX1 gate6531(.O (g14537), .I (g12208));
INVX1 gate6532(.O (g14541), .I (g13001));
INVX1 gate6533(.O (g14546), .I (g12213));
INVX1 gate6534(.O (g14551), .I (g12215));
INVX1 gate6535(.O (g14554), .I (g12216));
INVX1 gate6536(.O (g14558), .I (g12217));
INVX1 gate6537(.O (g14559), .I (g13002));
INVX1 gate6538(.O (g14565), .I (g12224));
INVX1 gate6539(.O (g14570), .I (g12232));
INVX1 gate6540(.O (g14573), .I (g12233));
INVX1 gate6541(.O (g14577), .I (g12234));
INVX1 gate6542(.O (g14580), .I (g12250));
INVX1 gate6543(.O (g14584), .I (g11811));
INVX1 gate6544(.O (g14592), .I (g12263));
INVX1 gate6545(.O (g14596), .I (g13022));
INVX1 gate6546(.O (g14601), .I (g12268));
INVX1 gate6547(.O (g14606), .I (g12270));
INVX1 gate6548(.O (g14609), .I (g12271));
INVX1 gate6549(.O (g14613), .I (g12272));
INVX1 gate6550(.O (g14614), .I (g12293));
INVX1 gate6551(.O (g14618), .I (g11844));
INVX1 gate6552(.O (g14626), .I (g12306));
INVX1 gate6553(.O (I21241), .I (g13378));
INVX1 gate6554(.O (g14630), .I (I21241));
INVX1 gate6555(.O (g14637), .I (g12329));
INVX1 gate6556(.O (g14641), .I (g11823));
INVX1 gate6557(.O (I21246), .I (g11624));
INVX1 gate6558(.O (g14642), .I (I21246));
INVX1 gate6559(.O (I21249), .I (g11600));
INVX1 gate6560(.O (g14650), .I (I21249));
INVX1 gate6561(.O (I21252), .I (g11644));
INVX1 gate6562(.O (g14657), .I (I21252));
INVX1 gate6563(.O (g14668), .I (g11865));
INVX1 gate6564(.O (I21256), .I (g11647));
INVX1 gate6565(.O (g14669), .I (I21256));
INVX1 gate6566(.O (I21259), .I (g11630));
INVX1 gate6567(.O (g14677), .I (I21259));
INVX1 gate6568(.O (I21262), .I (g11713));
INVX1 gate6569(.O (g14684), .I (I21262));
INVX1 gate6570(.O (g14685), .I (g12245));
INVX1 gate6571(.O (I21267), .I (g11663));
INVX1 gate6572(.O (g14691), .I (I21267));
INVX1 gate6573(.O (g14702), .I (g11907));
INVX1 gate6574(.O (I21271), .I (g11666));
INVX1 gate6575(.O (g14703), .I (I21271));
INVX1 gate6576(.O (I21274), .I (g11653));
INVX1 gate6577(.O (g14711), .I (I21274));
INVX1 gate6578(.O (I21277), .I (g12430));
INVX1 gate6579(.O (g14718), .I (I21277));
INVX1 gate6580(.O (g14719), .I (g12288));
INVX1 gate6581(.O (I21282), .I (g11675));
INVX1 gate6582(.O (g14725), .I (I21282));
INVX1 gate6583(.O (g14736), .I (g11957));
INVX1 gate6584(.O (I21286), .I (g11678));
INVX1 gate6585(.O (g14737), .I (I21286));
INVX1 gate6586(.O (I21289), .I (g12434));
INVX1 gate6587(.O (g14745), .I (I21289));
INVX1 gate6588(.O (I21292), .I (g11888));
INVX1 gate6589(.O (g14746), .I (I21292));
INVX1 gate6590(.O (g14747), .I (g12324));
INVX1 gate6591(.O (I21297), .I (g11687));
INVX1 gate6592(.O (g14753), .I (I21297));
INVX1 gate6593(.O (g14764), .I (g11791));
INVX1 gate6594(.O (I21301), .I (g12438));
INVX1 gate6595(.O (g14765), .I (I21301));
INVX1 gate6596(.O (I21304), .I (g11927));
INVX1 gate6597(.O (g14766), .I (I21304));
INVX1 gate6598(.O (g14768), .I (g12352));
INVX1 gate6599(.O (I21310), .I (g12332));
INVX1 gate6600(.O (g14774), .I (I21310));
INVX1 gate6601(.O (I21313), .I (g11743));
INVX1 gate6602(.O (g14775), .I (I21313));
INVX1 gate6603(.O (g14776), .I (g12033));
INVX1 gate6604(.O (g14794), .I (g11848));
INVX1 gate6605(.O (I21318), .I (g12362));
INVX1 gate6606(.O (g14795), .I (I21318));
INVX1 gate6607(.O (I21321), .I (g11758));
INVX1 gate6608(.O (g14796), .I (I21321));
INVX1 gate6609(.O (g14797), .I (g12080));
INVX1 gate6610(.O (g14811), .I (g12097));
INVX1 gate6611(.O (I21326), .I (g12378));
INVX1 gate6612(.O (g14829), .I (I21326));
INVX1 gate6613(.O (I21329), .I (g11766));
INVX1 gate6614(.O (g14830), .I (I21329));
INVX1 gate6615(.O (g14831), .I (g11828));
INVX1 gate6616(.O (g14837), .I (g12145));
INVX1 gate6617(.O (g14849), .I (g12152));
INVX1 gate6618(.O (g14863), .I (g12169));
INVX1 gate6619(.O (g14881), .I (g11923));
INVX1 gate6620(.O (I21337), .I (g12408));
INVX1 gate6621(.O (g14882), .I (I21337));
INVX1 gate6622(.O (I21340), .I (g11779));
INVX1 gate6623(.O (g14883), .I (I21340));
INVX1 gate6624(.O (g14885), .I (g11860));
INVX1 gate6625(.O (g14895), .I (g12193));
INVX1 gate6626(.O (g14904), .I (g11870));
INVX1 gate6627(.O (g14910), .I (g12207));
INVX1 gate6628(.O (g14922), .I (g12214));
INVX1 gate6629(.O (g14936), .I (g12231));
INVX1 gate6630(.O (I21351), .I (g12420));
INVX1 gate6631(.O (g14954), .I (I21351));
INVX1 gate6632(.O (I21354), .I (g11798));
INVX1 gate6633(.O (g14955), .I (I21354));
INVX1 gate6634(.O (g14959), .I (g11976));
INVX1 gate6635(.O (I21361), .I (g13026));
INVX1 gate6636(.O (g14960), .I (I21361));
INVX1 gate6637(.O (I21364), .I (g13028));
INVX1 gate6638(.O (g14963), .I (I21364));
INVX1 gate6639(.O (g14966), .I (g11902));
INVX1 gate6640(.O (g14976), .I (g12248));
INVX1 gate6641(.O (g14985), .I (g11912));
INVX1 gate6642(.O (g14991), .I (g12262));
INVX1 gate6643(.O (g15003), .I (g12269));
INVX1 gate6644(.O (g15017), .I (g12009));
INVX1 gate6645(.O (I21374), .I (g12424));
INVX1 gate6646(.O (g15018), .I (I21374));
INVX1 gate6647(.O (I21377), .I (g11821));
INVX1 gate6648(.O (g15019), .I (I21377));
INVX1 gate6649(.O (I21381), .I (g13157));
INVX1 gate6650(.O (g15021), .I (I21381));
INVX1 gate6651(.O (g15022), .I (g11781));
INVX1 gate6652(.O (g15032), .I (g12027));
INVX1 gate6653(.O (g15033), .I (g12030));
INVX1 gate6654(.O (I21389), .I (g12883));
INVX1 gate6655(.O (g15034), .I (I21389));
INVX1 gate6656(.O (I21392), .I (g13020));
INVX1 gate6657(.O (g15037), .I (I21392));
INVX1 gate6658(.O (I21395), .I (g13034));
INVX1 gate6659(.O (g15040), .I (I21395));
INVX1 gate6660(.O (I21398), .I (g13021));
INVX1 gate6661(.O (g15043), .I (I21398));
INVX1 gate6662(.O (g15048), .I (g12045));
INVX1 gate6663(.O (I21404), .I (g13037));
INVX1 gate6664(.O (g15049), .I (I21404));
INVX1 gate6665(.O (I21407), .I (g13039));
INVX1 gate6666(.O (g15052), .I (I21407));
INVX1 gate6667(.O (g15055), .I (g11952));
INVX1 gate6668(.O (g15065), .I (g12291));
INVX1 gate6669(.O (g15074), .I (g11962));
INVX1 gate6670(.O (g15080), .I (g12305));
INVX1 gate6671(.O (I21415), .I (g11854));
INVX1 gate6672(.O (g15092), .I (I21415));
INVX1 gate6673(.O (I21420), .I (g13166));
INVX1 gate6674(.O (g15095), .I (I21420));
INVX1 gate6675(.O (g15096), .I (g11800));
INVX1 gate6676(.O (I21426), .I (g11661));
INVX1 gate6677(.O (g15106), .I (I21426));
INVX1 gate6678(.O (I21429), .I (g13027));
INVX1 gate6679(.O (g15109), .I (I21429));
INVX1 gate6680(.O (I21432), .I (g13044));
INVX1 gate6681(.O (g15112), .I (I21432));
INVX1 gate6682(.O (I21435), .I (g11662));
INVX1 gate6683(.O (g15115), .I (I21435));
INVX1 gate6684(.O (g15118), .I (g11807));
INVX1 gate6685(.O (g15128), .I (g12091));
INVX1 gate6686(.O (g15129), .I (g12094));
INVX1 gate6687(.O (I21443), .I (g12923));
INVX1 gate6688(.O (g15130), .I (I21443));
INVX1 gate6689(.O (I21446), .I (g13029));
INVX1 gate6690(.O (g15133), .I (I21446));
INVX1 gate6691(.O (I21449), .I (g13047));
INVX1 gate6692(.O (g15136), .I (I21449));
INVX1 gate6693(.O (I21452), .I (g13030));
INVX1 gate6694(.O (g15139), .I (I21452));
INVX1 gate6695(.O (g15144), .I (g12109));
INVX1 gate6696(.O (I21458), .I (g13050));
INVX1 gate6697(.O (g15145), .I (I21458));
INVX1 gate6698(.O (I21461), .I (g13052));
INVX1 gate6699(.O (g15148), .I (I21461));
INVX1 gate6700(.O (g15151), .I (g12005));
INVX1 gate6701(.O (g15161), .I (g12327));
INVX1 gate6702(.O (g15170), .I (g12125));
INVX1 gate6703(.O (g15174), .I (g12136));
INVX1 gate6704(.O (g15175), .I (g12139));
INVX1 gate6705(.O (g15176), .I (g12142));
INVX1 gate6706(.O (g15177), .I (g12339));
INVX1 gate6707(.O (I21476), .I (g11672));
INVX1 gate6708(.O (g15179), .I (I21476));
INVX1 gate6709(.O (I21479), .I (g13035));
INVX1 gate6710(.O (g15182), .I (I21479));
INVX1 gate6711(.O (I21482), .I (g13058));
INVX1 gate6712(.O (g15185), .I (I21482));
INVX1 gate6713(.O (g15188), .I (g11833));
INVX1 gate6714(.O (I21488), .I (g11673));
INVX1 gate6715(.O (g15198), .I (I21488));
INVX1 gate6716(.O (I21491), .I (g13038));
INVX1 gate6717(.O (g15201), .I (I21491));
INVX1 gate6718(.O (I21494), .I (g13061));
INVX1 gate6719(.O (g15204), .I (I21494));
INVX1 gate6720(.O (I21497), .I (g11674));
INVX1 gate6721(.O (g15207), .I (I21497));
INVX1 gate6722(.O (g15210), .I (g11840));
INVX1 gate6723(.O (g15220), .I (g12163));
INVX1 gate6724(.O (g15221), .I (g12166));
INVX1 gate6725(.O (I21505), .I (g12952));
INVX1 gate6726(.O (g15222), .I (I21505));
INVX1 gate6727(.O (I21508), .I (g13040));
INVX1 gate6728(.O (g15225), .I (I21508));
INVX1 gate6729(.O (I21511), .I (g13064));
INVX1 gate6730(.O (g15228), .I (I21511));
INVX1 gate6731(.O (I21514), .I (g13041));
INVX1 gate6732(.O (g15231), .I (I21514));
INVX1 gate6733(.O (g15236), .I (g12181));
INVX1 gate6734(.O (I21520), .I (g13067));
INVX1 gate6735(.O (g15237), .I (I21520));
INVX1 gate6736(.O (I21523), .I (g13069));
INVX1 gate6737(.O (g15240), .I (I21523));
INVX1 gate6738(.O (I21531), .I (g11683));
INVX1 gate6739(.O (g15248), .I (I21531));
INVX1 gate6740(.O (I21534), .I (g13045));
INVX1 gate6741(.O (g15251), .I (I21534));
INVX1 gate6742(.O (I21537), .I (g13071));
INVX1 gate6743(.O (g15254), .I (I21537));
INVX1 gate6744(.O (g15260), .I (g12198));
INVX1 gate6745(.O (g15261), .I (g12201));
INVX1 gate6746(.O (g15262), .I (g12204));
INVX1 gate6747(.O (g15263), .I (g12369));
INVX1 gate6748(.O (I21548), .I (g11684));
INVX1 gate6749(.O (g15265), .I (I21548));
INVX1 gate6750(.O (I21551), .I (g13048));
INVX1 gate6751(.O (g15268), .I (I21551));
INVX1 gate6752(.O (I21554), .I (g13074));
INVX1 gate6753(.O (g15271), .I (I21554));
INVX1 gate6754(.O (g15274), .I (g11875));
INVX1 gate6755(.O (I21560), .I (g11685));
INVX1 gate6756(.O (g15284), .I (I21560));
INVX1 gate6757(.O (I21563), .I (g13051));
INVX1 gate6758(.O (g15287), .I (I21563));
INVX1 gate6759(.O (I21566), .I (g13077));
INVX1 gate6760(.O (g15290), .I (I21566));
INVX1 gate6761(.O (I21569), .I (g11686));
INVX1 gate6762(.O (g15293), .I (I21569));
INVX1 gate6763(.O (g15296), .I (g11882));
INVX1 gate6764(.O (g15306), .I (g12225));
INVX1 gate6765(.O (g15307), .I (g12228));
INVX1 gate6766(.O (I21577), .I (g12981));
INVX1 gate6767(.O (g15308), .I (I21577));
INVX1 gate6768(.O (I21580), .I (g13053));
INVX1 gate6769(.O (g15311), .I (I21580));
INVX1 gate6770(.O (I21583), .I (g13080));
INVX1 gate6771(.O (g15314), .I (I21583));
INVX1 gate6772(.O (I21586), .I (g13054));
INVX1 gate6773(.O (g15317), .I (I21586));
INVX1 gate6774(.O (g15322), .I (g12239));
INVX1 gate6775(.O (g15323), .I (g12242));
INVX1 gate6776(.O (I21595), .I (g11691));
INVX1 gate6777(.O (g15326), .I (I21595));
INVX1 gate6778(.O (I21598), .I (g13059));
INVX1 gate6779(.O (g15329), .I (I21598));
INVX1 gate6780(.O (I21601), .I (g13087));
INVX1 gate6781(.O (g15332), .I (I21601));
INVX1 gate6782(.O (I21609), .I (g11692));
INVX1 gate6783(.O (g15340), .I (I21609));
INVX1 gate6784(.O (I21612), .I (g13062));
INVX1 gate6785(.O (g15343), .I (I21612));
INVX1 gate6786(.O (I21615), .I (g13090));
INVX1 gate6787(.O (g15346), .I (I21615));
INVX1 gate6788(.O (g15352), .I (g12253));
INVX1 gate6789(.O (g15353), .I (g12256));
INVX1 gate6790(.O (g15354), .I (g12259));
INVX1 gate6791(.O (g15355), .I (g12388));
INVX1 gate6792(.O (I21626), .I (g11693));
INVX1 gate6793(.O (g15357), .I (I21626));
INVX1 gate6794(.O (I21629), .I (g13065));
INVX1 gate6795(.O (g15360), .I (I21629));
INVX1 gate6796(.O (I21632), .I (g13093));
INVX1 gate6797(.O (g15363), .I (I21632));
INVX1 gate6798(.O (g15366), .I (g11917));
INVX1 gate6799(.O (I21638), .I (g11694));
INVX1 gate6800(.O (g15376), .I (I21638));
INVX1 gate6801(.O (I21641), .I (g13068));
INVX1 gate6802(.O (g15379), .I (I21641));
INVX1 gate6803(.O (I21644), .I (g13096));
INVX1 gate6804(.O (g15382), .I (I21644));
INVX1 gate6805(.O (I21647), .I (g11695));
INVX1 gate6806(.O (g15385), .I (I21647));
INVX1 gate6807(.O (g15390), .I (g12279));
INVX1 gate6808(.O (I21655), .I (g11696));
INVX1 gate6809(.O (g15393), .I (I21655));
INVX1 gate6810(.O (I21658), .I (g13072));
INVX1 gate6811(.O (g15396), .I (I21658));
INVX1 gate6812(.O (I21661), .I (g13098));
INVX1 gate6813(.O (g15399), .I (I21661));
INVX1 gate6814(.O (I21666), .I (g13100));
INVX1 gate6815(.O (g15404), .I (I21666));
INVX1 gate6816(.O (g15408), .I (g12282));
INVX1 gate6817(.O (g15409), .I (g12285));
INVX1 gate6818(.O (I21674), .I (g11698));
INVX1 gate6819(.O (g15412), .I (I21674));
INVX1 gate6820(.O (I21677), .I (g13075));
INVX1 gate6821(.O (g15415), .I (I21677));
INVX1 gate6822(.O (I21680), .I (g13102));
INVX1 gate6823(.O (g15418), .I (I21680));
INVX1 gate6824(.O (I21688), .I (g11699));
INVX1 gate6825(.O (g15426), .I (I21688));
INVX1 gate6826(.O (I21691), .I (g13078));
INVX1 gate6827(.O (g15429), .I (I21691));
INVX1 gate6828(.O (I21694), .I (g13105));
INVX1 gate6829(.O (g15432), .I (I21694));
INVX1 gate6830(.O (g15438), .I (g12296));
INVX1 gate6831(.O (g15439), .I (g12299));
INVX1 gate6832(.O (g15440), .I (g12302));
INVX1 gate6833(.O (g15441), .I (g12418));
INVX1 gate6834(.O (I21705), .I (g11700));
INVX1 gate6835(.O (g15443), .I (I21705));
INVX1 gate6836(.O (I21708), .I (g13081));
INVX1 gate6837(.O (g15446), .I (I21708));
INVX1 gate6838(.O (I21711), .I (g13108));
INVX1 gate6839(.O (g15449), .I (I21711));
INVX1 gate6840(.O (g15458), .I (g12312));
INVX1 gate6841(.O (I21720), .I (g11701));
INVX1 gate6842(.O (g15461), .I (I21720));
INVX1 gate6843(.O (I21723), .I (g13088));
INVX1 gate6844(.O (g15464), .I (I21723));
INVX1 gate6845(.O (I21726), .I (g13112));
INVX1 gate6846(.O (g15467), .I (I21726));
INVX1 gate6847(.O (I21730), .I (g13089));
INVX1 gate6848(.O (g15471), .I (I21730));
INVX1 gate6849(.O (g15474), .I (g12315));
INVX1 gate6850(.O (I21736), .I (g11702));
INVX1 gate6851(.O (g15477), .I (I21736));
INVX1 gate6852(.O (I21739), .I (g13091));
INVX1 gate6853(.O (g15480), .I (I21739));
INVX1 gate6854(.O (I21742), .I (g13114));
INVX1 gate6855(.O (g15483), .I (I21742));
INVX1 gate6856(.O (I21747), .I (g13116));
INVX1 gate6857(.O (g15488), .I (I21747));
INVX1 gate6858(.O (g15492), .I (g12318));
INVX1 gate6859(.O (g15493), .I (g12321));
INVX1 gate6860(.O (I21755), .I (g11704));
INVX1 gate6861(.O (g15496), .I (I21755));
INVX1 gate6862(.O (I21758), .I (g13094));
INVX1 gate6863(.O (g15499), .I (I21758));
INVX1 gate6864(.O (I21761), .I (g13118));
INVX1 gate6865(.O (g15502), .I (I21761));
INVX1 gate6866(.O (I21769), .I (g11705));
INVX1 gate6867(.O (g15510), .I (I21769));
INVX1 gate6868(.O (I21772), .I (g13097));
INVX1 gate6869(.O (g15513), .I (I21772));
INVX1 gate6870(.O (I21775), .I (g13121));
INVX1 gate6871(.O (g15516), .I (I21775));
INVX1 gate6872(.O (I21780), .I (g13305));
INVX1 gate6873(.O (g15521), .I (I21780));
INVX1 gate6874(.O (g15524), .I (g12333));
INVX1 gate6875(.O (g15525), .I (g12336));
INVX1 gate6876(.O (I21787), .I (g11707));
INVX1 gate6877(.O (g15528), .I (I21787));
INVX1 gate6878(.O (I21790), .I (g13099));
INVX1 gate6879(.O (g15531), .I (I21790));
INVX1 gate6880(.O (I21793), .I (g13123));
INVX1 gate6881(.O (g15534), .I (I21793));
INVX1 gate6882(.O (I21796), .I (g11708));
INVX1 gate6883(.O (g15537), .I (I21796));
INVX1 gate6884(.O (g15544), .I (g12340));
INVX1 gate6885(.O (I21803), .I (g11709));
INVX1 gate6886(.O (g15547), .I (I21803));
INVX1 gate6887(.O (I21806), .I (g13103));
INVX1 gate6888(.O (g15550), .I (I21806));
INVX1 gate6889(.O (I21809), .I (g13125));
INVX1 gate6890(.O (g15553), .I (I21809));
INVX1 gate6891(.O (I21813), .I (g13104));
INVX1 gate6892(.O (g15557), .I (I21813));
INVX1 gate6893(.O (g15560), .I (g12343));
INVX1 gate6894(.O (I21819), .I (g11710));
INVX1 gate6895(.O (g15563), .I (I21819));
INVX1 gate6896(.O (I21822), .I (g13106));
INVX1 gate6897(.O (g15566), .I (I21822));
INVX1 gate6898(.O (I21825), .I (g13127));
INVX1 gate6899(.O (g15569), .I (I21825));
INVX1 gate6900(.O (I21830), .I (g13129));
INVX1 gate6901(.O (g15574), .I (I21830));
INVX1 gate6902(.O (g15578), .I (g12346));
INVX1 gate6903(.O (g15579), .I (g12349));
INVX1 gate6904(.O (I21838), .I (g11712));
INVX1 gate6905(.O (g15582), .I (I21838));
INVX1 gate6906(.O (I21841), .I (g13109));
INVX1 gate6907(.O (g15585), .I (I21841));
INVX1 gate6908(.O (I21844), .I (g13131));
INVX1 gate6909(.O (g15588), .I (I21844));
INVX1 gate6910(.O (I21852), .I (g11716));
INVX1 gate6911(.O (g15596), .I (I21852));
INVX1 gate6912(.O (I21855), .I (g13113));
INVX1 gate6913(.O (g15599), .I (I21855));
INVX1 gate6914(.O (g15602), .I (g12363));
INVX1 gate6915(.O (g15603), .I (g12366));
INVX1 gate6916(.O (I21862), .I (g11717));
INVX1 gate6917(.O (g15606), .I (I21862));
INVX1 gate6918(.O (I21865), .I (g13115));
INVX1 gate6919(.O (g15609), .I (I21865));
INVX1 gate6920(.O (I21868), .I (g13134));
INVX1 gate6921(.O (g15612), .I (I21868));
INVX1 gate6922(.O (I21871), .I (g11718));
INVX1 gate6923(.O (g15615), .I (I21871));
INVX1 gate6924(.O (g15622), .I (g12370));
INVX1 gate6925(.O (I21878), .I (g11719));
INVX1 gate6926(.O (g15625), .I (I21878));
INVX1 gate6927(.O (I21881), .I (g13119));
INVX1 gate6928(.O (g15628), .I (I21881));
INVX1 gate6929(.O (I21884), .I (g13136));
INVX1 gate6930(.O (g15631), .I (I21884));
INVX1 gate6931(.O (I21888), .I (g13120));
INVX1 gate6932(.O (g15635), .I (I21888));
INVX1 gate6933(.O (g15638), .I (g12373));
INVX1 gate6934(.O (I21894), .I (g11720));
INVX1 gate6935(.O (g15641), .I (I21894));
INVX1 gate6936(.O (I21897), .I (g13122));
INVX1 gate6937(.O (g15644), .I (I21897));
INVX1 gate6938(.O (I21900), .I (g13138));
INVX1 gate6939(.O (g15647), .I (I21900));
INVX1 gate6940(.O (I21905), .I (g13140));
INVX1 gate6941(.O (g15652), .I (I21905));
INVX1 gate6942(.O (I21908), .I (g13082));
INVX1 gate6943(.O (g15655), .I (I21908));
INVX1 gate6944(.O (g15659), .I (g11706));
INVX1 gate6945(.O (g15665), .I (g12379));
INVX1 gate6946(.O (I21918), .I (g11721));
INVX1 gate6947(.O (g15667), .I (I21918));
INVX1 gate6948(.O (I21923), .I (g11722));
INVX1 gate6949(.O (g15672), .I (I21923));
INVX1 gate6950(.O (I21926), .I (g13126));
INVX1 gate6951(.O (g15675), .I (I21926));
INVX1 gate6952(.O (g15678), .I (g12382));
INVX1 gate6953(.O (g15679), .I (g12385));
INVX1 gate6954(.O (I21933), .I (g11723));
INVX1 gate6955(.O (g15682), .I (I21933));
INVX1 gate6956(.O (I21936), .I (g13128));
INVX1 gate6957(.O (g15685), .I (I21936));
INVX1 gate6958(.O (I21939), .I (g13142));
INVX1 gate6959(.O (g15688), .I (I21939));
INVX1 gate6960(.O (I21942), .I (g11724));
INVX1 gate6961(.O (g15691), .I (I21942));
INVX1 gate6962(.O (g15698), .I (g12389));
INVX1 gate6963(.O (I21949), .I (g11725));
INVX1 gate6964(.O (g15701), .I (I21949));
INVX1 gate6965(.O (I21952), .I (g13132));
INVX1 gate6966(.O (g15704), .I (I21952));
INVX1 gate6967(.O (I21955), .I (g13144));
INVX1 gate6968(.O (g15707), .I (I21955));
INVX1 gate6969(.O (I21959), .I (g13133));
INVX1 gate6970(.O (g15711), .I (I21959));
INVX1 gate6971(.O (I21962), .I (g13004));
INVX1 gate6972(.O (g15714), .I (I21962));
INVX1 gate6973(.O (g15722), .I (g13011));
INVX1 gate6974(.O (g15724), .I (g12409));
INVX1 gate6975(.O (I21974), .I (g11726));
INVX1 gate6976(.O (g15726), .I (I21974));
INVX1 gate6977(.O (I21979), .I (g11727));
INVX1 gate6978(.O (g15731), .I (I21979));
INVX1 gate6979(.O (I21982), .I (g13137));
INVX1 gate6980(.O (g15734), .I (I21982));
INVX1 gate6981(.O (g15737), .I (g12412));
INVX1 gate6982(.O (g15738), .I (g12415));
INVX1 gate6983(.O (I21989), .I (g11728));
INVX1 gate6984(.O (g15741), .I (I21989));
INVX1 gate6985(.O (I21992), .I (g13139));
INVX1 gate6986(.O (g15744), .I (I21992));
INVX1 gate6987(.O (I21995), .I (g13146));
INVX1 gate6988(.O (g15747), .I (I21995));
INVX1 gate6989(.O (I21998), .I (g11729));
INVX1 gate6990(.O (g15750), .I (I21998));
INVX1 gate6991(.O (g15762), .I (g13011));
INVX1 gate6992(.O (g15764), .I (g12421));
INVX1 gate6993(.O (I22014), .I (g11730));
INVX1 gate6994(.O (g15766), .I (I22014));
INVX1 gate6995(.O (I22019), .I (g11731));
INVX1 gate6996(.O (g15771), .I (I22019));
INVX1 gate6997(.O (I22022), .I (g13145));
INVX1 gate6998(.O (g15774), .I (I22022));
INVX1 gate6999(.O (I22025), .I (g11617));
INVX1 gate7000(.O (g15777), .I (I22025));
INVX1 gate7001(.O (g15790), .I (g13011));
INVX1 gate7002(.O (g15792), .I (g12426));
INVX1 gate7003(.O (I22044), .I (g11733));
INVX1 gate7004(.O (g15794), .I (I22044));
INVX1 gate7005(.O (g15800), .I (g12909));
INVX1 gate7006(.O (g15813), .I (g13011));
INVX1 gate7007(.O (g15859), .I (g13378));
INVX1 gate7008(.O (I22120), .I (g12909));
INVX1 gate7009(.O (g15876), .I (I22120));
INVX1 gate7010(.O (g15880), .I (g11624));
INVX1 gate7011(.O (g15890), .I (g11600));
INVX1 gate7012(.O (g15904), .I (g11644));
INVX1 gate7013(.O (g15913), .I (g11647));
INVX1 gate7014(.O (g15923), .I (g11630));
INVX1 gate7015(.O (g15933), .I (g11663));
INVX1 gate7016(.O (g15942), .I (g11666));
INVX1 gate7017(.O (g15952), .I (g11653));
INVX1 gate7018(.O (g15962), .I (g11675));
INVX1 gate7019(.O (g15971), .I (g11678));
INVX1 gate7020(.O (g15981), .I (g11687));
INVX1 gate7021(.O (I22163), .I (g12433));
INVX1 gate7022(.O (g15989), .I (I22163));
INVX1 gate7023(.O (g15991), .I (g12548));
INVX1 gate7024(.O (g15994), .I (g12555));
INVX1 gate7025(.O (g15997), .I (g12561));
INVX1 gate7026(.O (g16001), .I (g12601));
INVX1 gate7027(.O (g16002), .I (g12604));
INVX1 gate7028(.O (g16005), .I (g12608));
INVX1 gate7029(.O (g16007), .I (g12647));
INVX1 gate7030(.O (g16011), .I (g12651));
INVX1 gate7031(.O (g16012), .I (g12654));
INVX1 gate7032(.O (g16013), .I (g12692));
INVX1 gate7033(.O (g16014), .I (g12695));
INVX1 gate7034(.O (g16023), .I (g12699));
INVX1 gate7035(.O (g16024), .I (g12702));
INVX1 gate7036(.O (g16025), .I (g12705));
INVX1 gate7037(.O (g16026), .I (g12708));
INVX1 gate7038(.O (g16027), .I (g12744));
INVX1 gate7039(.O (g16034), .I (g12749));
INVX1 gate7040(.O (g16035), .I (g12752));
INVX1 gate7041(.O (g16039), .I (g12756));
INVX1 gate7042(.O (g16040), .I (g12759));
INVX1 gate7043(.O (g16041), .I (g12762));
INVX1 gate7044(.O (g16042), .I (g12765));
INVX1 gate7045(.O (g16043), .I (g12769));
INVX1 gate7046(.O (g16044), .I (g12772));
INVX1 gate7047(.O (g16054), .I (g12783));
INVX1 gate7048(.O (g16055), .I (g12786));
INVX1 gate7049(.O (g16056), .I (g12791));
INVX1 gate7050(.O (g16057), .I (g12794));
INVX1 gate7051(.O (g16061), .I (g12798));
INVX1 gate7052(.O (g16062), .I (g12801));
INVX1 gate7053(.O (g16063), .I (g12804));
INVX1 gate7054(.O (g16064), .I (g12808));
INVX1 gate7055(.O (g16065), .I (g12811));
INVX1 gate7056(.O (g16075), .I (g11861));
INVX1 gate7057(.O (g16088), .I (g12816));
INVX1 gate7058(.O (g16090), .I (g12822));
INVX1 gate7059(.O (g16091), .I (g12825));
INVX1 gate7060(.O (g16092), .I (g12830));
INVX1 gate7061(.O (g16093), .I (g12833));
INVX1 gate7062(.O (g16097), .I (g12837));
INVX1 gate7063(.O (g16098), .I (g12840));
INVX1 gate7064(.O (g16099), .I (g12844));
INVX1 gate7065(.O (g16113), .I (g11903));
INVX1 gate7066(.O (g16126), .I (g12854));
INVX1 gate7067(.O (g16128), .I (g12860));
INVX1 gate7068(.O (g16129), .I (g12863));
INVX1 gate7069(.O (g16130), .I (g12868));
INVX1 gate7070(.O (g16131), .I (g12871));
INVX1 gate7071(.O (g16142), .I (g13057));
INVX1 gate7072(.O (g16154), .I (g12194));
INVX1 gate7073(.O (g16164), .I (g11953));
INVX1 gate7074(.O (g16177), .I (g12895));
INVX1 gate7075(.O (g16179), .I (g12901));
INVX1 gate7076(.O (g16180), .I (g12904));
INVX1 gate7077(.O (g16189), .I (g13043));
INVX1 gate7078(.O (g16201), .I (g13073));
INVX1 gate7079(.O (g16213), .I (g12249));
INVX1 gate7080(.O (g16223), .I (g12006));
INVX1 gate7081(.O (g16236), .I (g12935));
INVX1 gate7082(.O (g16243), .I (g13033));
INVX1 gate7083(.O (g16254), .I (g13060));
INVX1 gate7084(.O (g16266), .I (g13092));
INVX1 gate7085(.O (g16278), .I (g12292));
INVX1 gate7086(.O (g16287), .I (g12962));
INVX1 gate7087(.O (g16293), .I (g13025));
INVX1 gate7088(.O (I22382), .I (g520));
INVX1 gate7089(.O (g16297), .I (I22382));
INVX1 gate7090(.O (g16302), .I (g13046));
INVX1 gate7091(.O (g16313), .I (g13076));
INVX1 gate7092(.O (g16325), .I (g13107));
INVX1 gate7093(.O (g16337), .I (g12328));
INVX1 gate7094(.O (g16351), .I (g13036));
INVX1 gate7095(.O (I22414), .I (g1206));
INVX1 gate7096(.O (g16355), .I (I22414));
INVX1 gate7097(.O (g16360), .I (g13063));
INVX1 gate7098(.O (g16371), .I (g13095));
INVX1 gate7099(.O (g16395), .I (g13049));
INVX1 gate7100(.O (I22444), .I (g1900));
INVX1 gate7101(.O (g16399), .I (I22444));
INVX1 gate7102(.O (g16404), .I (g13079));
INVX1 gate7103(.O (g16433), .I (g13066));
INVX1 gate7104(.O (I22475), .I (g2594));
INVX1 gate7105(.O (g16437), .I (I22475));
INVX1 gate7106(.O (g16466), .I (g12017));
INVX1 gate7107(.O (I22503), .I (g13598));
INVX1 gate7108(.O (g16467), .I (I22503));
INVX1 gate7109(.O (I22506), .I (g13624));
INVX1 gate7110(.O (g16468), .I (I22506));
INVX1 gate7111(.O (I22509), .I (g13610));
INVX1 gate7112(.O (g16469), .I (I22509));
INVX1 gate7113(.O (I22512), .I (g13635));
INVX1 gate7114(.O (g16470), .I (I22512));
INVX1 gate7115(.O (I22515), .I (g13620));
INVX1 gate7116(.O (g16471), .I (I22515));
INVX1 gate7117(.O (I22518), .I (g13647));
INVX1 gate7118(.O (g16472), .I (I22518));
INVX1 gate7119(.O (I22521), .I (g13632));
INVX1 gate7120(.O (g16473), .I (I22521));
INVX1 gate7121(.O (I22524), .I (g13673));
INVX1 gate7122(.O (g16474), .I (I22524));
INVX1 gate7123(.O (I22527), .I (g13469));
INVX1 gate7124(.O (g16475), .I (I22527));
INVX1 gate7125(.O (I22530), .I (g14774));
INVX1 gate7126(.O (g16476), .I (I22530));
INVX1 gate7127(.O (I22533), .I (g14795));
INVX1 gate7128(.O (g16477), .I (I22533));
INVX1 gate7129(.O (I22536), .I (g14829));
INVX1 gate7130(.O (g16478), .I (I22536));
INVX1 gate7131(.O (I22539), .I (g14882));
INVX1 gate7132(.O (g16479), .I (I22539));
INVX1 gate7133(.O (I22542), .I (g14954));
INVX1 gate7134(.O (g16480), .I (I22542));
INVX1 gate7135(.O (I22545), .I (g15018));
INVX1 gate7136(.O (g16481), .I (I22545));
INVX1 gate7137(.O (I22548), .I (g14718));
INVX1 gate7138(.O (g16482), .I (I22548));
INVX1 gate7139(.O (I22551), .I (g14745));
INVX1 gate7140(.O (g16483), .I (I22551));
INVX1 gate7141(.O (I22554), .I (g14765));
INVX1 gate7142(.O (g16484), .I (I22554));
INVX1 gate7143(.O (I22557), .I (g14775));
INVX1 gate7144(.O (g16485), .I (I22557));
INVX1 gate7145(.O (I22560), .I (g14796));
INVX1 gate7146(.O (g16486), .I (I22560));
INVX1 gate7147(.O (I22563), .I (g14830));
INVX1 gate7148(.O (g16487), .I (I22563));
INVX1 gate7149(.O (I22566), .I (g14883));
INVX1 gate7150(.O (g16488), .I (I22566));
INVX1 gate7151(.O (I22569), .I (g14955));
INVX1 gate7152(.O (g16489), .I (I22569));
INVX1 gate7153(.O (I22572), .I (g15019));
INVX1 gate7154(.O (g16490), .I (I22572));
INVX1 gate7155(.O (I22575), .I (g15092));
INVX1 gate7156(.O (g16491), .I (I22575));
INVX1 gate7157(.O (I22578), .I (g14746));
INVX1 gate7158(.O (g16492), .I (I22578));
INVX1 gate7159(.O (I22581), .I (g14766));
INVX1 gate7160(.O (g16493), .I (I22581));
INVX1 gate7161(.O (I22584), .I (g15989));
INVX1 gate7162(.O (g16494), .I (I22584));
INVX1 gate7163(.O (I22587), .I (g14684));
INVX1 gate7164(.O (g16495), .I (I22587));
INVX1 gate7165(.O (I22590), .I (g13863));
INVX1 gate7166(.O (g16496), .I (I22590));
INVX1 gate7167(.O (I22593), .I (g15876));
INVX1 gate7168(.O (g16497), .I (I22593));
INVX1 gate7169(.O (g16501), .I (g14158));
INVX1 gate7170(.O (I22599), .I (g14966));
INVX1 gate7171(.O (g16506), .I (I22599));
INVX1 gate7172(.O (g16507), .I (g14186));
INVX1 gate7173(.O (I22604), .I (g15080));
INVX1 gate7174(.O (g16514), .I (I22604));
INVX1 gate7175(.O (g16515), .I (g14244));
INVX1 gate7176(.O (g16523), .I (g14273));
INVX1 gate7177(.O (I22611), .I (g15055));
INVX1 gate7178(.O (g16528), .I (I22611));
INVX1 gate7179(.O (g16529), .I (g14301));
INVX1 gate7180(.O (I22618), .I (g14630));
INVX1 gate7181(.O (g16540), .I (I22618));
INVX1 gate7182(.O (g16543), .I (g14347));
INVX1 gate7183(.O (g16546), .I (g14366));
INVX1 gate7184(.O (g16554), .I (g14395));
INVX1 gate7185(.O (I22626), .I (g15151));
INVX1 gate7186(.O (g16559), .I (I22626));
INVX1 gate7187(.O (g16560), .I (g14423));
INVX1 gate7188(.O (I22640), .I (g14650));
INVX1 gate7189(.O (g16572), .I (I22640));
INVX1 gate7190(.O (g16575), .I (g14459));
INVX1 gate7191(.O (g16578), .I (g14478));
INVX1 gate7192(.O (g16586), .I (g14507));
INVX1 gate7193(.O (I22651), .I (g14677));
INVX1 gate7194(.O (g16596), .I (I22651));
INVX1 gate7195(.O (g16599), .I (g14546));
INVX1 gate7196(.O (g16602), .I (g14565));
INVX1 gate7197(.O (I22657), .I (g14657));
INVX1 gate7198(.O (g16608), .I (I22657));
INVX1 gate7199(.O (I22663), .I (g14711));
INVX1 gate7200(.O (g16616), .I (I22663));
INVX1 gate7201(.O (g16619), .I (g14601));
INVX1 gate7202(.O (I22667), .I (g14642));
INVX1 gate7203(.O (g16622), .I (I22667));
INVX1 gate7204(.O (I22671), .I (g14691));
INVX1 gate7205(.O (g16626), .I (I22671));
INVX1 gate7206(.O (I22676), .I (g14630));
INVX1 gate7207(.O (g16633), .I (I22676));
INVX1 gate7208(.O (I22679), .I (g14669));
INVX1 gate7209(.O (g16636), .I (I22679));
INVX1 gate7210(.O (I22683), .I (g14725));
INVX1 gate7211(.O (g16640), .I (I22683));
INVX1 gate7212(.O (I22687), .I (g14650));
INVX1 gate7213(.O (g16644), .I (I22687));
INVX1 gate7214(.O (I22690), .I (g14703));
INVX1 gate7215(.O (g16647), .I (I22690));
INVX1 gate7216(.O (I22694), .I (g14753));
INVX1 gate7217(.O (g16651), .I (I22694));
INVX1 gate7218(.O (I22699), .I (g14677));
INVX1 gate7219(.O (g16656), .I (I22699));
INVX1 gate7220(.O (I22702), .I (g14737));
INVX1 gate7221(.O (g16659), .I (I22702));
INVX1 gate7222(.O (g16665), .I (g14776));
INVX1 gate7223(.O (I22715), .I (g14711));
INVX1 gate7224(.O (g16673), .I (I22715));
INVX1 gate7225(.O (I22718), .I (g14657));
INVX1 gate7226(.O (g16676), .I (I22718));
INVX1 gate7227(.O (g16682), .I (g14797));
INVX1 gate7228(.O (g16686), .I (g14811));
INVX1 gate7229(.O (I22726), .I (g14642));
INVX1 gate7230(.O (g16694), .I (I22726));
INVX1 gate7231(.O (g16697), .I (g14837));
INVX1 gate7232(.O (I22730), .I (g14691));
INVX1 gate7233(.O (g16702), .I (I22730));
INVX1 gate7234(.O (g16708), .I (g14849));
INVX1 gate7235(.O (g16712), .I (g14863));
INVX1 gate7236(.O (I22737), .I (g14630));
INVX1 gate7237(.O (g16719), .I (I22737));
INVX1 gate7238(.O (g16722), .I (g14895));
INVX1 gate7239(.O (I22741), .I (g14669));
INVX1 gate7240(.O (g16725), .I (I22741));
INVX1 gate7241(.O (g16728), .I (g14910));
INVX1 gate7242(.O (I22745), .I (g14725));
INVX1 gate7243(.O (g16733), .I (I22745));
INVX1 gate7244(.O (g16739), .I (g14922));
INVX1 gate7245(.O (g16743), .I (g14936));
INVX1 gate7246(.O (g16749), .I (g15782));
INVX1 gate7247(.O (I22752), .I (g14657));
INVX1 gate7248(.O (g16758), .I (I22752));
INVX1 gate7249(.O (I22755), .I (g14650));
INVX1 gate7250(.O (g16761), .I (I22755));
INVX1 gate7251(.O (g16764), .I (g14976));
INVX1 gate7252(.O (I22759), .I (g14703));
INVX1 gate7253(.O (g16767), .I (I22759));
INVX1 gate7254(.O (g16770), .I (g14991));
INVX1 gate7255(.O (I22763), .I (g14753));
INVX1 gate7256(.O (g16775), .I (I22763));
INVX1 gate7257(.O (g16781), .I (g15003));
INVX1 gate7258(.O (I22768), .I (g14691));
INVX1 gate7259(.O (g16785), .I (I22768));
INVX1 gate7260(.O (I22771), .I (g14677));
INVX1 gate7261(.O (g16788), .I (I22771));
INVX1 gate7262(.O (g16791), .I (g15065));
INVX1 gate7263(.O (I22775), .I (g14737));
INVX1 gate7264(.O (g16794), .I (I22775));
INVX1 gate7265(.O (g16797), .I (g15080));
INVX1 gate7266(.O (g16804), .I (g15803));
INVX1 gate7267(.O (g16809), .I (g15842));
INVX1 gate7268(.O (I22783), .I (g13572));
INVX1 gate7269(.O (g16813), .I (I22783));
INVX1 gate7270(.O (I22786), .I (g14725));
INVX1 gate7271(.O (g16814), .I (I22786));
INVX1 gate7272(.O (I22789), .I (g14711));
INVX1 gate7273(.O (g16817), .I (I22789));
INVX1 gate7274(.O (g16820), .I (g15161));
INVX1 gate7275(.O (g16825), .I (g15855));
INVX1 gate7276(.O (I22797), .I (g14165));
INVX1 gate7277(.O (g16830), .I (I22797));
INVX1 gate7278(.O (I22800), .I (g13581));
INVX1 gate7279(.O (g16831), .I (I22800));
INVX1 gate7280(.O (I22803), .I (g14753));
INVX1 gate7281(.O (g16832), .I (I22803));
INVX1 gate7282(.O (g16836), .I (g15818));
INVX1 gate7283(.O (g16840), .I (g15878));
INVX1 gate7284(.O (I22810), .I (g14280));
INVX1 gate7285(.O (g16842), .I (I22810));
INVX1 gate7286(.O (I22813), .I (g13601));
INVX1 gate7287(.O (g16843), .I (I22813));
INVX1 gate7288(.O (g16846), .I (g15903));
INVX1 gate7289(.O (I22820), .I (g14402));
INVX1 gate7290(.O (g16848), .I (I22820));
INVX1 gate7291(.O (I22823), .I (g13613));
INVX1 gate7292(.O (g16849), .I (I22823));
INVX1 gate7293(.O (I22828), .I (g14514));
INVX1 gate7294(.O (g16852), .I (I22828));
INVX1 gate7295(.O (I22836), .I (g13571));
INVX1 gate7296(.O (g16858), .I (I22836));
INVX1 gate7297(.O (I22842), .I (g13580));
INVX1 gate7298(.O (g16862), .I (I22842));
INVX1 gate7299(.O (I22845), .I (g13579));
INVX1 gate7300(.O (g16863), .I (I22845));
INVX1 gate7301(.O (g16867), .I (g13589));
INVX1 gate7302(.O (I22852), .I (g13600));
INVX1 gate7303(.O (g16877), .I (I22852));
INVX1 gate7304(.O (I22855), .I (g13588));
INVX1 gate7305(.O (g16878), .I (I22855));
INVX1 gate7306(.O (I22860), .I (g14885));
INVX1 gate7307(.O (g16881), .I (I22860));
INVX1 gate7308(.O (g16884), .I (g13589));
INVX1 gate7309(.O (g16895), .I (g13589));
INVX1 gate7310(.O (I22866), .I (g13612));
INVX1 gate7311(.O (g16905), .I (I22866));
INVX1 gate7312(.O (I22869), .I (g13608));
INVX1 gate7313(.O (g16906), .I (I22869));
INVX1 gate7314(.O (I22875), .I (g14966));
INVX1 gate7315(.O (g16910), .I (I22875));
INVX1 gate7316(.O (g16913), .I (g13589));
INVX1 gate7317(.O (g16924), .I (g13589));
INVX1 gate7318(.O (I22881), .I (g13622));
INVX1 gate7319(.O (g16934), .I (I22881));
INVX1 gate7320(.O (I22893), .I (g15055));
INVX1 gate7321(.O (g16940), .I (I22893));
INVX1 gate7322(.O (g16943), .I (g13589));
INVX1 gate7323(.O (g16954), .I (g13589));
INVX1 gate7324(.O (I22912), .I (g15151));
INVX1 gate7325(.O (g16971), .I (I22912));
INVX1 gate7326(.O (g16974), .I (g13589));
INVX1 gate7327(.O (g17029), .I (g14685));
INVX1 gate7328(.O (g17057), .I (g13519));
INVX1 gate7329(.O (g17063), .I (g14719));
INVX1 gate7330(.O (g17092), .I (g13530));
INVX1 gate7331(.O (g17098), .I (g14747));
INVX1 gate7332(.O (g17130), .I (g13541));
INVX1 gate7333(.O (g17136), .I (g14768));
INVX1 gate7334(.O (g17157), .I (g13552));
INVX1 gate7335(.O (I23253), .I (g13741));
INVX1 gate7336(.O (g17189), .I (I23253));
INVX1 gate7337(.O (I23274), .I (g13741));
INVX1 gate7338(.O (g17200), .I (I23274));
INVX1 gate7339(.O (g17203), .I (g13568));
INVX1 gate7340(.O (I23287), .I (g13741));
INVX1 gate7341(.O (g17207), .I (I23287));
INVX1 gate7342(.O (g17208), .I (g13576));
INVX1 gate7343(.O (I23292), .I (g13741));
INVX1 gate7344(.O (g17212), .I (I23292));
INVX1 gate7345(.O (g17214), .I (g13585));
INVX1 gate7346(.O (g17217), .I (g13605));
INVX1 gate7347(.O (I23309), .I (g16132));
INVX1 gate7348(.O (g17227), .I (I23309));
INVX1 gate7349(.O (I23314), .I (g15720));
INVX1 gate7350(.O (g17230), .I (I23314));
INVX1 gate7351(.O (I23317), .I (g16181));
INVX1 gate7352(.O (g17233), .I (I23317));
INVX1 gate7353(.O (I23323), .I (g15664));
INVX1 gate7354(.O (g17237), .I (I23323));
INVX1 gate7355(.O (I23326), .I (g15758));
INVX1 gate7356(.O (g17240), .I (I23326));
INVX1 gate7357(.O (I23329), .I (g15760));
INVX1 gate7358(.O (g17243), .I (I23329));
INVX1 gate7359(.O (I23335), .I (g16412));
INVX1 gate7360(.O (g17249), .I (I23335));
INVX1 gate7361(.O (I23338), .I (g15721));
INVX1 gate7362(.O (g17252), .I (I23338));
INVX1 gate7363(.O (I23341), .I (g15784));
INVX1 gate7364(.O (g17255), .I (I23341));
INVX1 gate7365(.O (g17258), .I (g16053));
INVX1 gate7366(.O (I23345), .I (g15723));
INVX1 gate7367(.O (g17259), .I (I23345));
INVX1 gate7368(.O (I23348), .I (g15786));
INVX1 gate7369(.O (g17262), .I (I23348));
INVX1 gate7370(.O (I23351), .I (g15788));
INVX1 gate7371(.O (g17265), .I (I23351));
INVX1 gate7372(.O (I23358), .I (g16442));
INVX1 gate7373(.O (g17272), .I (I23358));
INVX1 gate7374(.O (I23361), .I (g15759));
INVX1 gate7375(.O (g17275), .I (I23361));
INVX1 gate7376(.O (I23364), .I (g15805));
INVX1 gate7377(.O (g17278), .I (I23364));
INVX1 gate7378(.O (g17281), .I (g16081));
INVX1 gate7379(.O (I23368), .I (g16446));
INVX1 gate7380(.O (g17282), .I (I23368));
INVX1 gate7381(.O (I23371), .I (g15761));
INVX1 gate7382(.O (g17285), .I (I23371));
INVX1 gate7383(.O (I23374), .I (g15807));
INVX1 gate7384(.O (g17288), .I (I23374));
INVX1 gate7385(.O (I23377), .I (g15763));
INVX1 gate7386(.O (g17291), .I (I23377));
INVX1 gate7387(.O (I23380), .I (g15809));
INVX1 gate7388(.O (g17294), .I (I23380));
INVX1 gate7389(.O (I23383), .I (g15811));
INVX1 gate7390(.O (g17297), .I (I23383));
INVX1 gate7391(.O (I23386), .I (g13469));
INVX1 gate7392(.O (g17300), .I (I23386));
INVX1 gate7393(.O (I23392), .I (g13476));
INVX1 gate7394(.O (g17304), .I (I23392));
INVX1 gate7395(.O (I23395), .I (g15785));
INVX1 gate7396(.O (g17307), .I (I23395));
INVX1 gate7397(.O (I23398), .I (g15820));
INVX1 gate7398(.O (g17310), .I (I23398));
INVX1 gate7399(.O (g17313), .I (g16109));
INVX1 gate7400(.O (g17314), .I (g16110));
INVX1 gate7401(.O (I23403), .I (g13478));
INVX1 gate7402(.O (g17315), .I (I23403));
INVX1 gate7403(.O (I23406), .I (g15787));
INVX1 gate7404(.O (g17318), .I (I23406));
INVX1 gate7405(.O (I23409), .I (g15822));
INVX1 gate7406(.O (g17321), .I (I23409));
INVX1 gate7407(.O (I23412), .I (g13482));
INVX1 gate7408(.O (g17324), .I (I23412));
INVX1 gate7409(.O (I23415), .I (g15789));
INVX1 gate7410(.O (g17327), .I (I23415));
INVX1 gate7411(.O (I23418), .I (g15824));
INVX1 gate7412(.O (g17330), .I (I23418));
INVX1 gate7413(.O (I23421), .I (g15791));
INVX1 gate7414(.O (g17333), .I (I23421));
INVX1 gate7415(.O (I23424), .I (g15826));
INVX1 gate7416(.O (g17336), .I (I23424));
INVX1 gate7417(.O (I23430), .I (g13494));
INVX1 gate7418(.O (g17342), .I (I23430));
INVX1 gate7419(.O (I23433), .I (g15806));
INVX1 gate7420(.O (g17345), .I (I23433));
INVX1 gate7421(.O (I23436), .I (g15832));
INVX1 gate7422(.O (g17348), .I (I23436));
INVX1 gate7423(.O (g17351), .I (g16152));
INVX1 gate7424(.O (I23442), .I (g13495));
INVX1 gate7425(.O (g17354), .I (I23442));
INVX1 gate7426(.O (I23445), .I (g15808));
INVX1 gate7427(.O (g17357), .I (I23445));
INVX1 gate7428(.O (I23448), .I (g15834));
INVX1 gate7429(.O (g17360), .I (I23448));
INVX1 gate7430(.O (I23451), .I (g13497));
INVX1 gate7431(.O (g17363), .I (I23451));
INVX1 gate7432(.O (I23454), .I (g15810));
INVX1 gate7433(.O (g17366), .I (I23454));
INVX1 gate7434(.O (I23457), .I (g15836));
INVX1 gate7435(.O (g17369), .I (I23457));
INVX1 gate7436(.O (I23460), .I (g13501));
INVX1 gate7437(.O (g17372), .I (I23460));
INVX1 gate7438(.O (I23463), .I (g15812));
INVX1 gate7439(.O (g17375), .I (I23463));
INVX1 gate7440(.O (I23466), .I (g15838));
INVX1 gate7441(.O (g17378), .I (I23466));
INVX1 gate7442(.O (I23472), .I (g13510));
INVX1 gate7443(.O (g17384), .I (I23472));
INVX1 gate7444(.O (I23475), .I (g15821));
INVX1 gate7445(.O (g17387), .I (I23475));
INVX1 gate7446(.O (I23478), .I (g15844));
INVX1 gate7447(.O (g17390), .I (I23478));
INVX1 gate7448(.O (g17394), .I (g16197));
INVX1 gate7449(.O (I23487), .I (g13511));
INVX1 gate7450(.O (g17399), .I (I23487));
INVX1 gate7451(.O (I23490), .I (g15823));
INVX1 gate7452(.O (g17402), .I (I23490));
INVX1 gate7453(.O (I23493), .I (g15846));
INVX1 gate7454(.O (g17405), .I (I23493));
INVX1 gate7455(.O (I23498), .I (g13512));
INVX1 gate7456(.O (g17410), .I (I23498));
INVX1 gate7457(.O (I23501), .I (g15825));
INVX1 gate7458(.O (g17413), .I (I23501));
INVX1 gate7459(.O (I23504), .I (g15848));
INVX1 gate7460(.O (g17416), .I (I23504));
INVX1 gate7461(.O (I23507), .I (g13514));
INVX1 gate7462(.O (g17419), .I (I23507));
INVX1 gate7463(.O (I23510), .I (g15827));
INVX1 gate7464(.O (g17422), .I (I23510));
INVX1 gate7465(.O (I23513), .I (g15850));
INVX1 gate7466(.O (g17425), .I (I23513));
INVX1 gate7467(.O (I23518), .I (g15856));
INVX1 gate7468(.O (g17430), .I (I23518));
INVX1 gate7469(.O (I23521), .I (g13518));
INVX1 gate7470(.O (g17433), .I (I23521));
INVX1 gate7471(.O (I23524), .I (g15833));
INVX1 gate7472(.O (g17436), .I (I23524));
INVX1 gate7473(.O (I23527), .I (g15858));
INVX1 gate7474(.O (g17439), .I (I23527));
INVX1 gate7475(.O (I23530), .I (g14885));
INVX1 gate7476(.O (g17442), .I (I23530));
INVX1 gate7477(.O (g17445), .I (g16250));
INVX1 gate7478(.O (I23539), .I (g13524));
INVX1 gate7479(.O (g17451), .I (I23539));
INVX1 gate7480(.O (I23542), .I (g15835));
INVX1 gate7481(.O (g17454), .I (I23542));
INVX1 gate7482(.O (I23545), .I (g15867));
INVX1 gate7483(.O (g17457), .I (I23545));
INVX1 gate7484(.O (I23553), .I (g13525));
INVX1 gate7485(.O (g17465), .I (I23553));
INVX1 gate7486(.O (I23556), .I (g15837));
INVX1 gate7487(.O (g17468), .I (I23556));
INVX1 gate7488(.O (I23559), .I (g15869));
INVX1 gate7489(.O (g17471), .I (I23559));
INVX1 gate7490(.O (I23564), .I (g13526));
INVX1 gate7491(.O (g17476), .I (I23564));
INVX1 gate7492(.O (I23567), .I (g15839));
INVX1 gate7493(.O (g17479), .I (I23567));
INVX1 gate7494(.O (I23570), .I (g15871));
INVX1 gate7495(.O (g17482), .I (I23570));
INVX1 gate7496(.O (I23575), .I (g15843));
INVX1 gate7497(.O (g17487), .I (I23575));
INVX1 gate7498(.O (I23578), .I (g15879));
INVX1 gate7499(.O (g17490), .I (I23578));
INVX1 gate7500(.O (I23581), .I (g13528));
INVX1 gate7501(.O (g17493), .I (I23581));
INVX1 gate7502(.O (I23584), .I (g15845));
INVX1 gate7503(.O (g17496), .I (I23584));
INVX1 gate7504(.O (g17499), .I (g16292));
INVX1 gate7505(.O (I23588), .I (g14885));
INVX1 gate7506(.O (g17500), .I (I23588));
INVX1 gate7507(.O (I23591), .I (g14885));
INVX1 gate7508(.O (g17503), .I (I23591));
INVX1 gate7509(.O (I23599), .I (g15887));
INVX1 gate7510(.O (g17511), .I (I23599));
INVX1 gate7511(.O (I23602), .I (g13529));
INVX1 gate7512(.O (g17514), .I (I23602));
INVX1 gate7513(.O (I23605), .I (g15847));
INVX1 gate7514(.O (g17517), .I (I23605));
INVX1 gate7515(.O (I23608), .I (g15889));
INVX1 gate7516(.O (g17520), .I (I23608));
INVX1 gate7517(.O (I23611), .I (g14966));
INVX1 gate7518(.O (g17523), .I (I23611));
INVX1 gate7519(.O (I23619), .I (g13535));
INVX1 gate7520(.O (g17531), .I (I23619));
INVX1 gate7521(.O (I23622), .I (g15849));
INVX1 gate7522(.O (g17534), .I (I23622));
INVX1 gate7523(.O (I23625), .I (g15898));
INVX1 gate7524(.O (g17537), .I (I23625));
INVX1 gate7525(.O (I23633), .I (g13536));
INVX1 gate7526(.O (g17545), .I (I23633));
INVX1 gate7527(.O (I23636), .I (g15851));
INVX1 gate7528(.O (g17548), .I (I23636));
INVX1 gate7529(.O (I23639), .I (g15900));
INVX1 gate7530(.O (g17551), .I (I23639));
INVX1 gate7531(.O (I23645), .I (g13537));
INVX1 gate7532(.O (g17557), .I (I23645));
INVX1 gate7533(.O (I23648), .I (g15857));
INVX1 gate7534(.O (g17560), .I (I23648));
INVX1 gate7535(.O (I23651), .I (g13538));
INVX1 gate7536(.O (g17563), .I (I23651));
INVX1 gate7537(.O (g17566), .I (g16346));
INVX1 gate7538(.O (I23655), .I (g14831));
INVX1 gate7539(.O (g17567), .I (I23655));
INVX1 gate7540(.O (I23658), .I (g14885));
INVX1 gate7541(.O (g17570), .I (I23658));
INVX1 gate7542(.O (I23661), .I (g16085));
INVX1 gate7543(.O (g17573), .I (I23661));
INVX1 gate7544(.O (I23667), .I (g15866));
INVX1 gate7545(.O (g17579), .I (I23667));
INVX1 gate7546(.O (I23670), .I (g15912));
INVX1 gate7547(.O (g17582), .I (I23670));
INVX1 gate7548(.O (I23673), .I (g13539));
INVX1 gate7549(.O (g17585), .I (I23673));
INVX1 gate7550(.O (I23676), .I (g15868));
INVX1 gate7551(.O (g17588), .I (I23676));
INVX1 gate7552(.O (I23679), .I (g14966));
INVX1 gate7553(.O (g17591), .I (I23679));
INVX1 gate7554(.O (I23682), .I (g14966));
INVX1 gate7555(.O (g17594), .I (I23682));
INVX1 gate7556(.O (I23689), .I (g15920));
INVX1 gate7557(.O (g17601), .I (I23689));
INVX1 gate7558(.O (I23692), .I (g13540));
INVX1 gate7559(.O (g17604), .I (I23692));
INVX1 gate7560(.O (I23695), .I (g15870));
INVX1 gate7561(.O (g17607), .I (I23695));
INVX1 gate7562(.O (I23698), .I (g15922));
INVX1 gate7563(.O (g17610), .I (I23698));
INVX1 gate7564(.O (I23701), .I (g15055));
INVX1 gate7565(.O (g17613), .I (I23701));
INVX1 gate7566(.O (I23709), .I (g13546));
INVX1 gate7567(.O (g17621), .I (I23709));
INVX1 gate7568(.O (I23712), .I (g15872));
INVX1 gate7569(.O (g17624), .I (I23712));
INVX1 gate7570(.O (I23715), .I (g15931));
INVX1 gate7571(.O (g17627), .I (I23715));
INVX1 gate7572(.O (I23725), .I (g13547));
INVX1 gate7573(.O (g17637), .I (I23725));
INVX1 gate7574(.O (g17640), .I (g13873));
INVX1 gate7575(.O (I23729), .I (g14337));
INVX1 gate7576(.O (g17645), .I (I23729));
INVX1 gate7577(.O (g17648), .I (g16384));
INVX1 gate7578(.O (I23733), .I (g14831));
INVX1 gate7579(.O (g17649), .I (I23733));
INVX1 gate7580(.O (I23739), .I (g13548));
INVX1 gate7581(.O (g17655), .I (I23739));
INVX1 gate7582(.O (I23742), .I (g15888));
INVX1 gate7583(.O (g17658), .I (I23742));
INVX1 gate7584(.O (I23745), .I (g13549));
INVX1 gate7585(.O (g17661), .I (I23745));
INVX1 gate7586(.O (I23748), .I (g14904));
INVX1 gate7587(.O (g17664), .I (I23748));
INVX1 gate7588(.O (I23751), .I (g14966));
INVX1 gate7589(.O (g17667), .I (I23751));
INVX1 gate7590(.O (I23754), .I (g16123));
INVX1 gate7591(.O (g17670), .I (I23754));
INVX1 gate7592(.O (I23760), .I (g15897));
INVX1 gate7593(.O (g17676), .I (I23760));
INVX1 gate7594(.O (I23763), .I (g15941));
INVX1 gate7595(.O (g17679), .I (I23763));
INVX1 gate7596(.O (I23766), .I (g13550));
INVX1 gate7597(.O (g17682), .I (I23766));
INVX1 gate7598(.O (I23769), .I (g15899));
INVX1 gate7599(.O (g17685), .I (I23769));
INVX1 gate7600(.O (I23772), .I (g15055));
INVX1 gate7601(.O (g17688), .I (I23772));
INVX1 gate7602(.O (I23775), .I (g15055));
INVX1 gate7603(.O (g17691), .I (I23775));
INVX1 gate7604(.O (I23782), .I (g15949));
INVX1 gate7605(.O (g17698), .I (I23782));
INVX1 gate7606(.O (I23785), .I (g13551));
INVX1 gate7607(.O (g17701), .I (I23785));
INVX1 gate7608(.O (I23788), .I (g15901));
INVX1 gate7609(.O (g17704), .I (I23788));
INVX1 gate7610(.O (I23791), .I (g15951));
INVX1 gate7611(.O (g17707), .I (I23791));
INVX1 gate7612(.O (I23794), .I (g15151));
INVX1 gate7613(.O (g17710), .I (I23794));
INVX1 gate7614(.O (g17720), .I (g15853));
INVX1 gate7615(.O (g17724), .I (g13886));
INVX1 gate7616(.O (I23817), .I (g13557));
INVX1 gate7617(.O (g17738), .I (I23817));
INVX1 gate7618(.O (g17741), .I (g13895));
INVX1 gate7619(.O (I23821), .I (g14337));
INVX1 gate7620(.O (g17746), .I (I23821));
INVX1 gate7621(.O (I23824), .I (g14904));
INVX1 gate7622(.O (g17749), .I (I23824));
INVX1 gate7623(.O (I23830), .I (g13558));
INVX1 gate7624(.O (g17755), .I (I23830));
INVX1 gate7625(.O (I23833), .I (g15921));
INVX1 gate7626(.O (g17758), .I (I23833));
INVX1 gate7627(.O (I23836), .I (g13559));
INVX1 gate7628(.O (g17761), .I (I23836));
INVX1 gate7629(.O (I23839), .I (g14985));
INVX1 gate7630(.O (g17764), .I (I23839));
INVX1 gate7631(.O (I23842), .I (g15055));
INVX1 gate7632(.O (g17767), .I (I23842));
INVX1 gate7633(.O (I23845), .I (g16174));
INVX1 gate7634(.O (g17770), .I (I23845));
INVX1 gate7635(.O (I23851), .I (g15930));
INVX1 gate7636(.O (g17776), .I (I23851));
INVX1 gate7637(.O (I23854), .I (g15970));
INVX1 gate7638(.O (g17779), .I (I23854));
INVX1 gate7639(.O (I23857), .I (g13560));
INVX1 gate7640(.O (g17782), .I (I23857));
INVX1 gate7641(.O (I23860), .I (g15932));
INVX1 gate7642(.O (g17785), .I (I23860));
INVX1 gate7643(.O (I23863), .I (g15151));
INVX1 gate7644(.O (g17788), .I (I23863));
INVX1 gate7645(.O (I23866), .I (g15151));
INVX1 gate7646(.O (g17791), .I (I23866));
INVX1 gate7647(.O (I23874), .I (g15797));
INVX1 gate7648(.O (g17799), .I (I23874));
INVX1 gate7649(.O (g17802), .I (g13907));
INVX1 gate7650(.O (I23888), .I (g14685));
INVX1 gate7651(.O (g17815), .I (I23888));
INVX1 gate7652(.O (g17825), .I (g13927));
INVX1 gate7653(.O (I23904), .I (g13561));
INVX1 gate7654(.O (g17839), .I (I23904));
INVX1 gate7655(.O (g17842), .I (g13936));
INVX1 gate7656(.O (I23908), .I (g14337));
INVX1 gate7657(.O (g17847), .I (I23908));
INVX1 gate7658(.O (I23911), .I (g14985));
INVX1 gate7659(.O (g17850), .I (I23911));
INVX1 gate7660(.O (I23917), .I (g13562));
INVX1 gate7661(.O (g17856), .I (I23917));
INVX1 gate7662(.O (I23920), .I (g15950));
INVX1 gate7663(.O (g17859), .I (I23920));
INVX1 gate7664(.O (I23923), .I (g13563));
INVX1 gate7665(.O (g17862), .I (I23923));
INVX1 gate7666(.O (I23926), .I (g15074));
INVX1 gate7667(.O (g17865), .I (I23926));
INVX1 gate7668(.O (I23929), .I (g15151));
INVX1 gate7669(.O (g17868), .I (I23929));
INVX1 gate7670(.O (I23932), .I (g16233));
INVX1 gate7671(.O (g17871), .I (I23932));
INVX1 gate7672(.O (g17878), .I (g15830));
INVX1 gate7673(.O (g17882), .I (g13946));
INVX1 gate7674(.O (g17892), .I (g13954));
INVX1 gate7675(.O (g17893), .I (g14165));
INVX1 gate7676(.O (I23954), .I (g16154));
INVX1 gate7677(.O (g17903), .I (I23954));
INVX1 gate7678(.O (g17914), .I (g13963));
INVX1 gate7679(.O (I23976), .I (g14719));
INVX1 gate7680(.O (g17927), .I (I23976));
INVX1 gate7681(.O (g17937), .I (g13983));
INVX1 gate7682(.O (I23992), .I (g13564));
INVX1 gate7683(.O (g17951), .I (I23992));
INVX1 gate7684(.O (g17954), .I (g13992));
INVX1 gate7685(.O (I23996), .I (g14337));
INVX1 gate7686(.O (g17959), .I (I23996));
INVX1 gate7687(.O (I23999), .I (g15074));
INVX1 gate7688(.O (g17962), .I (I23999));
INVX1 gate7689(.O (g17969), .I (g15841));
INVX1 gate7690(.O (g17974), .I (g14001));
INVX1 gate7691(.O (g17984), .I (g14008));
INVX1 gate7692(.O (g17988), .I (g14685));
INVX1 gate7693(.O (g17991), .I (g14450));
INVX1 gate7694(.O (g17993), .I (g14016));
INVX1 gate7695(.O (g18003), .I (g14024));
INVX1 gate7696(.O (g18004), .I (g14280));
INVX1 gate7697(.O (I24049), .I (g16213));
INVX1 gate7698(.O (g18014), .I (I24049));
INVX1 gate7699(.O (g18025), .I (g14033));
INVX1 gate7700(.O (I24071), .I (g14747));
INVX1 gate7701(.O (g18038), .I (I24071));
INVX1 gate7702(.O (g18048), .I (g14053));
INVX1 gate7703(.O (g18063), .I (g15660));
INVX1 gate7704(.O (g18070), .I (g15854));
INVX1 gate7705(.O (g18074), .I (g14062));
INVX1 gate7706(.O (g18084), .I (g14068));
INVX1 gate7707(.O (g18089), .I (g14355));
INVX1 gate7708(.O (g18091), .I (g14092));
INVX1 gate7709(.O (g18101), .I (g14099));
INVX1 gate7710(.O (g18105), .I (g14719));
INVX1 gate7711(.O (g18108), .I (g14537));
INVX1 gate7712(.O (g18110), .I (g14107));
INVX1 gate7713(.O (g18120), .I (g14115));
INVX1 gate7714(.O (g18121), .I (g14402));
INVX1 gate7715(.O (I24144), .I (g16278));
INVX1 gate7716(.O (g18131), .I (I24144));
INVX1 gate7717(.O (g18142), .I (g14124));
INVX1 gate7718(.O (I24166), .I (g14768));
INVX1 gate7719(.O (g18155), .I (I24166));
INVX1 gate7720(.O (I24171), .I (g16439));
INVX1 gate7721(.O (g18166), .I (I24171));
INVX1 gate7722(.O (g18170), .I (g15877));
INVX1 gate7723(.O (g18174), .I (g14148));
INVX1 gate7724(.O (g18179), .I (g14153));
INVX1 gate7725(.O (g18188), .I (g14252));
INVX1 gate7726(.O (g18190), .I (g14177));
INVX1 gate7727(.O (g18200), .I (g14183));
INVX1 gate7728(.O (g18205), .I (g14467));
INVX1 gate7729(.O (g18207), .I (g14207));
INVX1 gate7730(.O (g18217), .I (g14214));
INVX1 gate7731(.O (g18221), .I (g14747));
INVX1 gate7732(.O (g18224), .I (g14592));
INVX1 gate7733(.O (g18226), .I (g14222));
INVX1 gate7734(.O (g18236), .I (g14230));
INVX1 gate7735(.O (g18237), .I (g14514));
INVX1 gate7736(.O (I24247), .I (g16337));
INVX1 gate7737(.O (g18247), .I (I24247));
INVX1 gate7738(.O (I24258), .I (g16463));
INVX1 gate7739(.O (g18258), .I (I24258));
INVX1 gate7740(.O (g18261), .I (g15719));
INVX1 gate7741(.O (g18265), .I (g14238));
INVX1 gate7742(.O (g18275), .I (g14171));
INVX1 gate7743(.O (I24285), .I (g15992));
INVX1 gate7744(.O (g18278), .I (I24285));
INVX1 gate7745(.O (g18281), .I (g14263));
INVX1 gate7746(.O (g18286), .I (g14268));
INVX1 gate7747(.O (g18295), .I (g14374));
INVX1 gate7748(.O (g18297), .I (g14292));
INVX1 gate7749(.O (g18307), .I (g14298));
INVX1 gate7750(.O (g18312), .I (g14554));
INVX1 gate7751(.O (g18314), .I (g14322));
INVX1 gate7752(.O (g18324), .I (g14329));
INVX1 gate7753(.O (g18328), .I (g14768));
INVX1 gate7754(.O (g18331), .I (g14626));
INVX1 gate7755(.O (I24346), .I (g15873));
INVX1 gate7756(.O (g18334), .I (I24346));
INVX1 gate7757(.O (g18337), .I (g15757));
INVX1 gate7758(.O (g18341), .I (g14342));
INVX1 gate7759(.O (g18351), .I (g13741));
INVX1 gate7760(.O (g18353), .I (g13918));
INVX1 gate7761(.O (I24368), .I (g15990));
INVX1 gate7762(.O (g18355), .I (I24368));
INVX1 gate7763(.O (g18358), .I (g14360));
INVX1 gate7764(.O (g18368), .I (g14286));
INVX1 gate7765(.O (I24394), .I (g15995));
INVX1 gate7766(.O (g18371), .I (I24394));
INVX1 gate7767(.O (g18374), .I (g14385));
INVX1 gate7768(.O (g18379), .I (g14390));
INVX1 gate7769(.O (g18388), .I (g14486));
INVX1 gate7770(.O (g18390), .I (g14414));
INVX1 gate7771(.O (g18400), .I (g14420));
INVX1 gate7772(.O (g18405), .I (g14609));
INVX1 gate7773(.O (g18407), .I (g15959));
INVX1 gate7774(.O (g18414), .I (g15718));
INVX1 gate7775(.O (g18415), .I (g15783));
INVX1 gate7776(.O (g18429), .I (g14831));
INVX1 gate7777(.O (I24459), .I (g13599));
INVX1 gate7778(.O (g18432), .I (I24459));
INVX1 gate7779(.O (g18435), .I (g14359));
INVX1 gate7780(.O (g18436), .I (g14454));
INVX1 gate7781(.O (g18446), .I (g13741));
INVX1 gate7782(.O (g18448), .I (g13974));
INVX1 gate7783(.O (I24481), .I (g15993));
INVX1 gate7784(.O (g18450), .I (I24481));
INVX1 gate7785(.O (g18453), .I (g14472));
INVX1 gate7786(.O (g18463), .I (g14408));
INVX1 gate7787(.O (I24507), .I (g15999));
INVX1 gate7788(.O (g18466), .I (I24507));
INVX1 gate7789(.O (g18469), .I (g14497));
INVX1 gate7790(.O (g18474), .I (g14502));
INVX1 gate7791(.O (g18483), .I (g14573));
INVX1 gate7792(.O (g18485), .I (g15756));
INVX1 gate7793(.O (g18486), .I (g15804));
INVX1 gate7794(.O (g18490), .I (g13565));
INVX1 gate7795(.O (g18502), .I (g14904));
INVX1 gate7796(.O (I24560), .I (g13611));
INVX1 gate7797(.O (g18505), .I (I24560));
INVX1 gate7798(.O (g18508), .I (g14471));
INVX1 gate7799(.O (g18509), .I (g14541));
INVX1 gate7800(.O (g18519), .I (g13741));
INVX1 gate7801(.O (g18521), .I (g14044));
INVX1 gate7802(.O (I24582), .I (g15996));
INVX1 gate7803(.O (g18523), .I (I24582));
INVX1 gate7804(.O (g18526), .I (g14559));
INVX1 gate7805(.O (g18536), .I (g14520));
INVX1 gate7806(.O (I24608), .I (g16006));
INVX1 gate7807(.O (g18539), .I (I24608));
INVX1 gate7808(.O (g18543), .I (g15819));
INVX1 gate7809(.O (g18552), .I (g16154));
INVX1 gate7810(.O (g18554), .I (g13573));
INVX1 gate7811(.O (g18566), .I (g14985));
INVX1 gate7812(.O (I24662), .I (g13621));
INVX1 gate7813(.O (g18569), .I (I24662));
INVX1 gate7814(.O (g18572), .I (g14558));
INVX1 gate7815(.O (g18573), .I (g14596));
INVX1 gate7816(.O (g18583), .I (g13741));
INVX1 gate7817(.O (g18585), .I (g14135));
INVX1 gate7818(.O (I24684), .I (g16000));
INVX1 gate7819(.O (g18587), .I (I24684));
INVX1 gate7820(.O (g18593), .I (g15831));
INVX1 gate7821(.O (g18602), .I (g16213));
INVX1 gate7822(.O (g18604), .I (g13582));
INVX1 gate7823(.O (g18616), .I (g15074));
INVX1 gate7824(.O (I24732), .I (g13633));
INVX1 gate7825(.O (g18619), .I (I24732));
INVX1 gate7826(.O (g18622), .I (g14613));
INVX1 gate7827(.O (g18634), .I (g16278));
INVX1 gate7828(.O (g18636), .I (g13602));
INVX1 gate7829(.O (g18643), .I (g16337));
INVX1 gate7830(.O (g18646), .I (g16341));
INVX1 gate7831(.O (g18656), .I (g14776));
INVX1 gate7832(.O (g18670), .I (g14797));
INVX1 gate7833(.O (g18679), .I (g14811));
INVX1 gate7834(.O (g18691), .I (g14885));
INVX1 gate7835(.O (g18692), .I (g14837));
INVX1 gate7836(.O (g18699), .I (g14849));
INVX1 gate7837(.O (g18708), .I (g14863));
INVX1 gate7838(.O (g18720), .I (g14895));
INVX1 gate7839(.O (g18725), .I (g13865));
INVX1 gate7840(.O (g18727), .I (g14966));
INVX1 gate7841(.O (g18728), .I (g14910));
INVX1 gate7842(.O (g18735), .I (g14922));
INVX1 gate7843(.O (g18744), .I (g14936));
INVX1 gate7844(.O (g18756), .I (g14960));
INVX1 gate7845(.O (g18757), .I (g14963));
INVX1 gate7846(.O (g18758), .I (g14976));
INVX1 gate7847(.O (g18764), .I (g15055));
INVX1 gate7848(.O (g18765), .I (g14991));
INVX1 gate7849(.O (g18772), .I (g15003));
INVX1 gate7850(.O (g18783), .I (g15034));
INVX1 gate7851(.O (g18784), .I (g15037));
INVX1 gate7852(.O (g18785), .I (g15040));
INVX1 gate7853(.O (g18786), .I (g15043));
INVX1 gate7854(.O (g18787), .I (g15049));
INVX1 gate7855(.O (g18788), .I (g15052));
INVX1 gate7856(.O (g18789), .I (g15065));
INVX1 gate7857(.O (g18795), .I (g15151));
INVX1 gate7858(.O (g18796), .I (g15080));
INVX1 gate7859(.O (g18805), .I (g15106));
INVX1 gate7860(.O (g18806), .I (g15109));
INVX1 gate7861(.O (g18807), .I (g15112));
INVX1 gate7862(.O (g18808), .I (g15115));
INVX1 gate7863(.O (g18809), .I (g15130));
INVX1 gate7864(.O (g18810), .I (g15133));
INVX1 gate7865(.O (g18811), .I (g15136));
INVX1 gate7866(.O (g18812), .I (g15139));
INVX1 gate7867(.O (g18813), .I (g15145));
INVX1 gate7868(.O (g18814), .I (g15148));
INVX1 gate7869(.O (g18815), .I (g15161));
INVX1 gate7870(.O (g18822), .I (g15179));
INVX1 gate7871(.O (g18823), .I (g15182));
INVX1 gate7872(.O (g18824), .I (g15185));
INVX1 gate7873(.O (g18825), .I (g15198));
INVX1 gate7874(.O (g18826), .I (g15201));
INVX1 gate7875(.O (g18827), .I (g15204));
INVX1 gate7876(.O (g18828), .I (g15207));
INVX1 gate7877(.O (g18829), .I (g15222));
INVX1 gate7878(.O (g18830), .I (g15225));
INVX1 gate7879(.O (g18831), .I (g15228));
INVX1 gate7880(.O (g18832), .I (g15231));
INVX1 gate7881(.O (g18833), .I (g15237));
INVX1 gate7882(.O (g18834), .I (g15240));
INVX1 gate7883(.O (g18838), .I (g15248));
INVX1 gate7884(.O (g18839), .I (g15251));
INVX1 gate7885(.O (g18840), .I (g15254));
INVX1 gate7886(.O (g18841), .I (g15265));
INVX1 gate7887(.O (g18842), .I (g15268));
INVX1 gate7888(.O (g18843), .I (g15271));
INVX1 gate7889(.O (g18844), .I (g15284));
INVX1 gate7890(.O (g18845), .I (g15287));
INVX1 gate7891(.O (g18846), .I (g15290));
INVX1 gate7892(.O (g18847), .I (g15293));
INVX1 gate7893(.O (g18848), .I (g15308));
INVX1 gate7894(.O (g18849), .I (g15311));
INVX1 gate7895(.O (g18850), .I (g15314));
INVX1 gate7896(.O (g18851), .I (g15317));
INVX1 gate7897(.O (g18853), .I (g15326));
INVX1 gate7898(.O (g18854), .I (g15329));
INVX1 gate7899(.O (g18855), .I (g15332));
INVX1 gate7900(.O (g18856), .I (g15340));
INVX1 gate7901(.O (g18857), .I (g15343));
INVX1 gate7902(.O (g18858), .I (g15346));
INVX1 gate7903(.O (g18859), .I (g15357));
INVX1 gate7904(.O (g18860), .I (g15360));
INVX1 gate7905(.O (g18861), .I (g15363));
INVX1 gate7906(.O (g18862), .I (g15376));
INVX1 gate7907(.O (g18863), .I (g15379));
INVX1 gate7908(.O (g18864), .I (g15382));
INVX1 gate7909(.O (g18865), .I (g15385));
INVX1 gate7910(.O (I24894), .I (g14797));
INVX1 gate7911(.O (g18869), .I (I24894));
INVX1 gate7912(.O (g18870), .I (g15393));
INVX1 gate7913(.O (g18871), .I (g15396));
INVX1 gate7914(.O (g18872), .I (g15399));
INVX1 gate7915(.O (g18873), .I (g15404));
INVX1 gate7916(.O (g18874), .I (g15412));
INVX1 gate7917(.O (g18875), .I (g15415));
INVX1 gate7918(.O (g18876), .I (g15418));
INVX1 gate7919(.O (g18877), .I (g15426));
INVX1 gate7920(.O (g18878), .I (g15429));
INVX1 gate7921(.O (g18879), .I (g15432));
INVX1 gate7922(.O (g18880), .I (g15443));
INVX1 gate7923(.O (g18881), .I (g15446));
INVX1 gate7924(.O (g18882), .I (g15449));
INVX1 gate7925(.O (g18884), .I (g13469));
INVX1 gate7926(.O (I24913), .I (g15800));
INVX1 gate7927(.O (g18886), .I (I24913));
INVX1 gate7928(.O (I24916), .I (g14776));
INVX1 gate7929(.O (g18890), .I (I24916));
INVX1 gate7930(.O (g18891), .I (g15461));
INVX1 gate7931(.O (g18892), .I (g15464));
INVX1 gate7932(.O (g18893), .I (g15467));
INVX1 gate7933(.O (g18894), .I (g15471));
INVX1 gate7934(.O (I24923), .I (g14849));
INVX1 gate7935(.O (g18895), .I (I24923));
INVX1 gate7936(.O (g18896), .I (g15477));
INVX1 gate7937(.O (g18897), .I (g15480));
INVX1 gate7938(.O (g18898), .I (g15483));
INVX1 gate7939(.O (g18899), .I (g15488));
INVX1 gate7940(.O (g18900), .I (g15496));
INVX1 gate7941(.O (g18901), .I (g15499));
INVX1 gate7942(.O (g18902), .I (g15502));
INVX1 gate7943(.O (g18903), .I (g15510));
INVX1 gate7944(.O (g18904), .I (g15513));
INVX1 gate7945(.O (g18905), .I (g15516));
INVX1 gate7946(.O (g18908), .I (g15521));
INVX1 gate7947(.O (g18909), .I (g15528));
INVX1 gate7948(.O (g18910), .I (g15531));
INVX1 gate7949(.O (g18911), .I (g15534));
INVX1 gate7950(.O (g18912), .I (g15537));
INVX1 gate7951(.O (I24943), .I (g14811));
INVX1 gate7952(.O (g18913), .I (I24943));
INVX1 gate7953(.O (g18914), .I (g15547));
INVX1 gate7954(.O (g18915), .I (g15550));
INVX1 gate7955(.O (g18916), .I (g15553));
INVX1 gate7956(.O (g18917), .I (g15557));
INVX1 gate7957(.O (I24950), .I (g14922));
INVX1 gate7958(.O (g18918), .I (I24950));
INVX1 gate7959(.O (g18919), .I (g15563));
INVX1 gate7960(.O (g18920), .I (g15566));
INVX1 gate7961(.O (g18921), .I (g15569));
INVX1 gate7962(.O (g18922), .I (g15574));
INVX1 gate7963(.O (g18923), .I (g15582));
INVX1 gate7964(.O (g18924), .I (g15585));
INVX1 gate7965(.O (g18925), .I (g15588));
INVX1 gate7966(.O (g18926), .I (g15596));
INVX1 gate7967(.O (g18927), .I (g15599));
INVX1 gate7968(.O (g18928), .I (g15606));
INVX1 gate7969(.O (g18929), .I (g15609));
INVX1 gate7970(.O (g18930), .I (g15612));
INVX1 gate7971(.O (g18931), .I (g15615));
INVX1 gate7972(.O (I24966), .I (g14863));
INVX1 gate7973(.O (g18932), .I (I24966));
INVX1 gate7974(.O (g18933), .I (g15625));
INVX1 gate7975(.O (g18934), .I (g15628));
INVX1 gate7976(.O (g18935), .I (g15631));
INVX1 gate7977(.O (g18936), .I (g15635));
INVX1 gate7978(.O (I24973), .I (g15003));
INVX1 gate7979(.O (g18937), .I (I24973));
INVX1 gate7980(.O (g18938), .I (g15641));
INVX1 gate7981(.O (g18939), .I (g15644));
INVX1 gate7982(.O (g18940), .I (g15647));
INVX1 gate7983(.O (g18941), .I (g15652));
INVX1 gate7984(.O (g18943), .I (g15655));
INVX1 gate7985(.O (I24982), .I (g14347));
INVX1 gate7986(.O (g18944), .I (I24982));
INVX1 gate7987(.O (g18945), .I (g15667));
INVX1 gate7988(.O (g18946), .I (g15672));
INVX1 gate7989(.O (g18947), .I (g15675));
INVX1 gate7990(.O (g18948), .I (g15682));
INVX1 gate7991(.O (g18949), .I (g15685));
INVX1 gate7992(.O (g18950), .I (g15688));
INVX1 gate7993(.O (g18951), .I (g15691));
INVX1 gate7994(.O (I24992), .I (g14936));
INVX1 gate7995(.O (g18952), .I (I24992));
INVX1 gate7996(.O (g18953), .I (g15701));
INVX1 gate7997(.O (g18954), .I (g15704));
INVX1 gate7998(.O (g18955), .I (g15707));
INVX1 gate7999(.O (g18956), .I (g15711));
INVX1 gate8000(.O (g18958), .I (g15714));
INVX1 gate8001(.O (I25001), .I (g14244));
INVX1 gate8002(.O (g18959), .I (I25001));
INVX1 gate8003(.O (I25004), .I (g14459));
INVX1 gate8004(.O (g18960), .I (I25004));
INVX1 gate8005(.O (g18961), .I (g15726));
INVX1 gate8006(.O (g18962), .I (g15731));
INVX1 gate8007(.O (g18963), .I (g15734));
INVX1 gate8008(.O (g18964), .I (g15741));
INVX1 gate8009(.O (g18965), .I (g15744));
INVX1 gate8010(.O (g18966), .I (g15747));
INVX1 gate8011(.O (g18967), .I (g15750));
INVX1 gate8012(.O (I25015), .I (g14158));
INVX1 gate8013(.O (g18969), .I (I25015));
INVX1 gate8014(.O (I25018), .I (g14366));
INVX1 gate8015(.O (g18970), .I (I25018));
INVX1 gate8016(.O (I25021), .I (g14546));
INVX1 gate8017(.O (g18971), .I (I25021));
INVX1 gate8018(.O (g18972), .I (g15766));
INVX1 gate8019(.O (g18973), .I (g15771));
INVX1 gate8020(.O (g18974), .I (g15774));
INVX1 gate8021(.O (g18976), .I (g15777));
INVX1 gate8022(.O (I25037), .I (g14071));
INVX1 gate8023(.O (g18981), .I (I25037));
INVX1 gate8024(.O (I25041), .I (g14895));
INVX1 gate8025(.O (g18983), .I (I25041));
INVX1 gate8026(.O (I25044), .I (g14273));
INVX1 gate8027(.O (g18984), .I (I25044));
INVX1 gate8028(.O (I25047), .I (g14478));
INVX1 gate8029(.O (g18985), .I (I25047));
INVX1 gate8030(.O (I25050), .I (g14601));
INVX1 gate8031(.O (g18986), .I (I25050));
INVX1 gate8032(.O (g18987), .I (g15794));
INVX1 gate8033(.O (I25054), .I (g14837));
INVX1 gate8034(.O (g18988), .I (I25054));
INVX1 gate8035(.O (I25057), .I (g14186));
INVX1 gate8036(.O (g18989), .I (I25057));
INVX1 gate8037(.O (I25061), .I (g14976));
INVX1 gate8038(.O (g18991), .I (I25061));
INVX1 gate8039(.O (I25064), .I (g14395));
INVX1 gate8040(.O (g18992), .I (I25064));
INVX1 gate8041(.O (I25067), .I (g14565));
INVX1 gate8042(.O (g18993), .I (I25067));
INVX1 gate8043(.O (I25071), .I (g14910));
INVX1 gate8044(.O (g18995), .I (I25071));
INVX1 gate8045(.O (I25074), .I (g14301));
INVX1 gate8046(.O (g18996), .I (I25074));
INVX1 gate8047(.O (I25078), .I (g15065));
INVX1 gate8048(.O (g18998), .I (I25078));
INVX1 gate8049(.O (I25081), .I (g14507));
INVX1 gate8050(.O (g18999), .I (I25081));
INVX1 gate8051(.O (I25084), .I (g14885));
INVX1 gate8052(.O (g19000), .I (I25084));
INVX1 gate8053(.O (g19001), .I (g14071));
INVX1 gate8054(.O (I25089), .I (g14991));
INVX1 gate8055(.O (g19008), .I (I25089));
INVX1 gate8056(.O (I25092), .I (g14423));
INVX1 gate8057(.O (g19009), .I (I25092));
INVX1 gate8058(.O (I25096), .I (g15161));
INVX1 gate8059(.O (g19011), .I (I25096));
INVX1 gate8060(.O (I25099), .I (g19000));
INVX1 gate8061(.O (g19012), .I (I25099));
INVX1 gate8062(.O (I25102), .I (g18944));
INVX1 gate8063(.O (g19013), .I (I25102));
INVX1 gate8064(.O (I25105), .I (g18959));
INVX1 gate8065(.O (g19014), .I (I25105));
INVX1 gate8066(.O (I25108), .I (g18969));
INVX1 gate8067(.O (g19015), .I (I25108));
INVX1 gate8068(.O (I25111), .I (g18981));
INVX1 gate8069(.O (g19016), .I (I25111));
INVX1 gate8070(.O (I25114), .I (g18983));
INVX1 gate8071(.O (g19017), .I (I25114));
INVX1 gate8072(.O (I25117), .I (g18988));
INVX1 gate8073(.O (g19018), .I (I25117));
INVX1 gate8074(.O (I25120), .I (g18869));
INVX1 gate8075(.O (g19019), .I (I25120));
INVX1 gate8076(.O (I25123), .I (g18890));
INVX1 gate8077(.O (g19020), .I (I25123));
INVX1 gate8078(.O (I25126), .I (g16858));
INVX1 gate8079(.O (g19021), .I (I25126));
INVX1 gate8080(.O (I25129), .I (g16813));
INVX1 gate8081(.O (g19022), .I (I25129));
INVX1 gate8082(.O (I25132), .I (g16862));
INVX1 gate8083(.O (g19023), .I (I25132));
INVX1 gate8084(.O (I25135), .I (g16506));
INVX1 gate8085(.O (g19024), .I (I25135));
INVX1 gate8086(.O (I25138), .I (g18960));
INVX1 gate8087(.O (g19025), .I (I25138));
INVX1 gate8088(.O (I25141), .I (g18970));
INVX1 gate8089(.O (g19026), .I (I25141));
INVX1 gate8090(.O (I25144), .I (g18984));
INVX1 gate8091(.O (g19027), .I (I25144));
INVX1 gate8092(.O (I25147), .I (g18989));
INVX1 gate8093(.O (g19028), .I (I25147));
INVX1 gate8094(.O (I25150), .I (g18991));
INVX1 gate8095(.O (g19029), .I (I25150));
INVX1 gate8096(.O (I25153), .I (g18995));
INVX1 gate8097(.O (g19030), .I (I25153));
INVX1 gate8098(.O (I25156), .I (g18895));
INVX1 gate8099(.O (g19031), .I (I25156));
INVX1 gate8100(.O (I25159), .I (g18913));
INVX1 gate8101(.O (g19032), .I (I25159));
INVX1 gate8102(.O (I25162), .I (g16863));
INVX1 gate8103(.O (g19033), .I (I25162));
INVX1 gate8104(.O (I25165), .I (g16831));
INVX1 gate8105(.O (g19034), .I (I25165));
INVX1 gate8106(.O (I25168), .I (g16877));
INVX1 gate8107(.O (g19035), .I (I25168));
INVX1 gate8108(.O (I25171), .I (g16528));
INVX1 gate8109(.O (g19036), .I (I25171));
INVX1 gate8110(.O (I25174), .I (g18971));
INVX1 gate8111(.O (g19037), .I (I25174));
INVX1 gate8112(.O (I25177), .I (g18985));
INVX1 gate8113(.O (g19038), .I (I25177));
INVX1 gate8114(.O (I25180), .I (g18992));
INVX1 gate8115(.O (g19039), .I (I25180));
INVX1 gate8116(.O (I25183), .I (g18996));
INVX1 gate8117(.O (g19040), .I (I25183));
INVX1 gate8118(.O (I25186), .I (g18998));
INVX1 gate8119(.O (g19041), .I (I25186));
INVX1 gate8120(.O (I25189), .I (g19008));
INVX1 gate8121(.O (g19042), .I (I25189));
INVX1 gate8122(.O (I25192), .I (g18918));
INVX1 gate8123(.O (g19043), .I (I25192));
INVX1 gate8124(.O (I25195), .I (g18932));
INVX1 gate8125(.O (g19044), .I (I25195));
INVX1 gate8126(.O (I25198), .I (g16878));
INVX1 gate8127(.O (g19045), .I (I25198));
INVX1 gate8128(.O (I25201), .I (g16843));
INVX1 gate8129(.O (g19046), .I (I25201));
INVX1 gate8130(.O (I25204), .I (g16905));
INVX1 gate8131(.O (g19047), .I (I25204));
INVX1 gate8132(.O (I25207), .I (g16559));
INVX1 gate8133(.O (g19048), .I (I25207));
INVX1 gate8134(.O (I25210), .I (g18986));
INVX1 gate8135(.O (g19049), .I (I25210));
INVX1 gate8136(.O (I25213), .I (g18993));
INVX1 gate8137(.O (g19050), .I (I25213));
INVX1 gate8138(.O (I25216), .I (g18999));
INVX1 gate8139(.O (g19051), .I (I25216));
INVX1 gate8140(.O (I25219), .I (g19009));
INVX1 gate8141(.O (g19052), .I (I25219));
INVX1 gate8142(.O (I25222), .I (g19011));
INVX1 gate8143(.O (g19053), .I (I25222));
INVX1 gate8144(.O (I25225), .I (g16514));
INVX1 gate8145(.O (g19054), .I (I25225));
INVX1 gate8146(.O (I25228), .I (g18937));
INVX1 gate8147(.O (g19055), .I (I25228));
INVX1 gate8148(.O (I25231), .I (g18952));
INVX1 gate8149(.O (g19056), .I (I25231));
INVX1 gate8150(.O (I25234), .I (g16906));
INVX1 gate8151(.O (g19057), .I (I25234));
INVX1 gate8152(.O (I25237), .I (g16849));
INVX1 gate8153(.O (g19058), .I (I25237));
INVX1 gate8154(.O (I25240), .I (g16934));
INVX1 gate8155(.O (g19059), .I (I25240));
INVX1 gate8156(.O (I25243), .I (g17227));
INVX1 gate8157(.O (g19060), .I (I25243));
INVX1 gate8158(.O (I25246), .I (g17233));
INVX1 gate8159(.O (g19061), .I (I25246));
INVX1 gate8160(.O (I25249), .I (g17300));
INVX1 gate8161(.O (g19062), .I (I25249));
INVX1 gate8162(.O (I25253), .I (g17124));
INVX1 gate8163(.O (g19064), .I (I25253));
INVX1 gate8164(.O (g19070), .I (g18583));
INVX1 gate8165(.O (I25258), .I (g16974));
INVX1 gate8166(.O (g19075), .I (I25258));
INVX1 gate8167(.O (g19078), .I (g18619));
INVX1 gate8168(.O (I25264), .I (g17151));
INVX1 gate8169(.O (g19081), .I (I25264));
INVX1 gate8170(.O (I25272), .I (g17051));
INVX1 gate8171(.O (g19091), .I (I25272));
INVX1 gate8172(.O (g19096), .I (g18980));
INVX1 gate8173(.O (I25283), .I (g17086));
INVX1 gate8174(.O (g19098), .I (I25283));
INVX1 gate8175(.O (I25294), .I (g17124));
INVX1 gate8176(.O (g19105), .I (I25294));
INVX1 gate8177(.O (I25303), .I (g17151));
INVX1 gate8178(.O (g19110), .I (I25303));
INVX1 gate8179(.O (I25308), .I (g16867));
INVX1 gate8180(.O (g19113), .I (I25308));
INVX1 gate8181(.O (I25315), .I (g16895));
INVX1 gate8182(.O (g19118), .I (I25315));
INVX1 gate8183(.O (I25320), .I (g16924));
INVX1 gate8184(.O (g19125), .I (I25320));
INVX1 gate8185(.O (I25325), .I (g16954));
INVX1 gate8186(.O (g19132), .I (I25325));
INVX1 gate8187(.O (I25334), .I (g17645));
INVX1 gate8188(.O (g19145), .I (I25334));
INVX1 gate8189(.O (I25338), .I (g17746));
INVX1 gate8190(.O (g19147), .I (I25338));
INVX1 gate8191(.O (I25344), .I (g17847));
INVX1 gate8192(.O (g19151), .I (I25344));
INVX1 gate8193(.O (I25351), .I (g17959));
INVX1 gate8194(.O (g19156), .I (I25351));
INVX1 gate8195(.O (I25355), .I (g18669));
INVX1 gate8196(.O (g19158), .I (I25355));
INVX1 gate8197(.O (I25358), .I (g18678));
INVX1 gate8198(.O (g19159), .I (I25358));
INVX1 gate8199(.O (I25365), .I (g18707));
INVX1 gate8200(.O (g19164), .I (I25365));
INVX1 gate8201(.O (I25371), .I (g18719));
INVX1 gate8202(.O (g19168), .I (I25371));
INVX1 gate8203(.O (I25374), .I (g18726));
INVX1 gate8204(.O (g19169), .I (I25374));
INVX1 gate8205(.O (I25377), .I (g18743));
INVX1 gate8206(.O (g19170), .I (I25377));
INVX1 gate8207(.O (I25383), .I (g18755));
INVX1 gate8208(.O (g19174), .I (I25383));
INVX1 gate8209(.O (I25386), .I (g18763));
INVX1 gate8210(.O (g19175), .I (I25386));
INVX1 gate8211(.O (I25389), .I (g18780));
INVX1 gate8212(.O (g19176), .I (I25389));
INVX1 gate8213(.O (I25395), .I (g18782));
INVX1 gate8214(.O (g19180), .I (I25395));
INVX1 gate8215(.O (I25399), .I (g18794));
INVX1 gate8216(.O (g19182), .I (I25399));
INVX1 gate8217(.O (I25402), .I (g18821));
INVX1 gate8218(.O (g19183), .I (I25402));
INVX1 gate8219(.O (I25406), .I (g18804));
INVX1 gate8220(.O (g19185), .I (I25406));
INVX1 gate8221(.O (I25412), .I (g18820));
INVX1 gate8222(.O (g19189), .I (I25412));
INVX1 gate8223(.O (I25415), .I (g18835));
INVX1 gate8224(.O (g19190), .I (I25415));
INVX1 gate8225(.O (I25423), .I (g18852));
INVX1 gate8226(.O (g19196), .I (I25423));
INVX1 gate8227(.O (I25426), .I (g18836));
INVX1 gate8228(.O (g19197), .I (I25426));
INVX1 gate8229(.O (I25429), .I (g18975));
INVX1 gate8230(.O (g19198), .I (I25429));
INVX1 gate8231(.O (I25432), .I (g18837));
INVX1 gate8232(.O (g19199), .I (I25432));
INVX1 gate8233(.O (I25442), .I (g18866));
INVX1 gate8234(.O (g19207), .I (I25442));
INVX1 gate8235(.O (I25445), .I (g18968));
INVX1 gate8236(.O (g19208), .I (I25445));
INVX1 gate8237(.O (I25456), .I (g18883));
INVX1 gate8238(.O (g19217), .I (I25456));
INVX1 gate8239(.O (I25459), .I (g18867));
INVX1 gate8240(.O (g19218), .I (I25459));
INVX1 gate8241(.O (I25463), .I (g18868));
INVX1 gate8242(.O (g19220), .I (I25463));
INVX1 gate8243(.O (I25474), .I (g18885));
INVX1 gate8244(.O (g19229), .I (I25474));
INVX1 gate8245(.O (I25486), .I (g18754));
INVX1 gate8246(.O (g19237), .I (I25486));
INVX1 gate8247(.O (I25489), .I (g18906));
INVX1 gate8248(.O (g19238), .I (I25489));
INVX1 gate8249(.O (I25492), .I (g18907));
INVX1 gate8250(.O (g19239), .I (I25492));
INVX1 gate8251(.O (I25506), .I (g18781));
INVX1 gate8252(.O (g19247), .I (I25506));
INVX1 gate8253(.O (I25510), .I (g18542));
INVX1 gate8254(.O (g19249), .I (I25510));
INVX1 gate8255(.O (g19251), .I (g16540));
INVX1 gate8256(.O (I25525), .I (g18803));
INVX1 gate8257(.O (g19258), .I (I25525));
INVX1 gate8258(.O (I25528), .I (g18942));
INVX1 gate8259(.O (g19259), .I (I25528));
INVX1 gate8260(.O (g19265), .I (g16572));
INVX1 gate8261(.O (I25557), .I (g18957));
INVX1 gate8262(.O (g19270), .I (I25557));
INVX1 gate8263(.O (I25567), .I (g17186));
INVX1 gate8264(.O (g19272), .I (I25567));
INVX1 gate8265(.O (g19280), .I (g16596));
INVX1 gate8266(.O (g19287), .I (g16608));
INVX1 gate8267(.O (I25612), .I (g17197));
INVX1 gate8268(.O (g19291), .I (I25612));
INVX1 gate8269(.O (g19299), .I (g16616));
INVX1 gate8270(.O (g19301), .I (g16622));
INVX1 gate8271(.O (g19302), .I (g17025));
INVX1 gate8272(.O (g19305), .I (g16626));
INVX1 gate8273(.O (I25660), .I (g17204));
INVX1 gate8274(.O (g19309), .I (I25660));
INVX1 gate8275(.O (g19319), .I (g16633));
INVX1 gate8276(.O (g19322), .I (g16636));
INVX1 gate8277(.O (g19323), .I (g17059));
INVX1 gate8278(.O (g19326), .I (g16640));
INVX1 gate8279(.O (I25717), .I (g17209));
INVX1 gate8280(.O (g19330), .I (I25717));
INVX1 gate8281(.O (I25728), .I (g17118));
INVX1 gate8282(.O (g19335), .I (I25728));
INVX1 gate8283(.O (g19346), .I (g16644));
INVX1 gate8284(.O (g19349), .I (g16647));
INVX1 gate8285(.O (g19350), .I (g17094));
INVX1 gate8286(.O (g19353), .I (g16651));
INVX1 gate8287(.O (I25768), .I (g17139));
INVX1 gate8288(.O (g19358), .I (I25768));
INVX1 gate8289(.O (I25778), .I (g17145));
INVX1 gate8290(.O (g19369), .I (I25778));
INVX1 gate8291(.O (g19380), .I (g16656));
INVX1 gate8292(.O (g19383), .I (g16659));
INVX1 gate8293(.O (g19384), .I (g17132));
INVX1 gate8294(.O (g19387), .I (g16567));
INVX1 gate8295(.O (g19388), .I (g17139));
INVX1 gate8296(.O (I25816), .I (g17162));
INVX1 gate8297(.O (g19390), .I (I25816));
INVX1 gate8298(.O (I25826), .I (g17168));
INVX1 gate8299(.O (g19401), .I (I25826));
INVX1 gate8300(.O (g19412), .I (g16673));
INVX1 gate8301(.O (g19415), .I (g16676));
INVX1 gate8302(.O (g19417), .I (g16591));
INVX1 gate8303(.O (g19418), .I (g17162));
INVX1 gate8304(.O (I25862), .I (g17177));
INVX1 gate8305(.O (g19420), .I (I25862));
INVX1 gate8306(.O (I25872), .I (g17183));
INVX1 gate8307(.O (g19431), .I (I25872));
INVX1 gate8308(.O (g19441), .I (g17213));
INVX1 gate8309(.O (g19444), .I (g17985));
INVX1 gate8310(.O (g19448), .I (g16694));
INVX1 gate8311(.O (g19452), .I (g16702));
INVX1 gate8312(.O (g19454), .I (g16611));
INVX1 gate8313(.O (g19455), .I (g17177));
INVX1 gate8314(.O (I25904), .I (g17194));
INVX1 gate8315(.O (g19457), .I (I25904));
INVX1 gate8316(.O (g19467), .I (g16719));
INVX1 gate8317(.O (g19468), .I (g17216));
INVX1 gate8318(.O (g19471), .I (g18102));
INVX1 gate8319(.O (g19475), .I (g16725));
INVX1 gate8320(.O (g19479), .I (g16733));
INVX1 gate8321(.O (g19481), .I (g16629));
INVX1 gate8322(.O (g19482), .I (g17194));
INVX1 gate8323(.O (g19483), .I (g16758));
INVX1 gate8324(.O (g19484), .I (g16867));
INVX1 gate8325(.O (g19490), .I (g16761));
INVX1 gate8326(.O (g19491), .I (g17219));
INVX1 gate8327(.O (g19494), .I (g18218));
INVX1 gate8328(.O (g19498), .I (g16767));
INVX1 gate8329(.O (g19502), .I (g16775));
INVX1 gate8330(.O (g19504), .I (g16785));
INVX1 gate8331(.O (g19505), .I (g16895));
INVX1 gate8332(.O (g19511), .I (g16788));
INVX1 gate8333(.O (g19512), .I (g17221));
INVX1 gate8334(.O (g19515), .I (g18325));
INVX1 gate8335(.O (g19519), .I (g16794));
INVX1 gate8336(.O (g19523), .I (g16814));
INVX1 gate8337(.O (g19524), .I (g16924));
INVX1 gate8338(.O (g19530), .I (g16817));
INVX1 gate8339(.O (g19533), .I (g16832));
INVX1 gate8340(.O (g19534), .I (g16954));
INVX1 gate8341(.O (I25966), .I (g16654));
INVX1 gate8342(.O (g19543), .I (I25966));
INVX1 gate8343(.O (I25971), .I (g16671));
INVX1 gate8344(.O (g19546), .I (I25971));
INVX1 gate8345(.O (I25977), .I (g16692));
INVX1 gate8346(.O (g19550), .I (I25977));
INVX1 gate8347(.O (I25985), .I (g16718));
INVX1 gate8348(.O (g19556), .I (I25985));
INVX1 gate8349(.O (I25994), .I (g16860));
INVX1 gate8350(.O (g19563), .I (I25994));
INVX1 gate8351(.O (I26006), .I (g16866));
INVX1 gate8352(.O (g19573), .I (I26006));
INVX1 gate8353(.O (g19577), .I (g16881));
INVX1 gate8354(.O (g19578), .I (g16884));
INVX1 gate8355(.O (I26025), .I (g16803));
INVX1 gate8356(.O (g19595), .I (I26025));
INVX1 gate8357(.O (I26028), .I (g16566));
INVX1 gate8358(.O (g19596), .I (I26028));
INVX1 gate8359(.O (g19607), .I (g16910));
INVX1 gate8360(.O (g19608), .I (g16913));
INVX1 gate8361(.O (I26051), .I (g16824));
INVX1 gate8362(.O (g19622), .I (I26051));
INVX1 gate8363(.O (g19640), .I (g16940));
INVX1 gate8364(.O (g19641), .I (g16943));
INVX1 gate8365(.O (I26078), .I (g16835));
INVX1 gate8366(.O (g19652), .I (I26078));
INVX1 gate8367(.O (I26085), .I (g18085));
INVX1 gate8368(.O (g19657), .I (I26085));
INVX1 gate8369(.O (g19680), .I (g16971));
INVX1 gate8370(.O (g19681), .I (g16974));
INVX1 gate8371(.O (I26112), .I (g16844));
INVX1 gate8372(.O (g19689), .I (I26112));
INVX1 gate8373(.O (I26115), .I (g16845));
INVX1 gate8374(.O (g19690), .I (I26115));
INVX1 gate8375(.O (I26123), .I (g17503));
INVX1 gate8376(.O (g19696), .I (I26123));
INVX1 gate8377(.O (I26134), .I (g18201));
INVX1 gate8378(.O (g19705), .I (I26134));
INVX1 gate8379(.O (I26154), .I (g16851));
INVX1 gate8380(.O (g19725), .I (I26154));
INVX1 gate8381(.O (I26171), .I (g17594));
INVX1 gate8382(.O (g19740), .I (I26171));
INVX1 gate8383(.O (I26182), .I (g18308));
INVX1 gate8384(.O (g19749), .I (I26182));
INVX1 gate8385(.O (I26195), .I (g16853));
INVX1 gate8386(.O (g19762), .I (I26195));
INVX1 gate8387(.O (I26198), .I (g16854));
INVX1 gate8388(.O (g19763), .I (I26198));
INVX1 gate8389(.O (I26220), .I (g17691));
INVX1 gate8390(.O (g19783), .I (I26220));
INVX1 gate8391(.O (I26231), .I (g18401));
INVX1 gate8392(.O (g19792), .I (I26231));
INVX1 gate8393(.O (I26237), .I (g16857));
INVX1 gate8394(.O (g19798), .I (I26237));
INVX1 gate8395(.O (I26266), .I (g17791));
INVX1 gate8396(.O (g19825), .I (I26266));
INVX1 gate8397(.O (g19830), .I (g18886));
INVX1 gate8398(.O (I26276), .I (g16861));
INVX1 gate8399(.O (g19838), .I (I26276));
INVX1 gate8400(.O (I26334), .I (g18977));
INVX1 gate8401(.O (g19890), .I (I26334));
INVX1 gate8402(.O (I26337), .I (g16880));
INVX1 gate8403(.O (g19893), .I (I26337));
INVX1 gate8404(.O (I26340), .I (g17025));
INVX1 gate8405(.O (g19894), .I (I26340));
INVX1 gate8406(.O (I26365), .I (g18626));
INVX1 gate8407(.O (g19915), .I (I26365));
INVX1 gate8408(.O (g19918), .I (g18646));
INVX1 gate8409(.O (I26369), .I (g17059));
INVX1 gate8410(.O (g19919), .I (I26369));
INVX1 gate8411(.O (g19933), .I (g18548));
INVX1 gate8412(.O (I26388), .I (g17094));
INVX1 gate8413(.O (g19934), .I (I26388));
INVX1 gate8414(.O (I26401), .I (g17012));
INVX1 gate8415(.O (g19945), .I (I26401));
INVX1 gate8416(.O (g19948), .I (g17896));
INVX1 gate8417(.O (g19950), .I (g18598));
INVX1 gate8418(.O (I26407), .I (g17132));
INVX1 gate8419(.O (g19951), .I (I26407));
INVX1 gate8420(.O (I26413), .I (g16643));
INVX1 gate8421(.O (g19957), .I (I26413));
INVX1 gate8422(.O (I26420), .I (g17042));
INVX1 gate8423(.O (g19972), .I (I26420));
INVX1 gate8424(.O (g19975), .I (g18007));
INVX1 gate8425(.O (g19977), .I (g18630));
INVX1 gate8426(.O (I26426), .I (g16536));
INVX1 gate8427(.O (g19978), .I (I26426));
INVX1 gate8428(.O (I26437), .I (g16655));
INVX1 gate8429(.O (g19987), .I (I26437));
INVX1 gate8430(.O (I26444), .I (g17076));
INVX1 gate8431(.O (g20002), .I (I26444));
INVX1 gate8432(.O (g20005), .I (g18124));
INVX1 gate8433(.O (g20007), .I (g18639));
INVX1 gate8434(.O (I26458), .I (g17985));
INVX1 gate8435(.O (g20016), .I (I26458));
INVX1 gate8436(.O (I26469), .I (g16672));
INVX1 gate8437(.O (g20025), .I (I26469));
INVX1 gate8438(.O (I26476), .I (g17111));
INVX1 gate8439(.O (g20040), .I (I26476));
INVX1 gate8440(.O (g20043), .I (g18240));
INVX1 gate8441(.O (I26481), .I (g18590));
INVX1 gate8442(.O (g20045), .I (I26481));
INVX1 gate8443(.O (I26494), .I (g18102));
INVX1 gate8444(.O (g20058), .I (I26494));
INVX1 gate8445(.O (I26505), .I (g16693));
INVX1 gate8446(.O (g20067), .I (I26505));
INVX1 gate8447(.O (I26512), .I (g16802));
INVX1 gate8448(.O (g20082), .I (I26512));
INVX1 gate8449(.O (g20083), .I (g17968));
INVX1 gate8450(.O (I26535), .I (g18218));
INVX1 gate8451(.O (g20099), .I (I26535));
INVX1 gate8452(.O (I26545), .I (g16823));
INVX1 gate8453(.O (g20105), .I (I26545));
INVX1 gate8454(.O (I26574), .I (g18325));
INVX1 gate8455(.O (g20124), .I (I26574));
INVX1 gate8456(.O (g20127), .I (g18623));
INVX1 gate8457(.O (g20140), .I (g16830));
INVX1 gate8458(.O (g20163), .I (g17973));
INVX1 gate8459(.O (I26612), .I (g17645));
INVX1 gate8460(.O (g20164), .I (I26612));
INVX1 gate8461(.O (g20178), .I (g16842));
INVX1 gate8462(.O (g20193), .I (g18691));
INVX1 gate8463(.O (I26642), .I (g17746));
INVX1 gate8464(.O (g20198), .I (I26642));
INVX1 gate8465(.O (g20212), .I (g16848));
INVX1 gate8466(.O (g20223), .I (g18727));
INVX1 gate8467(.O (I26664), .I (g17847));
INVX1 gate8468(.O (g20228), .I (I26664));
INVX1 gate8469(.O (g20242), .I (g16852));
INVX1 gate8470(.O (g20250), .I (g18764));
INVX1 gate8471(.O (I26679), .I (g17959));
INVX1 gate8472(.O (g20255), .I (I26679));
INVX1 gate8473(.O (g20269), .I (g17230));
INVX1 gate8474(.O (g20273), .I (g18795));
INVX1 gate8475(.O (g20278), .I (g17237));
INVX1 gate8476(.O (g20279), .I (g17240));
INVX1 gate8477(.O (g20281), .I (g17243));
INVX1 gate8478(.O (g20286), .I (g17249));
INVX1 gate8479(.O (g20287), .I (g17252));
INVX1 gate8480(.O (g20288), .I (g17255));
INVX1 gate8481(.O (g20289), .I (g17259));
INVX1 gate8482(.O (g20290), .I (g17262));
INVX1 gate8483(.O (g20292), .I (g17265));
INVX1 gate8484(.O (I26714), .I (g17720));
INVX1 gate8485(.O (g20295), .I (I26714));
INVX1 gate8486(.O (g20296), .I (g17272));
INVX1 gate8487(.O (g20297), .I (g17275));
INVX1 gate8488(.O (g20298), .I (g17278));
INVX1 gate8489(.O (g20302), .I (g17282));
INVX1 gate8490(.O (g20303), .I (g17285));
INVX1 gate8491(.O (g20304), .I (g17288));
INVX1 gate8492(.O (g20305), .I (g17291));
INVX1 gate8493(.O (g20306), .I (g17294));
INVX1 gate8494(.O (g20308), .I (g17297));
INVX1 gate8495(.O (g20311), .I (g17304));
INVX1 gate8496(.O (g20312), .I (g17307));
INVX1 gate8497(.O (g20313), .I (g17310));
INVX1 gate8498(.O (g20315), .I (g17315));
INVX1 gate8499(.O (g20316), .I (g17318));
INVX1 gate8500(.O (g20317), .I (g17321));
INVX1 gate8501(.O (g20321), .I (g17324));
INVX1 gate8502(.O (g20322), .I (g17327));
INVX1 gate8503(.O (g20323), .I (g17330));
INVX1 gate8504(.O (g20324), .I (g17333));
INVX1 gate8505(.O (g20325), .I (g17336));
INVX1 gate8506(.O (g20327), .I (g17342));
INVX1 gate8507(.O (g20328), .I (g17345));
INVX1 gate8508(.O (g20329), .I (g17348));
INVX1 gate8509(.O (g20330), .I (g17354));
INVX1 gate8510(.O (g20331), .I (g17357));
INVX1 gate8511(.O (g20332), .I (g17360));
INVX1 gate8512(.O (g20334), .I (g17363));
INVX1 gate8513(.O (g20335), .I (g17366));
INVX1 gate8514(.O (g20336), .I (g17369));
INVX1 gate8515(.O (g20340), .I (g17372));
INVX1 gate8516(.O (g20341), .I (g17375));
INVX1 gate8517(.O (g20342), .I (g17378));
INVX1 gate8518(.O (g20344), .I (g17384));
INVX1 gate8519(.O (g20345), .I (g17387));
INVX1 gate8520(.O (g20346), .I (g17390));
INVX1 gate8521(.O (g20347), .I (g17399));
INVX1 gate8522(.O (g20348), .I (g17402));
INVX1 gate8523(.O (g20349), .I (g17405));
INVX1 gate8524(.O (g20350), .I (g17410));
INVX1 gate8525(.O (g20351), .I (g17413));
INVX1 gate8526(.O (g20352), .I (g17416));
INVX1 gate8527(.O (g20354), .I (g17419));
INVX1 gate8528(.O (g20355), .I (g17422));
INVX1 gate8529(.O (g20356), .I (g17425));
INVX1 gate8530(.O (I26777), .I (g17222));
INVX1 gate8531(.O (g20360), .I (I26777));
INVX1 gate8532(.O (g20361), .I (g17430));
INVX1 gate8533(.O (g20362), .I (g17433));
INVX1 gate8534(.O (g20363), .I (g17436));
INVX1 gate8535(.O (g20364), .I (g17439));
INVX1 gate8536(.O (g20365), .I (g17442));
INVX1 gate8537(.O (g20366), .I (g17451));
INVX1 gate8538(.O (g20367), .I (g17454));
INVX1 gate8539(.O (g20368), .I (g17457));
INVX1 gate8540(.O (g20369), .I (g17465));
INVX1 gate8541(.O (g20370), .I (g17468));
INVX1 gate8542(.O (g20371), .I (g17471));
INVX1 gate8543(.O (g20372), .I (g17476));
INVX1 gate8544(.O (g20373), .I (g17479));
INVX1 gate8545(.O (g20374), .I (g17482));
INVX1 gate8546(.O (I26796), .I (g17224));
INVX1 gate8547(.O (g20377), .I (I26796));
INVX1 gate8548(.O (g20378), .I (g17487));
INVX1 gate8549(.O (g20379), .I (g17490));
INVX1 gate8550(.O (g20380), .I (g17493));
INVX1 gate8551(.O (g20381), .I (g17496));
INVX1 gate8552(.O (g20382), .I (g17500));
INVX1 gate8553(.O (g20383), .I (g17503));
INVX1 gate8554(.O (g20384), .I (g17511));
INVX1 gate8555(.O (g20385), .I (g17514));
INVX1 gate8556(.O (g20386), .I (g17517));
INVX1 gate8557(.O (g20387), .I (g17520));
INVX1 gate8558(.O (g20388), .I (g17523));
INVX1 gate8559(.O (g20389), .I (g17531));
INVX1 gate8560(.O (g20390), .I (g17534));
INVX1 gate8561(.O (g20391), .I (g17537));
INVX1 gate8562(.O (g20392), .I (g17545));
INVX1 gate8563(.O (g20393), .I (g17548));
INVX1 gate8564(.O (g20394), .I (g17551));
INVX1 gate8565(.O (I26816), .I (g17225));
INVX1 gate8566(.O (g20395), .I (I26816));
INVX1 gate8567(.O (I26819), .I (g17226));
INVX1 gate8568(.O (g20396), .I (I26819));
INVX1 gate8569(.O (g20397), .I (g17557));
INVX1 gate8570(.O (g20398), .I (g17560));
INVX1 gate8571(.O (g20399), .I (g17563));
INVX1 gate8572(.O (g20400), .I (g17567));
INVX1 gate8573(.O (g20401), .I (g17570));
INVX1 gate8574(.O (g20402), .I (g17573));
INVX1 gate8575(.O (g20403), .I (g17579));
INVX1 gate8576(.O (g20404), .I (g17582));
INVX1 gate8577(.O (g20405), .I (g17585));
INVX1 gate8578(.O (g20406), .I (g17588));
INVX1 gate8579(.O (g20407), .I (g17591));
INVX1 gate8580(.O (g20408), .I (g17594));
INVX1 gate8581(.O (g20409), .I (g17601));
INVX1 gate8582(.O (g20410), .I (g17604));
INVX1 gate8583(.O (g20411), .I (g17607));
INVX1 gate8584(.O (g20412), .I (g17610));
INVX1 gate8585(.O (g20413), .I (g17613));
INVX1 gate8586(.O (g20414), .I (g17621));
INVX1 gate8587(.O (g20415), .I (g17624));
INVX1 gate8588(.O (g20416), .I (g17627));
INVX1 gate8589(.O (I26843), .I (g17228));
INVX1 gate8590(.O (g20418), .I (I26843));
INVX1 gate8591(.O (I26846), .I (g17229));
INVX1 gate8592(.O (g20419), .I (I26846));
INVX1 gate8593(.O (g20420), .I (g17637));
INVX1 gate8594(.O (g20421), .I (g17649));
INVX1 gate8595(.O (g20422), .I (g17655));
INVX1 gate8596(.O (g20423), .I (g17658));
INVX1 gate8597(.O (g20424), .I (g17661));
INVX1 gate8598(.O (g20425), .I (g17664));
INVX1 gate8599(.O (g20426), .I (g17667));
INVX1 gate8600(.O (g20427), .I (g17670));
INVX1 gate8601(.O (g20428), .I (g17676));
INVX1 gate8602(.O (g20429), .I (g17679));
INVX1 gate8603(.O (g20430), .I (g17682));
INVX1 gate8604(.O (g20431), .I (g17685));
INVX1 gate8605(.O (g20432), .I (g17688));
INVX1 gate8606(.O (g20433), .I (g17691));
INVX1 gate8607(.O (g20434), .I (g17698));
INVX1 gate8608(.O (g20435), .I (g17701));
INVX1 gate8609(.O (g20436), .I (g17704));
INVX1 gate8610(.O (g20437), .I (g17707));
INVX1 gate8611(.O (g20438), .I (g17710));
INVX1 gate8612(.O (I26868), .I (g17234));
INVX1 gate8613(.O (g20439), .I (I26868));
INVX1 gate8614(.O (I26871), .I (g17235));
INVX1 gate8615(.O (g20440), .I (I26871));
INVX1 gate8616(.O (I26874), .I (g17236));
INVX1 gate8617(.O (g20441), .I (I26874));
INVX1 gate8618(.O (g20442), .I (g17738));
INVX1 gate8619(.O (g20443), .I (g17749));
INVX1 gate8620(.O (g20444), .I (g17755));
INVX1 gate8621(.O (g20445), .I (g17758));
INVX1 gate8622(.O (g20446), .I (g17761));
INVX1 gate8623(.O (g20447), .I (g17764));
INVX1 gate8624(.O (g20448), .I (g17767));
INVX1 gate8625(.O (g20449), .I (g17770));
INVX1 gate8626(.O (g20450), .I (g17776));
INVX1 gate8627(.O (g20451), .I (g17779));
INVX1 gate8628(.O (g20452), .I (g17782));
INVX1 gate8629(.O (g20453), .I (g17785));
INVX1 gate8630(.O (g20454), .I (g17788));
INVX1 gate8631(.O (g20455), .I (g17791));
INVX1 gate8632(.O (g20456), .I (g17799));
INVX1 gate8633(.O (I26892), .I (g17246));
INVX1 gate8634(.O (g20457), .I (I26892));
INVX1 gate8635(.O (I26895), .I (g17247));
INVX1 gate8636(.O (g20458), .I (I26895));
INVX1 gate8637(.O (I26898), .I (g17248));
INVX1 gate8638(.O (g20459), .I (I26898));
INVX1 gate8639(.O (g20461), .I (g17839));
INVX1 gate8640(.O (g20462), .I (g17850));
INVX1 gate8641(.O (g20463), .I (g17856));
INVX1 gate8642(.O (g20464), .I (g17859));
INVX1 gate8643(.O (g20465), .I (g17862));
INVX1 gate8644(.O (g20466), .I (g17865));
INVX1 gate8645(.O (g20467), .I (g17868));
INVX1 gate8646(.O (g20468), .I (g17871));
INVX1 gate8647(.O (I26910), .I (g17269));
INVX1 gate8648(.O (g20469), .I (I26910));
INVX1 gate8649(.O (I26913), .I (g17270));
INVX1 gate8650(.O (g20470), .I (I26913));
INVX1 gate8651(.O (I26916), .I (g17271));
INVX1 gate8652(.O (g20471), .I (I26916));
INVX1 gate8653(.O (g20476), .I (g17951));
INVX1 gate8654(.O (g20477), .I (g17962));
INVX1 gate8655(.O (I26923), .I (g17302));
INVX1 gate8656(.O (g20478), .I (I26923));
INVX1 gate8657(.O (I26926), .I (g17303));
INVX1 gate8658(.O (g20479), .I (I26926));
INVX1 gate8659(.O (I26931), .I (g17340));
INVX1 gate8660(.O (g20484), .I (I26931));
INVX1 gate8661(.O (I26934), .I (g17341));
INVX1 gate8662(.O (g20485), .I (I26934));
INVX1 gate8663(.O (g20490), .I (g18166));
INVX1 gate8664(.O (I26940), .I (g17383));
INVX1 gate8665(.O (g20491), .I (I26940));
INVX1 gate8666(.O (g20496), .I (g18258));
INVX1 gate8667(.O (I26947), .I (g17429));
INVX1 gate8668(.O (g20498), .I (I26947));
INVX1 gate8669(.O (g20500), .I (g18278));
INVX1 gate8670(.O (g20501), .I (g18334));
INVX1 gate8671(.O (g20504), .I (g18355));
INVX1 gate8672(.O (g20505), .I (g18371));
INVX1 gate8673(.O (g20507), .I (g18351));
INVX1 gate8674(.O (I26960), .I (g16884));
INVX1 gate8675(.O (g20513), .I (I26960));
INVX1 gate8676(.O (g20516), .I (g18432));
INVX1 gate8677(.O (g20517), .I (g18450));
INVX1 gate8678(.O (g20518), .I (g18466));
INVX1 gate8679(.O (I26966), .I (g17051));
INVX1 gate8680(.O (g20519), .I (I26966));
INVX1 gate8681(.O (g20526), .I (g18446));
INVX1 gate8682(.O (I26972), .I (g16913));
INVX1 gate8683(.O (g20531), .I (I26972));
INVX1 gate8684(.O (g20534), .I (g18505));
INVX1 gate8685(.O (g20535), .I (g18523));
INVX1 gate8686(.O (g20536), .I (g18539));
INVX1 gate8687(.O (I26980), .I (g17086));
INVX1 gate8688(.O (g20539), .I (I26980));
INVX1 gate8689(.O (g20545), .I (g18519));
INVX1 gate8690(.O (I26985), .I (g16943));
INVX1 gate8691(.O (g20550), .I (I26985));
INVX1 gate8692(.O (g20553), .I (g18569));
INVX1 gate8693(.O (g20554), .I (g18587));
INVX1 gate8694(.O (I26990), .I (g19145));
INVX1 gate8695(.O (g20555), .I (I26990));
INVX1 gate8696(.O (I26993), .I (g19159));
INVX1 gate8697(.O (g20556), .I (I26993));
INVX1 gate8698(.O (I26996), .I (g19169));
INVX1 gate8699(.O (g20557), .I (I26996));
INVX1 gate8700(.O (I26999), .I (g19543));
INVX1 gate8701(.O (g20558), .I (I26999));
INVX1 gate8702(.O (I27002), .I (g19147));
INVX1 gate8703(.O (g20559), .I (I27002));
INVX1 gate8704(.O (I27005), .I (g19164));
INVX1 gate8705(.O (g20560), .I (I27005));
INVX1 gate8706(.O (I27008), .I (g19175));
INVX1 gate8707(.O (g20561), .I (I27008));
INVX1 gate8708(.O (I27011), .I (g19546));
INVX1 gate8709(.O (g20562), .I (I27011));
INVX1 gate8710(.O (I27014), .I (g19151));
INVX1 gate8711(.O (g20563), .I (I27014));
INVX1 gate8712(.O (I27017), .I (g19170));
INVX1 gate8713(.O (g20564), .I (I27017));
INVX1 gate8714(.O (I27020), .I (g19182));
INVX1 gate8715(.O (g20565), .I (I27020));
INVX1 gate8716(.O (I27023), .I (g19550));
INVX1 gate8717(.O (g20566), .I (I27023));
INVX1 gate8718(.O (I27026), .I (g19156));
INVX1 gate8719(.O (g20567), .I (I27026));
INVX1 gate8720(.O (I27029), .I (g19176));
INVX1 gate8721(.O (g20568), .I (I27029));
INVX1 gate8722(.O (I27032), .I (g19189));
INVX1 gate8723(.O (g20569), .I (I27032));
INVX1 gate8724(.O (I27035), .I (g19556));
INVX1 gate8725(.O (g20570), .I (I27035));
INVX1 gate8726(.O (I27038), .I (g20082));
INVX1 gate8727(.O (g20571), .I (I27038));
INVX1 gate8728(.O (I27041), .I (g19237));
INVX1 gate8729(.O (g20572), .I (I27041));
INVX1 gate8730(.O (I27044), .I (g19247));
INVX1 gate8731(.O (g20573), .I (I27044));
INVX1 gate8732(.O (I27047), .I (g19258));
INVX1 gate8733(.O (g20574), .I (I27047));
INVX1 gate8734(.O (I27050), .I (g19183));
INVX1 gate8735(.O (g20575), .I (I27050));
INVX1 gate8736(.O (I27053), .I (g19190));
INVX1 gate8737(.O (g20576), .I (I27053));
INVX1 gate8738(.O (I27056), .I (g19196));
INVX1 gate8739(.O (g20577), .I (I27056));
INVX1 gate8740(.O (I27059), .I (g19207));
INVX1 gate8741(.O (g20578), .I (I27059));
INVX1 gate8742(.O (I27062), .I (g19217));
INVX1 gate8743(.O (g20579), .I (I27062));
INVX1 gate8744(.O (I27065), .I (g19270));
INVX1 gate8745(.O (g20580), .I (I27065));
INVX1 gate8746(.O (I27068), .I (g19197));
INVX1 gate8747(.O (g20581), .I (I27068));
INVX1 gate8748(.O (I27071), .I (g19218));
INVX1 gate8749(.O (g20582), .I (I27071));
INVX1 gate8750(.O (I27074), .I (g19238));
INVX1 gate8751(.O (g20583), .I (I27074));
INVX1 gate8752(.O (I27077), .I (g19259));
INVX1 gate8753(.O (g20584), .I (I27077));
INVX1 gate8754(.O (I27080), .I (g19198));
INVX1 gate8755(.O (g20585), .I (I27080));
INVX1 gate8756(.O (I27083), .I (g19208));
INVX1 gate8757(.O (g20586), .I (I27083));
INVX1 gate8758(.O (I27086), .I (g19229));
INVX1 gate8759(.O (g20587), .I (I27086));
INVX1 gate8760(.O (I27089), .I (g20105));
INVX1 gate8761(.O (g20588), .I (I27089));
INVX1 gate8762(.O (I27092), .I (g19174));
INVX1 gate8763(.O (g20589), .I (I27092));
INVX1 gate8764(.O (I27095), .I (g19185));
INVX1 gate8765(.O (g20590), .I (I27095));
INVX1 gate8766(.O (I27098), .I (g19199));
INVX1 gate8767(.O (g20591), .I (I27098));
INVX1 gate8768(.O (I27101), .I (g19220));
INVX1 gate8769(.O (g20592), .I (I27101));
INVX1 gate8770(.O (I27104), .I (g19239));
INVX1 gate8771(.O (g20593), .I (I27104));
INVX1 gate8772(.O (I27107), .I (g19249));
INVX1 gate8773(.O (g20594), .I (I27107));
INVX1 gate8774(.O (I27110), .I (g19622));
INVX1 gate8775(.O (g20595), .I (I27110));
INVX1 gate8776(.O (I27113), .I (g19689));
INVX1 gate8777(.O (g20596), .I (I27113));
INVX1 gate8778(.O (I27116), .I (g19762));
INVX1 gate8779(.O (g20597), .I (I27116));
INVX1 gate8780(.O (I27119), .I (g19563));
INVX1 gate8781(.O (g20598), .I (I27119));
INVX1 gate8782(.O (I27122), .I (g19595));
INVX1 gate8783(.O (g20599), .I (I27122));
INVX1 gate8784(.O (I27125), .I (g19652));
INVX1 gate8785(.O (g20600), .I (I27125));
INVX1 gate8786(.O (I27128), .I (g19725));
INVX1 gate8787(.O (g20601), .I (I27128));
INVX1 gate8788(.O (I27131), .I (g19798));
INVX1 gate8789(.O (g20602), .I (I27131));
INVX1 gate8790(.O (I27134), .I (g19573));
INVX1 gate8791(.O (g20603), .I (I27134));
INVX1 gate8792(.O (I27137), .I (g19596));
INVX1 gate8793(.O (g20604), .I (I27137));
INVX1 gate8794(.O (I27140), .I (g19690));
INVX1 gate8795(.O (g20605), .I (I27140));
INVX1 gate8796(.O (I27143), .I (g19763));
INVX1 gate8797(.O (g20606), .I (I27143));
INVX1 gate8798(.O (I27146), .I (g19838));
INVX1 gate8799(.O (g20607), .I (I27146));
INVX1 gate8800(.O (I27149), .I (g19893));
INVX1 gate8801(.O (g20608), .I (I27149));
INVX1 gate8802(.O (I27152), .I (g20360));
INVX1 gate8803(.O (g20609), .I (I27152));
INVX1 gate8804(.O (I27155), .I (g20395));
INVX1 gate8805(.O (g20610), .I (I27155));
INVX1 gate8806(.O (I27158), .I (g20439));
INVX1 gate8807(.O (g20611), .I (I27158));
INVX1 gate8808(.O (I27161), .I (g20377));
INVX1 gate8809(.O (g20612), .I (I27161));
INVX1 gate8810(.O (I27164), .I (g20418));
INVX1 gate8811(.O (g20613), .I (I27164));
INVX1 gate8812(.O (I27167), .I (g20457));
INVX1 gate8813(.O (g20614), .I (I27167));
INVX1 gate8814(.O (I27170), .I (g20396));
INVX1 gate8815(.O (g20615), .I (I27170));
INVX1 gate8816(.O (I27173), .I (g20440));
INVX1 gate8817(.O (g20616), .I (I27173));
INVX1 gate8818(.O (I27176), .I (g20469));
INVX1 gate8819(.O (g20617), .I (I27176));
INVX1 gate8820(.O (I27179), .I (g20419));
INVX1 gate8821(.O (g20618), .I (I27179));
INVX1 gate8822(.O (I27182), .I (g20458));
INVX1 gate8823(.O (g20619), .I (I27182));
INVX1 gate8824(.O (I27185), .I (g20478));
INVX1 gate8825(.O (g20620), .I (I27185));
INVX1 gate8826(.O (I27188), .I (g20441));
INVX1 gate8827(.O (g20621), .I (I27188));
INVX1 gate8828(.O (I27191), .I (g20470));
INVX1 gate8829(.O (g20622), .I (I27191));
INVX1 gate8830(.O (I27194), .I (g20484));
INVX1 gate8831(.O (g20623), .I (I27194));
INVX1 gate8832(.O (I27197), .I (g20459));
INVX1 gate8833(.O (g20624), .I (I27197));
INVX1 gate8834(.O (I27200), .I (g20479));
INVX1 gate8835(.O (g20625), .I (I27200));
INVX1 gate8836(.O (I27203), .I (g20491));
INVX1 gate8837(.O (g20626), .I (I27203));
INVX1 gate8838(.O (I27206), .I (g20471));
INVX1 gate8839(.O (g20627), .I (I27206));
INVX1 gate8840(.O (I27209), .I (g20485));
INVX1 gate8841(.O (g20628), .I (I27209));
INVX1 gate8842(.O (I27212), .I (g20498));
INVX1 gate8843(.O (g20629), .I (I27212));
INVX1 gate8844(.O (I27215), .I (g19158));
INVX1 gate8845(.O (g20630), .I (I27215));
INVX1 gate8846(.O (I27218), .I (g19168));
INVX1 gate8847(.O (g20631), .I (I27218));
INVX1 gate8848(.O (I27221), .I (g19180));
INVX1 gate8849(.O (g20632), .I (I27221));
INVX1 gate8850(.O (I27225), .I (g19358));
INVX1 gate8851(.O (g20634), .I (I27225));
INVX1 gate8852(.O (I27228), .I (g19390));
INVX1 gate8853(.O (g20637), .I (I27228));
INVX1 gate8854(.O (I27232), .I (g19401));
INVX1 gate8855(.O (g20641), .I (I27232));
INVX1 gate8856(.O (I27235), .I (g19420));
INVX1 gate8857(.O (g20644), .I (I27235));
INVX1 gate8858(.O (I27240), .I (g19335));
INVX1 gate8859(.O (g20649), .I (I27240));
INVX1 gate8860(.O (I27243), .I (g19335));
INVX1 gate8861(.O (g20652), .I (I27243));
INVX1 gate8862(.O (I27246), .I (g19335));
INVX1 gate8863(.O (g20655), .I (I27246));
INVX1 gate8864(.O (I27250), .I (g19390));
INVX1 gate8865(.O (g20659), .I (I27250));
INVX1 gate8866(.O (I27253), .I (g19420));
INVX1 gate8867(.O (g20662), .I (I27253));
INVX1 gate8868(.O (I27257), .I (g19431));
INVX1 gate8869(.O (g20666), .I (I27257));
INVX1 gate8870(.O (I27260), .I (g19457));
INVX1 gate8871(.O (g20669), .I (I27260));
INVX1 gate8872(.O (I27264), .I (g19358));
INVX1 gate8873(.O (g20673), .I (I27264));
INVX1 gate8874(.O (I27267), .I (g19358));
INVX1 gate8875(.O (g20676), .I (I27267));
INVX1 gate8876(.O (I27270), .I (g19335));
INVX1 gate8877(.O (g20679), .I (I27270));
INVX1 gate8878(.O (I27275), .I (g19369));
INVX1 gate8879(.O (g20684), .I (I27275));
INVX1 gate8880(.O (I27278), .I (g19369));
INVX1 gate8881(.O (g20687), .I (I27278));
INVX1 gate8882(.O (I27281), .I (g19369));
INVX1 gate8883(.O (g20690), .I (I27281));
INVX1 gate8884(.O (I27285), .I (g19420));
INVX1 gate8885(.O (g20694), .I (I27285));
INVX1 gate8886(.O (I27288), .I (g19457));
INVX1 gate8887(.O (g20697), .I (I27288));
INVX1 gate8888(.O (I27293), .I (g19335));
INVX1 gate8889(.O (g20704), .I (I27293));
INVX1 gate8890(.O (I27297), .I (g19390));
INVX1 gate8891(.O (g20708), .I (I27297));
INVX1 gate8892(.O (I27300), .I (g19390));
INVX1 gate8893(.O (g20711), .I (I27300));
INVX1 gate8894(.O (I27303), .I (g19369));
INVX1 gate8895(.O (g20714), .I (I27303));
INVX1 gate8896(.O (I27308), .I (g19401));
INVX1 gate8897(.O (g20719), .I (I27308));
INVX1 gate8898(.O (I27311), .I (g19401));
INVX1 gate8899(.O (g20722), .I (I27311));
INVX1 gate8900(.O (I27314), .I (g19401));
INVX1 gate8901(.O (g20725), .I (I27314));
INVX1 gate8902(.O (I27318), .I (g19457));
INVX1 gate8903(.O (g20729), .I (I27318));
INVX1 gate8904(.O (I27321), .I (g19335));
INVX1 gate8905(.O (g20732), .I (I27321));
INVX1 gate8906(.O (I27324), .I (g19358));
INVX1 gate8907(.O (g20735), .I (I27324));
INVX1 gate8908(.O (I27328), .I (g19369));
INVX1 gate8909(.O (g20739), .I (I27328));
INVX1 gate8910(.O (I27332), .I (g19420));
INVX1 gate8911(.O (g20743), .I (I27332));
INVX1 gate8912(.O (I27335), .I (g19420));
INVX1 gate8913(.O (g20746), .I (I27335));
INVX1 gate8914(.O (I27338), .I (g19401));
INVX1 gate8915(.O (g20749), .I (I27338));
INVX1 gate8916(.O (I27343), .I (g19431));
INVX1 gate8917(.O (g20754), .I (I27343));
INVX1 gate8918(.O (I27346), .I (g19431));
INVX1 gate8919(.O (g20757), .I (I27346));
INVX1 gate8920(.O (I27349), .I (g19431));
INVX1 gate8921(.O (g20760), .I (I27349));
INVX1 gate8922(.O (I27352), .I (g19358));
INVX1 gate8923(.O (g20763), .I (I27352));
INVX1 gate8924(.O (I27355), .I (g19335));
INVX1 gate8925(.O (g20766), .I (I27355));
INVX1 gate8926(.O (I27358), .I (g19369));
INVX1 gate8927(.O (g20769), .I (I27358));
INVX1 gate8928(.O (I27361), .I (g19390));
INVX1 gate8929(.O (g20772), .I (I27361));
INVX1 gate8930(.O (I27365), .I (g19401));
INVX1 gate8931(.O (g20776), .I (I27365));
INVX1 gate8932(.O (I27369), .I (g19457));
INVX1 gate8933(.O (g20780), .I (I27369));
INVX1 gate8934(.O (I27372), .I (g19457));
INVX1 gate8935(.O (g20783), .I (I27372));
INVX1 gate8936(.O (I27375), .I (g19431));
INVX1 gate8937(.O (g20786), .I (I27375));
INVX1 gate8938(.O (I27379), .I (g19358));
INVX1 gate8939(.O (g20790), .I (I27379));
INVX1 gate8940(.O (I27382), .I (g19390));
INVX1 gate8941(.O (g20793), .I (I27382));
INVX1 gate8942(.O (I27385), .I (g19369));
INVX1 gate8943(.O (g20796), .I (I27385));
INVX1 gate8944(.O (I27388), .I (g19401));
INVX1 gate8945(.O (g20799), .I (I27388));
INVX1 gate8946(.O (I27391), .I (g19420));
INVX1 gate8947(.O (g20802), .I (I27391));
INVX1 gate8948(.O (I27395), .I (g19431));
INVX1 gate8949(.O (g20806), .I (I27395));
INVX1 gate8950(.O (I27399), .I (g19390));
INVX1 gate8951(.O (g20810), .I (I27399));
INVX1 gate8952(.O (I27402), .I (g19420));
INVX1 gate8953(.O (g20813), .I (I27402));
INVX1 gate8954(.O (I27405), .I (g19401));
INVX1 gate8955(.O (g20816), .I (I27405));
INVX1 gate8956(.O (I27408), .I (g19431));
INVX1 gate8957(.O (g20819), .I (I27408));
INVX1 gate8958(.O (I27411), .I (g19457));
INVX1 gate8959(.O (g20822), .I (I27411));
INVX1 gate8960(.O (I27416), .I (g19420));
INVX1 gate8961(.O (g20827), .I (I27416));
INVX1 gate8962(.O (I27419), .I (g19457));
INVX1 gate8963(.O (g20830), .I (I27419));
INVX1 gate8964(.O (I27422), .I (g19431));
INVX1 gate8965(.O (g20833), .I (I27422));
INVX1 gate8966(.O (I27426), .I (g19457));
INVX1 gate8967(.O (g20837), .I (I27426));
INVX1 gate8968(.O (g20842), .I (g19441));
INVX1 gate8969(.O (g20850), .I (g19468));
INVX1 gate8970(.O (g20858), .I (g19491));
INVX1 gate8971(.O (g20866), .I (g19512));
INVX1 gate8972(.O (g20885), .I (g19865));
INVX1 gate8973(.O (g20904), .I (g19896));
INVX1 gate8974(.O (g20928), .I (g19921));
INVX1 gate8975(.O (I27488), .I (g20310));
INVX1 gate8976(.O (g20942), .I (I27488));
INVX1 gate8977(.O (I27491), .I (g20314));
INVX1 gate8978(.O (g20943), .I (I27491));
INVX1 gate8979(.O (g20956), .I (g19936));
INVX1 gate8980(.O (I27516), .I (g20333));
INVX1 gate8981(.O (g20971), .I (I27516));
INVX1 gate8982(.O (I27531), .I (g20343));
INVX1 gate8983(.O (g20984), .I (I27531));
INVX1 gate8984(.O (I27534), .I (g20083));
INVX1 gate8985(.O (g20985), .I (I27534));
INVX1 gate8986(.O (I27537), .I (g19957));
INVX1 gate8987(.O (g20986), .I (I27537));
INVX1 gate8988(.O (I27549), .I (g20353));
INVX1 gate8989(.O (g20998), .I (I27549));
INVX1 gate8990(.O (I27565), .I (g19987));
INVX1 gate8991(.O (g21012), .I (I27565));
INVX1 gate8992(.O (I27577), .I (g20375));
INVX1 gate8993(.O (g21024), .I (I27577));
INVX1 gate8994(.O (I27585), .I (g20376));
INVX1 gate8995(.O (g21030), .I (I27585));
INVX1 gate8996(.O (I27593), .I (g20025));
INVX1 gate8997(.O (g21036), .I (I27593));
INVX1 gate8998(.O (g21050), .I (g20513));
INVX1 gate8999(.O (I27614), .I (g20067));
INVX1 gate9000(.O (g21057), .I (I27614));
INVX1 gate9001(.O (I27621), .I (g20417));
INVX1 gate9002(.O (g21064), .I (I27621));
INVX1 gate9003(.O (g21066), .I (g20519));
INVX1 gate9004(.O (g21069), .I (g20531));
INVX1 gate9005(.O (g21076), .I (g20539));
INVX1 gate9006(.O (g21079), .I (g20550));
INVX1 gate9007(.O (I27646), .I (g20507));
INVX1 gate9008(.O (g21087), .I (I27646));
INVX1 gate9009(.O (g21090), .I (g19064));
INVX1 gate9010(.O (g21093), .I (g19075));
INVX1 gate9011(.O (I27658), .I (g20526));
INVX1 gate9012(.O (g21099), .I (I27658));
INVX1 gate9013(.O (g21102), .I (g19081));
INVX1 gate9014(.O (I27667), .I (g20507));
INVX1 gate9015(.O (g21108), .I (I27667));
INVX1 gate9016(.O (I27672), .I (g20545));
INVX1 gate9017(.O (g21113), .I (I27672));
INVX1 gate9018(.O (I27684), .I (g20526));
INVX1 gate9019(.O (g21125), .I (I27684));
INVX1 gate9020(.O (I27689), .I (g19070));
INVX1 gate9021(.O (g21130), .I (I27689));
INVX1 gate9022(.O (I27705), .I (g20545));
INVX1 gate9023(.O (g21144), .I (I27705));
INVX1 gate9024(.O (I27727), .I (g19070));
INVX1 gate9025(.O (g21164), .I (I27727));
INVX1 gate9026(.O (I27749), .I (g19954));
INVX1 gate9027(.O (g21184), .I (I27749));
INVX1 gate9028(.O (g21187), .I (g19113));
INVX1 gate9029(.O (I27766), .I (g19984));
INVX1 gate9030(.O (g21199), .I (I27766));
INVX1 gate9031(.O (g21202), .I (g19118));
INVX1 gate9032(.O (I27779), .I (g20022));
INVX1 gate9033(.O (g21214), .I (I27779));
INVX1 gate9034(.O (g21217), .I (g19125));
INVX1 gate9035(.O (I27785), .I (g20064));
INVX1 gate9036(.O (g21222), .I (I27785));
INVX1 gate9037(.O (g21225), .I (g19132));
INVX1 gate9038(.O (g21241), .I (g19945));
INVX1 gate9039(.O (g21249), .I (g19972));
INVX1 gate9040(.O (g21258), .I (g20002));
INVX1 gate9041(.O (g21266), .I (g20040));
INVX1 gate9042(.O (I27822), .I (g19865));
INVX1 gate9043(.O (g21271), .I (I27822));
INVX1 gate9044(.O (I27827), .I (g19896));
INVX1 gate9045(.O (g21278), .I (I27827));
INVX1 gate9046(.O (I27832), .I (g19921));
INVX1 gate9047(.O (g21285), .I (I27832));
INVX1 gate9048(.O (I27838), .I (g19936));
INVX1 gate9049(.O (g21293), .I (I27838));
INVX1 gate9050(.O (I27868), .I (g19144));
INVX1 gate9051(.O (g21327), .I (I27868));
INVX1 gate9052(.O (I27897), .I (g19149));
INVX1 gate9053(.O (g21358), .I (I27897));
INVX1 gate9054(.O (I27900), .I (g19096));
INVX1 gate9055(.O (g21359), .I (I27900));
INVX1 gate9056(.O (I27917), .I (g19153));
INVX1 gate9057(.O (g21376), .I (I27917));
INVX1 gate9058(.O (I27920), .I (g19154));
INVX1 gate9059(.O (g21377), .I (I27920));
INVX1 gate9060(.O (I27927), .I (g19957));
INVX1 gate9061(.O (g21382), .I (I27927));
INVX1 gate9062(.O (I27942), .I (g19157));
INVX1 gate9063(.O (g21399), .I (I27942));
INVX1 gate9064(.O (g21400), .I (g19918));
INVX1 gate9065(.O (I27949), .I (g19957));
INVX1 gate9066(.O (g21404), .I (I27949));
INVX1 gate9067(.O (I27958), .I (g19987));
INVX1 gate9068(.O (g21415), .I (I27958));
INVX1 gate9069(.O (I27969), .I (g19162));
INVX1 gate9070(.O (g21426), .I (I27969));
INVX1 gate9071(.O (I27972), .I (g19163));
INVX1 gate9072(.O (g21427), .I (I27972));
INVX1 gate9073(.O (I27976), .I (g19957));
INVX1 gate9074(.O (g21429), .I (I27976));
INVX1 gate9075(.O (I27984), .I (g19987));
INVX1 gate9076(.O (g21441), .I (I27984));
INVX1 gate9077(.O (I27992), .I (g20025));
INVX1 gate9078(.O (g21449), .I (I27992));
INVX1 gate9079(.O (I28000), .I (g19167));
INVX1 gate9080(.O (g21457), .I (I28000));
INVX1 gate9081(.O (I28003), .I (g19957));
INVX1 gate9082(.O (g21458), .I (I28003));
INVX1 gate9083(.O (g21461), .I (g19957));
INVX1 gate9084(.O (I28009), .I (g20473));
INVX1 gate9085(.O (g21473), .I (I28009));
INVX1 gate9086(.O (I28013), .I (g19987));
INVX1 gate9087(.O (g21477), .I (I28013));
INVX1 gate9088(.O (I28019), .I (g20025));
INVX1 gate9089(.O (g21483), .I (I28019));
INVX1 gate9090(.O (I28027), .I (g20067));
INVX1 gate9091(.O (g21491), .I (I28027));
INVX1 gate9092(.O (I28031), .I (g19172));
INVX1 gate9093(.O (g21495), .I (I28031));
INVX1 gate9094(.O (I28034), .I (g19173));
INVX1 gate9095(.O (g21496), .I (I28034));
INVX1 gate9096(.O (I28038), .I (g19957));
INVX1 gate9097(.O (g21498), .I (I28038));
INVX1 gate9098(.O (I28043), .I (g19987));
INVX1 gate9099(.O (g21505), .I (I28043));
INVX1 gate9100(.O (g21508), .I (g19987));
INVX1 gate9101(.O (I28047), .I (g20481));
INVX1 gate9102(.O (g21514), .I (I28047));
INVX1 gate9103(.O (I28051), .I (g20025));
INVX1 gate9104(.O (g21518), .I (I28051));
INVX1 gate9105(.O (I28057), .I (g20067));
INVX1 gate9106(.O (g21524), .I (I28057));
INVX1 gate9107(.O (I28061), .I (g19178));
INVX1 gate9108(.O (g21528), .I (I28061));
INVX1 gate9109(.O (g21529), .I (g19272));
INVX1 gate9110(.O (I28065), .I (g19957));
INVX1 gate9111(.O (g21530), .I (I28065));
INVX1 gate9112(.O (I28072), .I (g19987));
INVX1 gate9113(.O (g21537), .I (I28072));
INVX1 gate9114(.O (I28076), .I (g20025));
INVX1 gate9115(.O (g21541), .I (I28076));
INVX1 gate9116(.O (g21544), .I (g20025));
INVX1 gate9117(.O (I28080), .I (g20487));
INVX1 gate9118(.O (g21550), .I (I28080));
INVX1 gate9119(.O (I28084), .I (g20067));
INVX1 gate9120(.O (g21554), .I (I28084));
INVX1 gate9121(.O (I28087), .I (g19184));
INVX1 gate9122(.O (g21557), .I (I28087));
INVX1 gate9123(.O (I28090), .I (g20008));
INVX1 gate9124(.O (g21558), .I (I28090));
INVX1 gate9125(.O (I28093), .I (g19957));
INVX1 gate9126(.O (g21561), .I (I28093));
INVX1 gate9127(.O (g21565), .I (g19291));
INVX1 gate9128(.O (I28100), .I (g19987));
INVX1 gate9129(.O (g21566), .I (I28100));
INVX1 gate9130(.O (I28107), .I (g20025));
INVX1 gate9131(.O (g21573), .I (I28107));
INVX1 gate9132(.O (I28111), .I (g20067));
INVX1 gate9133(.O (g21577), .I (I28111));
INVX1 gate9134(.O (g21580), .I (g20067));
INVX1 gate9135(.O (I28115), .I (g20493));
INVX1 gate9136(.O (g21586), .I (I28115));
INVX1 gate9137(.O (I28119), .I (g19957));
INVX1 gate9138(.O (g21590), .I (I28119));
INVX1 gate9139(.O (I28123), .I (g19987));
INVX1 gate9140(.O (g21594), .I (I28123));
INVX1 gate9141(.O (g21598), .I (g19309));
INVX1 gate9142(.O (I28130), .I (g20025));
INVX1 gate9143(.O (g21599), .I (I28130));
INVX1 gate9144(.O (I28137), .I (g20067));
INVX1 gate9145(.O (g21606), .I (I28137));
INVX1 gate9146(.O (I28143), .I (g19957));
INVX1 gate9147(.O (g21612), .I (I28143));
INVX1 gate9148(.O (I28148), .I (g19987));
INVX1 gate9149(.O (g21619), .I (I28148));
INVX1 gate9150(.O (I28152), .I (g20025));
INVX1 gate9151(.O (g21623), .I (I28152));
INVX1 gate9152(.O (g21627), .I (g19330));
INVX1 gate9153(.O (I28159), .I (g20067));
INVX1 gate9154(.O (g21628), .I (I28159));
INVX1 gate9155(.O (I28169), .I (g19987));
INVX1 gate9156(.O (g21640), .I (I28169));
INVX1 gate9157(.O (I28174), .I (g20025));
INVX1 gate9158(.O (g21647), .I (I28174));
INVX1 gate9159(.O (I28178), .I (g20067));
INVX1 gate9160(.O (g21651), .I (I28178));
INVX1 gate9161(.O (I28184), .I (g19103));
INVX1 gate9162(.O (g21655), .I (I28184));
INVX1 gate9163(.O (g21661), .I (g19091));
INVX1 gate9164(.O (I28201), .I (g20025));
INVX1 gate9165(.O (g21671), .I (I28201));
INVX1 gate9166(.O (I28206), .I (g20067));
INVX1 gate9167(.O (g21678), .I (I28206));
INVX1 gate9168(.O (I28210), .I (g20537));
INVX1 gate9169(.O (g21682), .I (I28210));
INVX1 gate9170(.O (g21690), .I (g19098));
INVX1 gate9171(.O (I28229), .I (g20067));
INVX1 gate9172(.O (g21700), .I (I28229));
INVX1 gate9173(.O (I28235), .I (g20153));
INVX1 gate9174(.O (g21708), .I (I28235));
INVX1 gate9175(.O (g21716), .I (g19894));
INVX1 gate9176(.O (g21726), .I (g19105));
INVX1 gate9177(.O (g21742), .I (g19919));
INVX1 gate9178(.O (g21752), .I (g19110));
INVX1 gate9179(.O (g21766), .I (g19934));
INVX1 gate9180(.O (g21782), .I (g19951));
INVX1 gate9181(.O (I28314), .I (g19152));
INVX1 gate9182(.O (g21795), .I (I28314));
INVX1 gate9183(.O (I28357), .I (g20497));
INVX1 gate9184(.O (g21824), .I (I28357));
INVX1 gate9185(.O (I28360), .I (g20163));
INVX1 gate9186(.O (g21825), .I (I28360));
INVX1 gate9187(.O (g21861), .I (g19657));
INVX1 gate9188(.O (g21867), .I (g19705));
INVX1 gate9189(.O (g21872), .I (g19749));
INVX1 gate9190(.O (g21876), .I (g19792));
INVX1 gate9191(.O (g21883), .I (g19890));
INVX1 gate9192(.O (g21886), .I (g19915));
INVX1 gate9193(.O (g21895), .I (g19945));
INVX1 gate9194(.O (g21902), .I (g19978));
INVX1 gate9195(.O (g21907), .I (g19972));
INVX1 gate9196(.O (I28432), .I (g19335));
INVX1 gate9197(.O (g21914), .I (I28432));
INVX1 gate9198(.O (I28435), .I (g19358));
INVX1 gate9199(.O (g21917), .I (I28435));
INVX1 gate9200(.O (g21921), .I (g20002));
INVX1 gate9201(.O (g21927), .I (g20045));
INVX1 gate9202(.O (I28443), .I (g19358));
INVX1 gate9203(.O (g21928), .I (I28443));
INVX1 gate9204(.O (I28447), .I (g19369));
INVX1 gate9205(.O (g21932), .I (I28447));
INVX1 gate9206(.O (I28450), .I (g19390));
INVX1 gate9207(.O (g21935), .I (I28450));
INVX1 gate9208(.O (g21939), .I (g20040));
INVX1 gate9209(.O (I28455), .I (g20943));
INVX1 gate9210(.O (g21943), .I (I28455));
INVX1 gate9211(.O (I28458), .I (g20971));
INVX1 gate9212(.O (g21944), .I (I28458));
INVX1 gate9213(.O (I28461), .I (g20998));
INVX1 gate9214(.O (g21945), .I (I28461));
INVX1 gate9215(.O (I28464), .I (g21024));
INVX1 gate9216(.O (g21946), .I (I28464));
INVX1 gate9217(.O (I28467), .I (g20942));
INVX1 gate9218(.O (g21947), .I (I28467));
INVX1 gate9219(.O (I28470), .I (g20984));
INVX1 gate9220(.O (g21948), .I (I28470));
INVX1 gate9221(.O (I28473), .I (g21030));
INVX1 gate9222(.O (g21949), .I (I28473));
INVX1 gate9223(.O (I28476), .I (g21064));
INVX1 gate9224(.O (g21950), .I (I28476));
INVX1 gate9225(.O (I28479), .I (g21795));
INVX1 gate9226(.O (g21951), .I (I28479));
INVX1 gate9227(.O (I28482), .I (g21376));
INVX1 gate9228(.O (g21952), .I (I28482));
INVX1 gate9229(.O (I28485), .I (g21426));
INVX1 gate9230(.O (g21953), .I (I28485));
INVX1 gate9231(.O (I28488), .I (g21495));
INVX1 gate9232(.O (g21954), .I (I28488));
INVX1 gate9233(.O (I28491), .I (g21327));
INVX1 gate9234(.O (g21955), .I (I28491));
INVX1 gate9235(.O (I28494), .I (g21358));
INVX1 gate9236(.O (g21956), .I (I28494));
INVX1 gate9237(.O (I28497), .I (g21399));
INVX1 gate9238(.O (g21957), .I (I28497));
INVX1 gate9239(.O (I28500), .I (g21457));
INVX1 gate9240(.O (g21958), .I (I28500));
INVX1 gate9241(.O (I28503), .I (g21528));
INVX1 gate9242(.O (g21959), .I (I28503));
INVX1 gate9243(.O (I28506), .I (g21377));
INVX1 gate9244(.O (g21960), .I (I28506));
INVX1 gate9245(.O (I28509), .I (g21427));
INVX1 gate9246(.O (g21961), .I (I28509));
INVX1 gate9247(.O (I28512), .I (g21496));
INVX1 gate9248(.O (g21962), .I (I28512));
INVX1 gate9249(.O (I28515), .I (g21557));
INVX1 gate9250(.O (g21963), .I (I28515));
INVX1 gate9251(.O (I28518), .I (g20985));
INVX1 gate9252(.O (g21964), .I (I28518));
INVX1 gate9253(.O (I28521), .I (g21824));
INVX1 gate9254(.O (g21965), .I (I28521));
INVX1 gate9255(.O (I28524), .I (g21359));
INVX1 gate9256(.O (g21966), .I (I28524));
INVX1 gate9257(.O (I28527), .I (g21407));
INVX1 gate9258(.O (g21967), .I (I28527));
INVX1 gate9259(.O (I28541), .I (g21467));
INVX1 gate9260(.O (g21982), .I (I28541));
INVX1 gate9261(.O (I28550), .I (g21432));
INVX1 gate9262(.O (g21995), .I (I28550));
INVX1 gate9263(.O (I28557), .I (g21407));
INVX1 gate9264(.O (g22003), .I (I28557));
INVX1 gate9265(.O (I28564), .I (g21385));
INVX1 gate9266(.O (g22014), .I (I28564));
INVX1 gate9267(.O (I28628), .I (g21842));
INVX1 gate9268(.O (g22082), .I (I28628));
INVX1 gate9269(.O (I28649), .I (g21843));
INVX1 gate9270(.O (g22107), .I (I28649));
INVX1 gate9271(.O (I28671), .I (g21845));
INVX1 gate9272(.O (g22133), .I (I28671));
INVX1 gate9273(.O (I28693), .I (g21847));
INVX1 gate9274(.O (g22156), .I (I28693));
INVX1 gate9275(.O (I28712), .I (g21851));
INVX1 gate9276(.O (g22176), .I (I28712));
INVX1 gate9277(.O (g22212), .I (g21914));
INVX1 gate9278(.O (g22213), .I (g21917));
INVX1 gate9279(.O (g22217), .I (g21928));
INVX1 gate9280(.O (I28781), .I (g21331));
INVX1 gate9281(.O (g22219), .I (I28781));
INVX1 gate9282(.O (g22221), .I (g21932));
INVX1 gate9283(.O (g22222), .I (g21935));
INVX1 gate9284(.O (I28789), .I (g21878));
INVX1 gate9285(.O (g22225), .I (I28789));
INVX1 gate9286(.O (I28792), .I (g21880));
INVX1 gate9287(.O (g22226), .I (I28792));
INVX1 gate9288(.O (g22230), .I (g20634));
INVX1 gate9289(.O (I28800), .I (g21316));
INVX1 gate9290(.O (g22232), .I (I28800));
INVX1 gate9291(.O (g22233), .I (g20637));
INVX1 gate9292(.O (g22236), .I (g20641));
INVX1 gate9293(.O (g22237), .I (g20644));
INVX1 gate9294(.O (g22239), .I (g20649));
INVX1 gate9295(.O (g22240), .I (g20652));
INVX1 gate9296(.O (g22241), .I (g20655));
INVX1 gate9297(.O (I28813), .I (g21502));
INVX1 gate9298(.O (g22243), .I (I28813));
INVX1 gate9299(.O (g22246), .I (g20659));
INVX1 gate9300(.O (g22248), .I (g20662));
INVX1 gate9301(.O (g22251), .I (g20666));
INVX1 gate9302(.O (g22252), .I (g20669));
INVX1 gate9303(.O (I28825), .I (g21882));
INVX1 gate9304(.O (g22253), .I (I28825));
INVX1 gate9305(.O (g22256), .I (g20673));
INVX1 gate9306(.O (g22257), .I (g20676));
INVX1 gate9307(.O (g22258), .I (g20679));
INVX1 gate9308(.O (I28833), .I (g21470));
INVX1 gate9309(.O (g22259), .I (I28833));
INVX1 gate9310(.O (g22260), .I (g20684));
INVX1 gate9311(.O (g22261), .I (g20687));
INVX1 gate9312(.O (g22262), .I (g20690));
INVX1 gate9313(.O (g22266), .I (g20694));
INVX1 gate9314(.O (g22268), .I (g20697));
INVX1 gate9315(.O (g22271), .I (g20704));
INVX1 gate9316(.O (g22274), .I (g20708));
INVX1 gate9317(.O (g22275), .I (g20711));
INVX1 gate9318(.O (g22276), .I (g20714));
INVX1 gate9319(.O (g22277), .I (g20719));
INVX1 gate9320(.O (g22278), .I (g20722));
INVX1 gate9321(.O (g22279), .I (g20725));
INVX1 gate9322(.O (g22283), .I (g20729));
INVX1 gate9323(.O (g22286), .I (g20732));
INVX1 gate9324(.O (g22287), .I (g20735));
INVX1 gate9325(.O (g22290), .I (g20739));
INVX1 gate9326(.O (g22293), .I (g20743));
INVX1 gate9327(.O (g22294), .I (g20746));
INVX1 gate9328(.O (g22295), .I (g20749));
INVX1 gate9329(.O (g22296), .I (g20754));
INVX1 gate9330(.O (g22297), .I (g20757));
INVX1 gate9331(.O (g22298), .I (g20760));
INVX1 gate9332(.O (I28876), .I (g21238));
INVX1 gate9333(.O (g22300), .I (I28876));
INVX1 gate9334(.O (g22303), .I (g20763));
INVX1 gate9335(.O (g22304), .I (g20766));
INVX1 gate9336(.O (g22306), .I (g20769));
INVX1 gate9337(.O (g22307), .I (g20772));
INVX1 gate9338(.O (g22310), .I (g20776));
INVX1 gate9339(.O (g22313), .I (g20780));
INVX1 gate9340(.O (g22314), .I (g20783));
INVX1 gate9341(.O (g22315), .I (g20786));
INVX1 gate9342(.O (g22316), .I (g21149));
INVX1 gate9343(.O (g22318), .I (g20790));
INVX1 gate9344(.O (g22319), .I (g21228));
INVX1 gate9345(.O (I28896), .I (g21246));
INVX1 gate9346(.O (g22328), .I (I28896));
INVX1 gate9347(.O (g22331), .I (g20793));
INVX1 gate9348(.O (g22332), .I (g20796));
INVX1 gate9349(.O (g22334), .I (g20799));
INVX1 gate9350(.O (g22335), .I (g20802));
INVX1 gate9351(.O (g22338), .I (g20806));
INVX1 gate9352(.O (g22341), .I (g21169));
INVX1 gate9353(.O (g22343), .I (g20810));
INVX1 gate9354(.O (g22344), .I (g21233));
INVX1 gate9355(.O (I28913), .I (g21255));
INVX1 gate9356(.O (g22353), .I (I28913));
INVX1 gate9357(.O (g22356), .I (g20813));
INVX1 gate9358(.O (g22357), .I (g20816));
INVX1 gate9359(.O (g22359), .I (g20819));
INVX1 gate9360(.O (g22360), .I (g20822));
INVX1 gate9361(.O (g22364), .I (g21189));
INVX1 gate9362(.O (g22366), .I (g20827));
INVX1 gate9363(.O (g22367), .I (g21242));
INVX1 gate9364(.O (I28928), .I (g21263));
INVX1 gate9365(.O (g22376), .I (I28928));
INVX1 gate9366(.O (g22379), .I (g20830));
INVX1 gate9367(.O (g22380), .I (g20833));
INVX1 gate9368(.O (g22384), .I (g21204));
INVX1 gate9369(.O (g22386), .I (g20837));
INVX1 gate9370(.O (g22387), .I (g21250));
INVX1 gate9371(.O (g22401), .I (g21533));
INVX1 gate9372(.O (g22402), .I (g21569));
INVX1 gate9373(.O (g22403), .I (g21602));
INVX1 gate9374(.O (g22404), .I (g21631));
INVX1 gate9375(.O (I28949), .I (g21685));
INVX1 gate9376(.O (g22405), .I (I28949));
INVX1 gate9377(.O (g22408), .I (g20986));
INVX1 gate9378(.O (I28953), .I (g21659));
INVX1 gate9379(.O (g22409), .I (I28953));
INVX1 gate9380(.O (I28956), .I (g21714));
INVX1 gate9381(.O (g22412), .I (I28956));
INVX1 gate9382(.O (I28959), .I (g21636));
INVX1 gate9383(.O (g22415), .I (I28959));
INVX1 gate9384(.O (I28962), .I (g21721));
INVX1 gate9385(.O (g22418), .I (I28962));
INVX1 gate9386(.O (g22421), .I (g21012));
INVX1 gate9387(.O (I28966), .I (g20633));
INVX1 gate9388(.O (g22422), .I (I28966));
INVX1 gate9389(.O (I28969), .I (g21686));
INVX1 gate9390(.O (g22425), .I (I28969));
INVX1 gate9391(.O (I28972), .I (g21736));
INVX1 gate9392(.O (g22428), .I (I28972));
INVX1 gate9393(.O (I28975), .I (g21688));
INVX1 gate9394(.O (g22431), .I (I28975));
INVX1 gate9395(.O (I28978), .I (g21740));
INVX1 gate9396(.O (g22434), .I (I28978));
INVX1 gate9397(.O (I28981), .I (g21667));
INVX1 gate9398(.O (g22437), .I (I28981));
INVX1 gate9399(.O (I28984), .I (g21747));
INVX1 gate9400(.O (g22440), .I (I28984));
INVX1 gate9401(.O (g22443), .I (g21036));
INVX1 gate9402(.O (I28988), .I (g20874));
INVX1 gate9403(.O (g22444), .I (I28988));
INVX1 gate9404(.O (I28991), .I (g20648));
INVX1 gate9405(.O (g22445), .I (I28991));
INVX1 gate9406(.O (I28994), .I (g21715));
INVX1 gate9407(.O (g22448), .I (I28994));
INVX1 gate9408(.O (I28997), .I (g21759));
INVX1 gate9409(.O (g22451), .I (I28997));
INVX1 gate9410(.O (I29001), .I (g20658));
INVX1 gate9411(.O (g22455), .I (I29001));
INVX1 gate9412(.O (I29004), .I (g21722));
INVX1 gate9413(.O (g22458), .I (I29004));
INVX1 gate9414(.O (I29007), .I (g21760));
INVX1 gate9415(.O (g22461), .I (I29007));
INVX1 gate9416(.O (I29010), .I (g21724));
INVX1 gate9417(.O (g22464), .I (I29010));
INVX1 gate9418(.O (I29013), .I (g21764));
INVX1 gate9419(.O (g22467), .I (I29013));
INVX1 gate9420(.O (I29016), .I (g21696));
INVX1 gate9421(.O (g22470), .I (I29016));
INVX1 gate9422(.O (I29019), .I (g21771));
INVX1 gate9423(.O (g22473), .I (I29019));
INVX1 gate9424(.O (g22476), .I (g21057));
INVX1 gate9425(.O (I29023), .I (g20672));
INVX1 gate9426(.O (g22477), .I (I29023));
INVX1 gate9427(.O (I29026), .I (g21737));
INVX1 gate9428(.O (g22480), .I (I29026));
INVX1 gate9429(.O (I29030), .I (g20683));
INVX1 gate9430(.O (g22484), .I (I29030));
INVX1 gate9431(.O (I29033), .I (g21741));
INVX1 gate9432(.O (g22487), .I (I29033));
INVX1 gate9433(.O (I29036), .I (g21775));
INVX1 gate9434(.O (g22490), .I (I29036));
INVX1 gate9435(.O (I29040), .I (g20693));
INVX1 gate9436(.O (g22494), .I (I29040));
INVX1 gate9437(.O (I29043), .I (g21748));
INVX1 gate9438(.O (g22497), .I (I29043));
INVX1 gate9439(.O (I29046), .I (g21776));
INVX1 gate9440(.O (g22500), .I (I29046));
INVX1 gate9441(.O (I29049), .I (g21750));
INVX1 gate9442(.O (g22503), .I (I29049));
INVX1 gate9443(.O (I29052), .I (g21780));
INVX1 gate9444(.O (g22506), .I (I29052));
INVX1 gate9445(.O (I29055), .I (g21732));
INVX1 gate9446(.O (g22509), .I (I29055));
INVX1 gate9447(.O (I29058), .I (g20703));
INVX1 gate9448(.O (g22512), .I (I29058));
INVX1 gate9449(.O (I29064), .I (g20875));
INVX1 gate9450(.O (g22518), .I (I29064));
INVX1 gate9451(.O (I29067), .I (g20876));
INVX1 gate9452(.O (g22519), .I (I29067));
INVX1 gate9453(.O (I29070), .I (g20707));
INVX1 gate9454(.O (g22520), .I (I29070));
INVX1 gate9455(.O (I29073), .I (g21761));
INVX1 gate9456(.O (g22523), .I (I29073));
INVX1 gate9457(.O (I29077), .I (g20718));
INVX1 gate9458(.O (g22527), .I (I29077));
INVX1 gate9459(.O (I29080), .I (g21765));
INVX1 gate9460(.O (g22530), .I (I29080));
INVX1 gate9461(.O (I29083), .I (g21790));
INVX1 gate9462(.O (g22533), .I (I29083));
INVX1 gate9463(.O (I29087), .I (g20728));
INVX1 gate9464(.O (g22537), .I (I29087));
INVX1 gate9465(.O (I29090), .I (g21772));
INVX1 gate9466(.O (g22540), .I (I29090));
INVX1 gate9467(.O (I29093), .I (g21791));
INVX1 gate9468(.O (g22543), .I (I29093));
INVX1 gate9469(.O (g22547), .I (g21087));
INVX1 gate9470(.O (I29098), .I (g20879));
INVX1 gate9471(.O (g22548), .I (I29098));
INVX1 gate9472(.O (I29101), .I (g20880));
INVX1 gate9473(.O (g22549), .I (I29101));
INVX1 gate9474(.O (I29104), .I (g20881));
INVX1 gate9475(.O (g22550), .I (I29104));
INVX1 gate9476(.O (I29107), .I (g21435));
INVX1 gate9477(.O (g22551), .I (I29107));
INVX1 gate9478(.O (I29110), .I (g20738));
INVX1 gate9479(.O (g22552), .I (I29110));
INVX1 gate9480(.O (I29116), .I (g20882));
INVX1 gate9481(.O (g22558), .I (I29116));
INVX1 gate9482(.O (I29119), .I (g20883));
INVX1 gate9483(.O (g22559), .I (I29119));
INVX1 gate9484(.O (I29122), .I (g20742));
INVX1 gate9485(.O (g22560), .I (I29122));
INVX1 gate9486(.O (I29125), .I (g21777));
INVX1 gate9487(.O (g22563), .I (I29125));
INVX1 gate9488(.O (I29129), .I (g20753));
INVX1 gate9489(.O (g22567), .I (I29129));
INVX1 gate9490(.O (I29132), .I (g21781));
INVX1 gate9491(.O (g22570), .I (I29132));
INVX1 gate9492(.O (I29135), .I (g21804));
INVX1 gate9493(.O (g22573), .I (I29135));
INVX1 gate9494(.O (I29142), .I (g20682));
INVX1 gate9495(.O (g22582), .I (I29142));
INVX1 gate9496(.O (I29145), .I (g20891));
INVX1 gate9497(.O (g22583), .I (I29145));
INVX1 gate9498(.O (I29148), .I (g20892));
INVX1 gate9499(.O (g22584), .I (I29148));
INVX1 gate9500(.O (I29151), .I (g20893));
INVX1 gate9501(.O (g22585), .I (I29151));
INVX1 gate9502(.O (I29154), .I (g20894));
INVX1 gate9503(.O (g22586), .I (I29154));
INVX1 gate9504(.O (g22588), .I (g21099));
INVX1 gate9505(.O (I29159), .I (g20896));
INVX1 gate9506(.O (g22589), .I (I29159));
INVX1 gate9507(.O (I29162), .I (g20897));
INVX1 gate9508(.O (g22590), .I (I29162));
INVX1 gate9509(.O (I29165), .I (g20898));
INVX1 gate9510(.O (g22591), .I (I29165));
INVX1 gate9511(.O (I29168), .I (g20775));
INVX1 gate9512(.O (g22592), .I (I29168));
INVX1 gate9513(.O (I29174), .I (g20899));
INVX1 gate9514(.O (g22598), .I (I29174));
INVX1 gate9515(.O (I29177), .I (g20900));
INVX1 gate9516(.O (g22599), .I (I29177));
INVX1 gate9517(.O (I29180), .I (g20779));
INVX1 gate9518(.O (g22600), .I (I29180));
INVX1 gate9519(.O (I29183), .I (g21792));
INVX1 gate9520(.O (g22603), .I (I29183));
INVX1 gate9521(.O (g22609), .I (g21108));
INVX1 gate9522(.O (I29191), .I (g20901));
INVX1 gate9523(.O (g22611), .I (I29191));
INVX1 gate9524(.O (I29194), .I (g20902));
INVX1 gate9525(.O (g22612), .I (I29194));
INVX1 gate9526(.O (I29197), .I (g20903));
INVX1 gate9527(.O (g22613), .I (I29197));
INVX1 gate9528(.O (I29203), .I (g20717));
INVX1 gate9529(.O (g22619), .I (I29203));
INVX1 gate9530(.O (I29206), .I (g20910));
INVX1 gate9531(.O (g22620), .I (I29206));
INVX1 gate9532(.O (I29209), .I (g20911));
INVX1 gate9533(.O (g22621), .I (I29209));
INVX1 gate9534(.O (I29212), .I (g20912));
INVX1 gate9535(.O (g22622), .I (I29212));
INVX1 gate9536(.O (I29215), .I (g20913));
INVX1 gate9537(.O (g22623), .I (I29215));
INVX1 gate9538(.O (g22625), .I (g21113));
INVX1 gate9539(.O (I29220), .I (g20915));
INVX1 gate9540(.O (g22626), .I (I29220));
INVX1 gate9541(.O (I29223), .I (g20916));
INVX1 gate9542(.O (g22627), .I (I29223));
INVX1 gate9543(.O (I29226), .I (g20917));
INVX1 gate9544(.O (g22628), .I (I29226));
INVX1 gate9545(.O (I29229), .I (g20805));
INVX1 gate9546(.O (g22629), .I (I29229));
INVX1 gate9547(.O (I29235), .I (g20918));
INVX1 gate9548(.O (g22635), .I (I29235));
INVX1 gate9549(.O (I29238), .I (g20919));
INVX1 gate9550(.O (g22636), .I (I29238));
INVX1 gate9551(.O (I29243), .I (g20921));
INVX1 gate9552(.O (g22639), .I (I29243));
INVX1 gate9553(.O (I29246), .I (g20922));
INVX1 gate9554(.O (g22640), .I (I29246));
INVX1 gate9555(.O (I29249), .I (g20923));
INVX1 gate9556(.O (g22641), .I (I29249));
INVX1 gate9557(.O (I29252), .I (g20924));
INVX1 gate9558(.O (g22642), .I (I29252));
INVX1 gate9559(.O (g22645), .I (g21125));
INVX1 gate9560(.O (I29259), .I (g20925));
INVX1 gate9561(.O (g22647), .I (I29259));
INVX1 gate9562(.O (I29262), .I (g20926));
INVX1 gate9563(.O (g22648), .I (I29262));
INVX1 gate9564(.O (I29265), .I (g20927));
INVX1 gate9565(.O (g22649), .I (I29265));
INVX1 gate9566(.O (I29271), .I (g20752));
INVX1 gate9567(.O (g22655), .I (I29271));
INVX1 gate9568(.O (I29274), .I (g20934));
INVX1 gate9569(.O (g22656), .I (I29274));
INVX1 gate9570(.O (I29277), .I (g20935));
INVX1 gate9571(.O (g22657), .I (I29277));
INVX1 gate9572(.O (I29280), .I (g20936));
INVX1 gate9573(.O (g22658), .I (I29280));
INVX1 gate9574(.O (I29283), .I (g20937));
INVX1 gate9575(.O (g22659), .I (I29283));
INVX1 gate9576(.O (g22661), .I (g21130));
INVX1 gate9577(.O (I29288), .I (g20939));
INVX1 gate9578(.O (g22662), .I (I29288));
INVX1 gate9579(.O (I29291), .I (g20940));
INVX1 gate9580(.O (g22663), .I (I29291));
INVX1 gate9581(.O (I29294), .I (g20941));
INVX1 gate9582(.O (g22664), .I (I29294));
INVX1 gate9583(.O (I29301), .I (g20944));
INVX1 gate9584(.O (g22669), .I (I29301));
INVX1 gate9585(.O (I29304), .I (g20945));
INVX1 gate9586(.O (g22670), .I (I29304));
INVX1 gate9587(.O (I29307), .I (g20946));
INVX1 gate9588(.O (g22671), .I (I29307));
INVX1 gate9589(.O (I29310), .I (g20947));
INVX1 gate9590(.O (g22672), .I (I29310));
INVX1 gate9591(.O (I29313), .I (g20948));
INVX1 gate9592(.O (g22673), .I (I29313));
INVX1 gate9593(.O (I29317), .I (g20949));
INVX1 gate9594(.O (g22675), .I (I29317));
INVX1 gate9595(.O (I29320), .I (g20950));
INVX1 gate9596(.O (g22676), .I (I29320));
INVX1 gate9597(.O (I29323), .I (g20951));
INVX1 gate9598(.O (g22677), .I (I29323));
INVX1 gate9599(.O (I29326), .I (g20952));
INVX1 gate9600(.O (g22678), .I (I29326));
INVX1 gate9601(.O (g22681), .I (g21144));
INVX1 gate9602(.O (I29333), .I (g20953));
INVX1 gate9603(.O (g22683), .I (I29333));
INVX1 gate9604(.O (I29336), .I (g20954));
INVX1 gate9605(.O (g22684), .I (I29336));
INVX1 gate9606(.O (I29339), .I (g20955));
INVX1 gate9607(.O (g22685), .I (I29339));
INVX1 gate9608(.O (I29345), .I (g20789));
INVX1 gate9609(.O (g22691), .I (I29345));
INVX1 gate9610(.O (I29348), .I (g20962));
INVX1 gate9611(.O (g22692), .I (I29348));
INVX1 gate9612(.O (I29351), .I (g20963));
INVX1 gate9613(.O (g22693), .I (I29351));
INVX1 gate9614(.O (I29354), .I (g20964));
INVX1 gate9615(.O (g22694), .I (I29354));
INVX1 gate9616(.O (I29357), .I (g20965));
INVX1 gate9617(.O (g22695), .I (I29357));
INVX1 gate9618(.O (I29360), .I (g21796));
INVX1 gate9619(.O (g22696), .I (I29360));
INVX1 gate9620(.O (I29366), .I (g20966));
INVX1 gate9621(.O (g22702), .I (I29366));
INVX1 gate9622(.O (I29369), .I (g20967));
INVX1 gate9623(.O (g22703), .I (I29369));
INVX1 gate9624(.O (I29372), .I (g20968));
INVX1 gate9625(.O (g22704), .I (I29372));
INVX1 gate9626(.O (I29375), .I (g20969));
INVX1 gate9627(.O (g22705), .I (I29375));
INVX1 gate9628(.O (I29378), .I (g20970));
INVX1 gate9629(.O (g22706), .I (I29378));
INVX1 gate9630(.O (I29383), .I (g20972));
INVX1 gate9631(.O (g22709), .I (I29383));
INVX1 gate9632(.O (I29386), .I (g20973));
INVX1 gate9633(.O (g22710), .I (I29386));
INVX1 gate9634(.O (I29389), .I (g20974));
INVX1 gate9635(.O (g22711), .I (I29389));
INVX1 gate9636(.O (I29392), .I (g20975));
INVX1 gate9637(.O (g22712), .I (I29392));
INVX1 gate9638(.O (I29395), .I (g20976));
INVX1 gate9639(.O (g22713), .I (I29395));
INVX1 gate9640(.O (I29399), .I (g20977));
INVX1 gate9641(.O (g22715), .I (I29399));
INVX1 gate9642(.O (I29402), .I (g20978));
INVX1 gate9643(.O (g22716), .I (I29402));
INVX1 gate9644(.O (I29405), .I (g20979));
INVX1 gate9645(.O (g22717), .I (I29405));
INVX1 gate9646(.O (I29408), .I (g20980));
INVX1 gate9647(.O (g22718), .I (I29408));
INVX1 gate9648(.O (g22721), .I (g21164));
INVX1 gate9649(.O (I29415), .I (g20981));
INVX1 gate9650(.O (g22723), .I (I29415));
INVX1 gate9651(.O (I29418), .I (g20982));
INVX1 gate9652(.O (g22724), .I (I29418));
INVX1 gate9653(.O (I29421), .I (g20983));
INVX1 gate9654(.O (g22725), .I (I29421));
INVX1 gate9655(.O (I29426), .I (g20989));
INVX1 gate9656(.O (g22728), .I (I29426));
INVX1 gate9657(.O (I29429), .I (g20990));
INVX1 gate9658(.O (g22729), .I (I29429));
INVX1 gate9659(.O (I29432), .I (g20991));
INVX1 gate9660(.O (g22730), .I (I29432));
INVX1 gate9661(.O (I29435), .I (g20992));
INVX1 gate9662(.O (g22731), .I (I29435));
INVX1 gate9663(.O (I29439), .I (g20993));
INVX1 gate9664(.O (g22733), .I (I29439));
INVX1 gate9665(.O (I29442), .I (g20994));
INVX1 gate9666(.O (g22734), .I (I29442));
INVX1 gate9667(.O (I29445), .I (g20995));
INVX1 gate9668(.O (g22735), .I (I29445));
INVX1 gate9669(.O (I29448), .I (g20996));
INVX1 gate9670(.O (g22736), .I (I29448));
INVX1 gate9671(.O (I29451), .I (g20997));
INVX1 gate9672(.O (g22737), .I (I29451));
INVX1 gate9673(.O (I29456), .I (g20999));
INVX1 gate9674(.O (g22740), .I (I29456));
INVX1 gate9675(.O (I29459), .I (g21000));
INVX1 gate9676(.O (g22741), .I (I29459));
INVX1 gate9677(.O (I29462), .I (g21001));
INVX1 gate9678(.O (g22742), .I (I29462));
INVX1 gate9679(.O (I29465), .I (g21002));
INVX1 gate9680(.O (g22743), .I (I29465));
INVX1 gate9681(.O (I29468), .I (g21003));
INVX1 gate9682(.O (g22744), .I (I29468));
INVX1 gate9683(.O (I29472), .I (g21004));
INVX1 gate9684(.O (g22746), .I (I29472));
INVX1 gate9685(.O (I29475), .I (g21005));
INVX1 gate9686(.O (g22747), .I (I29475));
INVX1 gate9687(.O (I29478), .I (g21006));
INVX1 gate9688(.O (g22748), .I (I29478));
INVX1 gate9689(.O (I29481), .I (g21007));
INVX1 gate9690(.O (g22749), .I (I29481));
INVX1 gate9691(.O (I29484), .I (g21903));
INVX1 gate9692(.O (g22750), .I (I29484));
INVX1 gate9693(.O (g22753), .I (g21184));
INVX1 gate9694(.O (I29490), .I (g21009));
INVX1 gate9695(.O (g22756), .I (I29490));
INVX1 gate9696(.O (I29493), .I (g21010));
INVX1 gate9697(.O (g22757), .I (I29493));
INVX1 gate9698(.O (I29496), .I (g21011));
INVX1 gate9699(.O (g22758), .I (I29496));
INVX1 gate9700(.O (I29500), .I (g21015));
INVX1 gate9701(.O (g22760), .I (I29500));
INVX1 gate9702(.O (I29503), .I (g21016));
INVX1 gate9703(.O (g22761), .I (I29503));
INVX1 gate9704(.O (I29506), .I (g21017));
INVX1 gate9705(.O (g22762), .I (I29506));
INVX1 gate9706(.O (I29509), .I (g21018));
INVX1 gate9707(.O (g22763), .I (I29509));
INVX1 gate9708(.O (I29513), .I (g21019));
INVX1 gate9709(.O (g22765), .I (I29513));
INVX1 gate9710(.O (I29516), .I (g21020));
INVX1 gate9711(.O (g22766), .I (I29516));
INVX1 gate9712(.O (I29519), .I (g21021));
INVX1 gate9713(.O (g22767), .I (I29519));
INVX1 gate9714(.O (I29522), .I (g21022));
INVX1 gate9715(.O (g22768), .I (I29522));
INVX1 gate9716(.O (I29525), .I (g21023));
INVX1 gate9717(.O (g22769), .I (I29525));
INVX1 gate9718(.O (I29530), .I (g21025));
INVX1 gate9719(.O (g22772), .I (I29530));
INVX1 gate9720(.O (I29533), .I (g21026));
INVX1 gate9721(.O (g22773), .I (I29533));
INVX1 gate9722(.O (I29536), .I (g21027));
INVX1 gate9723(.O (g22774), .I (I29536));
INVX1 gate9724(.O (I29539), .I (g21028));
INVX1 gate9725(.O (g22775), .I (I29539));
INVX1 gate9726(.O (I29542), .I (g21029));
INVX1 gate9727(.O (g22776), .I (I29542));
INVX1 gate9728(.O (g22777), .I (g21796));
INVX1 gate9729(.O (I29547), .I (g21031));
INVX1 gate9730(.O (g22785), .I (I29547));
INVX1 gate9731(.O (I29550), .I (g21032));
INVX1 gate9732(.O (g22786), .I (I29550));
INVX1 gate9733(.O (g22787), .I (g21199));
INVX1 gate9734(.O (I29556), .I (g21033));
INVX1 gate9735(.O (g22790), .I (I29556));
INVX1 gate9736(.O (I29559), .I (g21034));
INVX1 gate9737(.O (g22791), .I (I29559));
INVX1 gate9738(.O (I29562), .I (g21035));
INVX1 gate9739(.O (g22792), .I (I29562));
INVX1 gate9740(.O (I29566), .I (g21039));
INVX1 gate9741(.O (g22794), .I (I29566));
INVX1 gate9742(.O (I29569), .I (g21040));
INVX1 gate9743(.O (g22795), .I (I29569));
INVX1 gate9744(.O (I29572), .I (g21041));
INVX1 gate9745(.O (g22796), .I (I29572));
INVX1 gate9746(.O (I29575), .I (g21042));
INVX1 gate9747(.O (g22797), .I (I29575));
INVX1 gate9748(.O (I29579), .I (g21043));
INVX1 gate9749(.O (g22799), .I (I29579));
INVX1 gate9750(.O (I29582), .I (g21044));
INVX1 gate9751(.O (g22800), .I (I29582));
INVX1 gate9752(.O (I29585), .I (g21045));
INVX1 gate9753(.O (g22801), .I (I29585));
INVX1 gate9754(.O (I29588), .I (g21046));
INVX1 gate9755(.O (g22802), .I (I29588));
INVX1 gate9756(.O (I29591), .I (g21047));
INVX1 gate9757(.O (g22803), .I (I29591));
INVX1 gate9758(.O (g22805), .I (g21894));
INVX1 gate9759(.O (g22806), .I (g21615));
INVX1 gate9760(.O (I29600), .I (g21720));
INVX1 gate9761(.O (g22812), .I (I29600));
INVX1 gate9762(.O (I29603), .I (g21051));
INVX1 gate9763(.O (g22824), .I (I29603));
INVX1 gate9764(.O (I29606), .I (g21364));
INVX1 gate9765(.O (g22825), .I (I29606));
INVX1 gate9766(.O (I29610), .I (g21052));
INVX1 gate9767(.O (g22827), .I (I29610));
INVX1 gate9768(.O (I29613), .I (g21053));
INVX1 gate9769(.O (g22828), .I (I29613));
INVX1 gate9770(.O (g22829), .I (g21214));
INVX1 gate9771(.O (I29619), .I (g21054));
INVX1 gate9772(.O (g22832), .I (I29619));
INVX1 gate9773(.O (I29622), .I (g21055));
INVX1 gate9774(.O (g22833), .I (I29622));
INVX1 gate9775(.O (I29625), .I (g21056));
INVX1 gate9776(.O (g22834), .I (I29625));
INVX1 gate9777(.O (I29629), .I (g21060));
INVX1 gate9778(.O (g22836), .I (I29629));
INVX1 gate9779(.O (I29632), .I (g21061));
INVX1 gate9780(.O (g22837), .I (I29632));
INVX1 gate9781(.O (I29635), .I (g21062));
INVX1 gate9782(.O (g22838), .I (I29635));
INVX1 gate9783(.O (I29638), .I (g21063));
INVX1 gate9784(.O (g22839), .I (I29638));
INVX1 gate9785(.O (I29641), .I (g20825));
INVX1 gate9786(.O (g22840), .I (I29641));
INVX1 gate9787(.O (g22843), .I (g21889));
INVX1 gate9788(.O (g22847), .I (g21643));
INVX1 gate9789(.O (I29653), .I (g21746));
INVX1 gate9790(.O (g22852), .I (I29653));
INVX1 gate9791(.O (I29656), .I (g21070));
INVX1 gate9792(.O (g22864), .I (I29656));
INVX1 gate9793(.O (I29660), .I (g21071));
INVX1 gate9794(.O (g22866), .I (I29660));
INVX1 gate9795(.O (I29663), .I (g21072));
INVX1 gate9796(.O (g22867), .I (I29663));
INVX1 gate9797(.O (g22868), .I (g21222));
INVX1 gate9798(.O (I29669), .I (g21073));
INVX1 gate9799(.O (g22871), .I (I29669));
INVX1 gate9800(.O (I29672), .I (g21074));
INVX1 gate9801(.O (g22872), .I (I29672));
INVX1 gate9802(.O (I29675), .I (g21075));
INVX1 gate9803(.O (g22873), .I (I29675));
INVX1 gate9804(.O (g22875), .I (g21884));
INVX1 gate9805(.O (g22882), .I (g21674));
INVX1 gate9806(.O (I29687), .I (g21770));
INVX1 gate9807(.O (g22887), .I (I29687));
INVX1 gate9808(.O (I29690), .I (g21080));
INVX1 gate9809(.O (g22899), .I (I29690));
INVX1 gate9810(.O (I29694), .I (g21081));
INVX1 gate9811(.O (g22901), .I (I29694));
INVX1 gate9812(.O (I29697), .I (g21082));
INVX1 gate9813(.O (g22902), .I (I29697));
INVX1 gate9814(.O (I29700), .I (g20700));
INVX1 gate9815(.O (g22903), .I (I29700));
INVX1 gate9816(.O (g22907), .I (g21711));
INVX1 gate9817(.O (g22917), .I (g21703));
INVX1 gate9818(.O (I29712), .I (g21786));
INVX1 gate9819(.O (g22922), .I (I29712));
INVX1 gate9820(.O (I29715), .I (g21094));
INVX1 gate9821(.O (g22934), .I (I29715));
INVX1 gate9822(.O (I29724), .I (g21851));
INVX1 gate9823(.O (g22945), .I (I29724));
INVX1 gate9824(.O (I29727), .I (g20877));
INVX1 gate9825(.O (g22948), .I (I29727));
INVX1 gate9826(.O (g22949), .I (g21665));
INVX1 gate9827(.O (g22954), .I (g21739));
INVX1 gate9828(.O (g22958), .I (g21694));
INVX1 gate9829(.O (g22962), .I (g21763));
INVX1 gate9830(.O (g22966), .I (g21730));
INVX1 gate9831(.O (I29736), .I (g20884));
INVX1 gate9832(.O (g22970), .I (I29736));
INVX1 gate9833(.O (g22971), .I (g21779));
INVX1 gate9834(.O (g22975), .I (g21756));
INVX1 gate9835(.O (I29741), .I (g21346));
INVX1 gate9836(.O (g22979), .I (I29741));
INVX1 gate9837(.O (g22980), .I (g21794));
INVX1 gate9838(.O (g22986), .I (g21382));
INVX1 gate9839(.O (g22988), .I (g21404));
INVX1 gate9840(.O (g22989), .I (g21415));
INVX1 gate9841(.O (g22991), .I (g21429));
INVX1 gate9842(.O (g22995), .I (g21441));
INVX1 gate9843(.O (g22996), .I (g21449));
INVX1 gate9844(.O (g22998), .I (g21458));
INVX1 gate9845(.O (g23001), .I (g21473));
INVX1 gate9846(.O (g23002), .I (g21477));
INVX1 gate9847(.O (g23006), .I (g21483));
INVX1 gate9848(.O (g23007), .I (g21491));
INVX1 gate9849(.O (g23008), .I (g21498));
INVX1 gate9850(.O (g23012), .I (g21505));
INVX1 gate9851(.O (g23015), .I (g21514));
INVX1 gate9852(.O (g23016), .I (g21518));
INVX1 gate9853(.O (g23020), .I (g21524));
INVX1 gate9854(.O (g23021), .I (g21530));
INVX1 gate9855(.O (g23024), .I (g21537));
INVX1 gate9856(.O (g23028), .I (g21541));
INVX1 gate9857(.O (g23031), .I (g21550));
INVX1 gate9858(.O (g23032), .I (g21554));
INVX1 gate9859(.O (g23036), .I (g21558));
INVX1 gate9860(.O (g23037), .I (g21561));
INVX1 gate9861(.O (g23038), .I (g21566));
INVX1 gate9862(.O (g23041), .I (g21573));
INVX1 gate9863(.O (g23045), .I (g21577));
INVX1 gate9864(.O (g23048), .I (g21586));
INVX1 gate9865(.O (g23049), .I (g21590));
INVX1 gate9866(.O (I29797), .I (g21432));
INVX1 gate9867(.O (g23050), .I (I29797));
INVX1 gate9868(.O (I29802), .I (g21435));
INVX1 gate9869(.O (g23055), .I (I29802));
INVX1 gate9870(.O (g23056), .I (g21594));
INVX1 gate9871(.O (g23057), .I (g21599));
INVX1 gate9872(.O (g23060), .I (g21606));
INVX1 gate9873(.O (g23064), .I (g21612));
INVX1 gate9874(.O (I29812), .I (g21467));
INVX1 gate9875(.O (g23065), .I (I29812));
INVX1 gate9876(.O (I29817), .I (g21470));
INVX1 gate9877(.O (g23068), .I (I29817));
INVX1 gate9878(.O (g23069), .I (g21619));
INVX1 gate9879(.O (g23074), .I (g21623));
INVX1 gate9880(.O (g23075), .I (g21628));
INVX1 gate9881(.O (I29827), .I (g21502));
INVX1 gate9882(.O (g23078), .I (I29827));
INVX1 gate9883(.O (g23079), .I (g21640));
INVX1 gate9884(.O (g23082), .I (g21647));
INVX1 gate9885(.O (g23087), .I (g21651));
INVX1 gate9886(.O (g23088), .I (g21655));
INVX1 gate9887(.O (I29841), .I (g21316));
INVX1 gate9888(.O (g23094), .I (I29841));
INVX1 gate9889(.O (g23095), .I (g21671));
INVX1 gate9890(.O (g23098), .I (g21678));
INVX1 gate9891(.O (g23103), .I (g21682));
INVX1 gate9892(.O (I29852), .I (g21331));
INVX1 gate9893(.O (g23105), .I (I29852));
INVX1 gate9894(.O (g23112), .I (g21700));
INVX1 gate9895(.O (g23115), .I (g21708));
INVX1 gate9896(.O (I29863), .I (g21346));
INVX1 gate9897(.O (g23116), .I (I29863));
INVX1 gate9898(.O (I29872), .I (g21364));
INVX1 gate9899(.O (g23125), .I (I29872));
INVX1 gate9900(.O (I29881), .I (g21385));
INVX1 gate9901(.O (g23134), .I (I29881));
INVX1 gate9902(.O (g23140), .I (g21825));
INVX1 gate9903(.O (g23141), .I (g21825));
INVX1 gate9904(.O (g23142), .I (g21825));
INVX1 gate9905(.O (g23143), .I (g21825));
INVX1 gate9906(.O (g23144), .I (g21825));
INVX1 gate9907(.O (g23145), .I (g21825));
INVX1 gate9908(.O (g23146), .I (g21825));
INVX1 gate9909(.O (g23147), .I (g21825));
INVX1 gate9910(.O (I29897), .I (g23116));
INVX1 gate9911(.O (g23148), .I (I29897));
INVX1 gate9912(.O (I29900), .I (g23125));
INVX1 gate9913(.O (g23149), .I (I29900));
INVX1 gate9914(.O (I29903), .I (g23134));
INVX1 gate9915(.O (g23150), .I (I29903));
INVX1 gate9916(.O (I29906), .I (g21967));
INVX1 gate9917(.O (g23151), .I (I29906));
INVX1 gate9918(.O (I29909), .I (g23050));
INVX1 gate9919(.O (g23152), .I (I29909));
INVX1 gate9920(.O (I29912), .I (g23065));
INVX1 gate9921(.O (g23153), .I (I29912));
INVX1 gate9922(.O (I29915), .I (g23055));
INVX1 gate9923(.O (g23154), .I (I29915));
INVX1 gate9924(.O (I29918), .I (g23068));
INVX1 gate9925(.O (g23155), .I (I29918));
INVX1 gate9926(.O (I29921), .I (g23078));
INVX1 gate9927(.O (g23156), .I (I29921));
INVX1 gate9928(.O (I29924), .I (g23094));
INVX1 gate9929(.O (g23157), .I (I29924));
INVX1 gate9930(.O (I29927), .I (g23105));
INVX1 gate9931(.O (g23158), .I (I29927));
INVX1 gate9932(.O (I29930), .I (g22176));
INVX1 gate9933(.O (g23159), .I (I29930));
INVX1 gate9934(.O (I29933), .I (g22082));
INVX1 gate9935(.O (g23160), .I (I29933));
INVX1 gate9936(.O (I29936), .I (g22582));
INVX1 gate9937(.O (g23161), .I (I29936));
INVX1 gate9938(.O (I29939), .I (g22518));
INVX1 gate9939(.O (g23162), .I (I29939));
INVX1 gate9940(.O (I29942), .I (g22548));
INVX1 gate9941(.O (g23163), .I (I29942));
INVX1 gate9942(.O (I29945), .I (g22583));
INVX1 gate9943(.O (g23164), .I (I29945));
INVX1 gate9944(.O (I29948), .I (g22549));
INVX1 gate9945(.O (g23165), .I (I29948));
INVX1 gate9946(.O (I29951), .I (g22584));
INVX1 gate9947(.O (g23166), .I (I29951));
INVX1 gate9948(.O (I29954), .I (g22611));
INVX1 gate9949(.O (g23167), .I (I29954));
INVX1 gate9950(.O (I29957), .I (g22585));
INVX1 gate9951(.O (g23168), .I (I29957));
INVX1 gate9952(.O (I29960), .I (g22612));
INVX1 gate9953(.O (g23169), .I (I29960));
INVX1 gate9954(.O (I29963), .I (g22639));
INVX1 gate9955(.O (g23170), .I (I29963));
INVX1 gate9956(.O (I29966), .I (g22613));
INVX1 gate9957(.O (g23171), .I (I29966));
INVX1 gate9958(.O (I29969), .I (g22640));
INVX1 gate9959(.O (g23172), .I (I29969));
INVX1 gate9960(.O (I29972), .I (g22669));
INVX1 gate9961(.O (g23173), .I (I29972));
INVX1 gate9962(.O (I29975), .I (g22641));
INVX1 gate9963(.O (g23174), .I (I29975));
INVX1 gate9964(.O (I29978), .I (g22670));
INVX1 gate9965(.O (g23175), .I (I29978));
INVX1 gate9966(.O (I29981), .I (g22702));
INVX1 gate9967(.O (g23176), .I (I29981));
INVX1 gate9968(.O (I29984), .I (g22671));
INVX1 gate9969(.O (g23177), .I (I29984));
INVX1 gate9970(.O (I29987), .I (g22703));
INVX1 gate9971(.O (g23178), .I (I29987));
INVX1 gate9972(.O (I29990), .I (g22728));
INVX1 gate9973(.O (g23179), .I (I29990));
INVX1 gate9974(.O (I29993), .I (g22704));
INVX1 gate9975(.O (g23180), .I (I29993));
INVX1 gate9976(.O (I29996), .I (g22729));
INVX1 gate9977(.O (g23181), .I (I29996));
INVX1 gate9978(.O (I29999), .I (g22756));
INVX1 gate9979(.O (g23182), .I (I29999));
INVX1 gate9980(.O (I30002), .I (g22730));
INVX1 gate9981(.O (g23183), .I (I30002));
INVX1 gate9982(.O (I30005), .I (g22757));
INVX1 gate9983(.O (g23184), .I (I30005));
INVX1 gate9984(.O (I30008), .I (g22785));
INVX1 gate9985(.O (g23185), .I (I30008));
INVX1 gate9986(.O (I30011), .I (g22758));
INVX1 gate9987(.O (g23186), .I (I30011));
INVX1 gate9988(.O (I30014), .I (g22786));
INVX1 gate9989(.O (g23187), .I (I30014));
INVX1 gate9990(.O (I30017), .I (g22824));
INVX1 gate9991(.O (g23188), .I (I30017));
INVX1 gate9992(.O (I30020), .I (g22519));
INVX1 gate9993(.O (g23189), .I (I30020));
INVX1 gate9994(.O (I30023), .I (g22550));
INVX1 gate9995(.O (g23190), .I (I30023));
INVX1 gate9996(.O (I30026), .I (g22586));
INVX1 gate9997(.O (g23191), .I (I30026));
INVX1 gate9998(.O (I30029), .I (g22642));
INVX1 gate9999(.O (g23192), .I (I30029));
INVX1 gate10000(.O (I30032), .I (g22672));
INVX1 gate10001(.O (g23193), .I (I30032));
INVX1 gate10002(.O (I30035), .I (g22705));
INVX1 gate10003(.O (g23194), .I (I30035));
INVX1 gate10004(.O (I30038), .I (g22673));
INVX1 gate10005(.O (g23195), .I (I30038));
INVX1 gate10006(.O (I30041), .I (g22706));
INVX1 gate10007(.O (g23196), .I (I30041));
INVX1 gate10008(.O (I30044), .I (g22731));
INVX1 gate10009(.O (g23197), .I (I30044));
INVX1 gate10010(.O (I30047), .I (g22107));
INVX1 gate10011(.O (g23198), .I (I30047));
INVX1 gate10012(.O (I30050), .I (g22619));
INVX1 gate10013(.O (g23199), .I (I30050));
INVX1 gate10014(.O (I30053), .I (g22558));
INVX1 gate10015(.O (g23200), .I (I30053));
INVX1 gate10016(.O (I30056), .I (g22589));
INVX1 gate10017(.O (g23201), .I (I30056));
INVX1 gate10018(.O (I30059), .I (g22620));
INVX1 gate10019(.O (g23202), .I (I30059));
INVX1 gate10020(.O (I30062), .I (g22590));
INVX1 gate10021(.O (g23203), .I (I30062));
INVX1 gate10022(.O (I30065), .I (g22621));
INVX1 gate10023(.O (g23204), .I (I30065));
INVX1 gate10024(.O (I30068), .I (g22647));
INVX1 gate10025(.O (g23205), .I (I30068));
INVX1 gate10026(.O (I30071), .I (g22622));
INVX1 gate10027(.O (g23206), .I (I30071));
INVX1 gate10028(.O (I30074), .I (g22648));
INVX1 gate10029(.O (g23207), .I (I30074));
INVX1 gate10030(.O (I30077), .I (g22675));
INVX1 gate10031(.O (g23208), .I (I30077));
INVX1 gate10032(.O (I30080), .I (g22649));
INVX1 gate10033(.O (g23209), .I (I30080));
INVX1 gate10034(.O (I30083), .I (g22676));
INVX1 gate10035(.O (g23210), .I (I30083));
INVX1 gate10036(.O (I30086), .I (g22709));
INVX1 gate10037(.O (g23211), .I (I30086));
INVX1 gate10038(.O (I30089), .I (g22677));
INVX1 gate10039(.O (g23212), .I (I30089));
INVX1 gate10040(.O (I30092), .I (g22710));
INVX1 gate10041(.O (g23213), .I (I30092));
INVX1 gate10042(.O (I30095), .I (g22733));
INVX1 gate10043(.O (g23214), .I (I30095));
INVX1 gate10044(.O (I30098), .I (g22711));
INVX1 gate10045(.O (g23215), .I (I30098));
INVX1 gate10046(.O (I30101), .I (g22734));
INVX1 gate10047(.O (g23216), .I (I30101));
INVX1 gate10048(.O (I30104), .I (g22760));
INVX1 gate10049(.O (g23217), .I (I30104));
INVX1 gate10050(.O (I30107), .I (g22735));
INVX1 gate10051(.O (g23218), .I (I30107));
INVX1 gate10052(.O (I30110), .I (g22761));
INVX1 gate10053(.O (g23219), .I (I30110));
INVX1 gate10054(.O (I30113), .I (g22790));
INVX1 gate10055(.O (g23220), .I (I30113));
INVX1 gate10056(.O (I30116), .I (g22762));
INVX1 gate10057(.O (g23221), .I (I30116));
INVX1 gate10058(.O (I30119), .I (g22791));
INVX1 gate10059(.O (g23222), .I (I30119));
INVX1 gate10060(.O (I30122), .I (g22827));
INVX1 gate10061(.O (g23223), .I (I30122));
INVX1 gate10062(.O (I30125), .I (g22792));
INVX1 gate10063(.O (g23224), .I (I30125));
INVX1 gate10064(.O (I30128), .I (g22828));
INVX1 gate10065(.O (g23225), .I (I30128));
INVX1 gate10066(.O (I30131), .I (g22864));
INVX1 gate10067(.O (g23226), .I (I30131));
INVX1 gate10068(.O (I30134), .I (g22559));
INVX1 gate10069(.O (g23227), .I (I30134));
INVX1 gate10070(.O (I30137), .I (g22591));
INVX1 gate10071(.O (g23228), .I (I30137));
INVX1 gate10072(.O (I30140), .I (g22623));
INVX1 gate10073(.O (g23229), .I (I30140));
INVX1 gate10074(.O (I30143), .I (g22678));
INVX1 gate10075(.O (g23230), .I (I30143));
INVX1 gate10076(.O (I30146), .I (g22712));
INVX1 gate10077(.O (g23231), .I (I30146));
INVX1 gate10078(.O (I30149), .I (g22736));
INVX1 gate10079(.O (g23232), .I (I30149));
INVX1 gate10080(.O (I30152), .I (g22713));
INVX1 gate10081(.O (g23233), .I (I30152));
INVX1 gate10082(.O (I30155), .I (g22737));
INVX1 gate10083(.O (g23234), .I (I30155));
INVX1 gate10084(.O (I30158), .I (g22763));
INVX1 gate10085(.O (g23235), .I (I30158));
INVX1 gate10086(.O (I30161), .I (g22133));
INVX1 gate10087(.O (g23236), .I (I30161));
INVX1 gate10088(.O (I30164), .I (g22655));
INVX1 gate10089(.O (g23237), .I (I30164));
INVX1 gate10090(.O (I30167), .I (g22598));
INVX1 gate10091(.O (g23238), .I (I30167));
INVX1 gate10092(.O (I30170), .I (g22626));
INVX1 gate10093(.O (g23239), .I (I30170));
INVX1 gate10094(.O (I30173), .I (g22656));
INVX1 gate10095(.O (g23240), .I (I30173));
INVX1 gate10096(.O (I30176), .I (g22627));
INVX1 gate10097(.O (g23241), .I (I30176));
INVX1 gate10098(.O (I30179), .I (g22657));
INVX1 gate10099(.O (g23242), .I (I30179));
INVX1 gate10100(.O (I30182), .I (g22683));
INVX1 gate10101(.O (g23243), .I (I30182));
INVX1 gate10102(.O (I30185), .I (g22658));
INVX1 gate10103(.O (g23244), .I (I30185));
INVX1 gate10104(.O (I30188), .I (g22684));
INVX1 gate10105(.O (g23245), .I (I30188));
INVX1 gate10106(.O (I30191), .I (g22715));
INVX1 gate10107(.O (g23246), .I (I30191));
INVX1 gate10108(.O (I30194), .I (g22685));
INVX1 gate10109(.O (g23247), .I (I30194));
INVX1 gate10110(.O (I30197), .I (g22716));
INVX1 gate10111(.O (g23248), .I (I30197));
INVX1 gate10112(.O (I30200), .I (g22740));
INVX1 gate10113(.O (g23249), .I (I30200));
INVX1 gate10114(.O (I30203), .I (g22717));
INVX1 gate10115(.O (g23250), .I (I30203));
INVX1 gate10116(.O (I30206), .I (g22741));
INVX1 gate10117(.O (g23251), .I (I30206));
INVX1 gate10118(.O (I30209), .I (g22765));
INVX1 gate10119(.O (g23252), .I (I30209));
INVX1 gate10120(.O (I30212), .I (g22742));
INVX1 gate10121(.O (g23253), .I (I30212));
INVX1 gate10122(.O (I30215), .I (g22766));
INVX1 gate10123(.O (g23254), .I (I30215));
INVX1 gate10124(.O (I30218), .I (g22794));
INVX1 gate10125(.O (g23255), .I (I30218));
INVX1 gate10126(.O (I30221), .I (g22767));
INVX1 gate10127(.O (g23256), .I (I30221));
INVX1 gate10128(.O (I30224), .I (g22795));
INVX1 gate10129(.O (g23257), .I (I30224));
INVX1 gate10130(.O (I30227), .I (g22832));
INVX1 gate10131(.O (g23258), .I (I30227));
INVX1 gate10132(.O (I30230), .I (g22796));
INVX1 gate10133(.O (g23259), .I (I30230));
INVX1 gate10134(.O (I30233), .I (g22833));
INVX1 gate10135(.O (g23260), .I (I30233));
INVX1 gate10136(.O (I30236), .I (g22866));
INVX1 gate10137(.O (g23261), .I (I30236));
INVX1 gate10138(.O (I30239), .I (g22834));
INVX1 gate10139(.O (g23262), .I (I30239));
INVX1 gate10140(.O (I30242), .I (g22867));
INVX1 gate10141(.O (g23263), .I (I30242));
INVX1 gate10142(.O (I30245), .I (g22899));
INVX1 gate10143(.O (g23264), .I (I30245));
INVX1 gate10144(.O (I30248), .I (g22599));
INVX1 gate10145(.O (g23265), .I (I30248));
INVX1 gate10146(.O (I30251), .I (g22628));
INVX1 gate10147(.O (g23266), .I (I30251));
INVX1 gate10148(.O (I30254), .I (g22659));
INVX1 gate10149(.O (g23267), .I (I30254));
INVX1 gate10150(.O (I30257), .I (g22718));
INVX1 gate10151(.O (g23268), .I (I30257));
INVX1 gate10152(.O (I30260), .I (g22743));
INVX1 gate10153(.O (g23269), .I (I30260));
INVX1 gate10154(.O (I30263), .I (g22768));
INVX1 gate10155(.O (g23270), .I (I30263));
INVX1 gate10156(.O (I30266), .I (g22744));
INVX1 gate10157(.O (g23271), .I (I30266));
INVX1 gate10158(.O (I30269), .I (g22769));
INVX1 gate10159(.O (g23272), .I (I30269));
INVX1 gate10160(.O (I30272), .I (g22797));
INVX1 gate10161(.O (g23273), .I (I30272));
INVX1 gate10162(.O (I30275), .I (g22156));
INVX1 gate10163(.O (g23274), .I (I30275));
INVX1 gate10164(.O (I30278), .I (g22691));
INVX1 gate10165(.O (g23275), .I (I30278));
INVX1 gate10166(.O (I30281), .I (g22635));
INVX1 gate10167(.O (g23276), .I (I30281));
INVX1 gate10168(.O (I30284), .I (g22662));
INVX1 gate10169(.O (g23277), .I (I30284));
INVX1 gate10170(.O (I30287), .I (g22692));
INVX1 gate10171(.O (g23278), .I (I30287));
INVX1 gate10172(.O (I30290), .I (g22663));
INVX1 gate10173(.O (g23279), .I (I30290));
INVX1 gate10174(.O (I30293), .I (g22693));
INVX1 gate10175(.O (g23280), .I (I30293));
INVX1 gate10176(.O (I30296), .I (g22723));
INVX1 gate10177(.O (g23281), .I (I30296));
INVX1 gate10178(.O (I30299), .I (g22694));
INVX1 gate10179(.O (g23282), .I (I30299));
INVX1 gate10180(.O (I30302), .I (g22724));
INVX1 gate10181(.O (g23283), .I (I30302));
INVX1 gate10182(.O (I30305), .I (g22746));
INVX1 gate10183(.O (g23284), .I (I30305));
INVX1 gate10184(.O (I30308), .I (g22725));
INVX1 gate10185(.O (g23285), .I (I30308));
INVX1 gate10186(.O (I30311), .I (g22747));
INVX1 gate10187(.O (g23286), .I (I30311));
INVX1 gate10188(.O (I30314), .I (g22772));
INVX1 gate10189(.O (g23287), .I (I30314));
INVX1 gate10190(.O (I30317), .I (g22748));
INVX1 gate10191(.O (g23288), .I (I30317));
INVX1 gate10192(.O (I30320), .I (g22773));
INVX1 gate10193(.O (g23289), .I (I30320));
INVX1 gate10194(.O (I30323), .I (g22799));
INVX1 gate10195(.O (g23290), .I (I30323));
INVX1 gate10196(.O (I30326), .I (g22774));
INVX1 gate10197(.O (g23291), .I (I30326));
INVX1 gate10198(.O (I30329), .I (g22800));
INVX1 gate10199(.O (g23292), .I (I30329));
INVX1 gate10200(.O (I30332), .I (g22836));
INVX1 gate10201(.O (g23293), .I (I30332));
INVX1 gate10202(.O (I30335), .I (g22801));
INVX1 gate10203(.O (g23294), .I (I30335));
INVX1 gate10204(.O (I30338), .I (g22837));
INVX1 gate10205(.O (g23295), .I (I30338));
INVX1 gate10206(.O (I30341), .I (g22871));
INVX1 gate10207(.O (g23296), .I (I30341));
INVX1 gate10208(.O (I30344), .I (g22838));
INVX1 gate10209(.O (g23297), .I (I30344));
INVX1 gate10210(.O (I30347), .I (g22872));
INVX1 gate10211(.O (g23298), .I (I30347));
INVX1 gate10212(.O (I30350), .I (g22901));
INVX1 gate10213(.O (g23299), .I (I30350));
INVX1 gate10214(.O (I30353), .I (g22873));
INVX1 gate10215(.O (g23300), .I (I30353));
INVX1 gate10216(.O (I30356), .I (g22902));
INVX1 gate10217(.O (g23301), .I (I30356));
INVX1 gate10218(.O (I30359), .I (g22934));
INVX1 gate10219(.O (g23302), .I (I30359));
INVX1 gate10220(.O (I30362), .I (g22636));
INVX1 gate10221(.O (g23303), .I (I30362));
INVX1 gate10222(.O (I30365), .I (g22664));
INVX1 gate10223(.O (g23304), .I (I30365));
INVX1 gate10224(.O (I30368), .I (g22695));
INVX1 gate10225(.O (g23305), .I (I30368));
INVX1 gate10226(.O (I30371), .I (g22749));
INVX1 gate10227(.O (g23306), .I (I30371));
INVX1 gate10228(.O (I30374), .I (g22775));
INVX1 gate10229(.O (g23307), .I (I30374));
INVX1 gate10230(.O (I30377), .I (g22802));
INVX1 gate10231(.O (g23308), .I (I30377));
INVX1 gate10232(.O (I30380), .I (g22776));
INVX1 gate10233(.O (g23309), .I (I30380));
INVX1 gate10234(.O (I30383), .I (g22803));
INVX1 gate10235(.O (g23310), .I (I30383));
INVX1 gate10236(.O (I30386), .I (g22839));
INVX1 gate10237(.O (g23311), .I (I30386));
INVX1 gate10238(.O (I30389), .I (g22225));
INVX1 gate10239(.O (g23312), .I (I30389));
INVX1 gate10240(.O (I30392), .I (g22226));
INVX1 gate10241(.O (g23313), .I (I30392));
INVX1 gate10242(.O (I30395), .I (g22253));
INVX1 gate10243(.O (g23314), .I (I30395));
INVX1 gate10244(.O (I30398), .I (g22840));
INVX1 gate10245(.O (g23315), .I (I30398));
INVX1 gate10246(.O (I30401), .I (g22444));
INVX1 gate10247(.O (g23316), .I (I30401));
INVX1 gate10248(.O (I30404), .I (g22948));
INVX1 gate10249(.O (g23317), .I (I30404));
INVX1 gate10250(.O (I30407), .I (g22970));
INVX1 gate10251(.O (g23318), .I (I30407));
INVX1 gate10252(.O (g23403), .I (g23052));
INVX1 gate10253(.O (g23410), .I (g23071));
INVX1 gate10254(.O (g23415), .I (g23084));
INVX1 gate10255(.O (g23420), .I (g23089));
INVX1 gate10256(.O (g23424), .I (g23100));
INVX1 gate10257(.O (g23429), .I (g23107));
INVX1 gate10258(.O (g23435), .I (g23120));
INVX1 gate10259(.O (I30467), .I (g23000));
INVX1 gate10260(.O (g23438), .I (I30467));
INVX1 gate10261(.O (I30470), .I (g23117));
INVX1 gate10262(.O (g23439), .I (I30470));
INVX1 gate10263(.O (g23441), .I (g23129));
INVX1 gate10264(.O (g23444), .I (g22945));
INVX1 gate10265(.O (I30476), .I (g22876));
INVX1 gate10266(.O (g23448), .I (I30476));
INVX1 gate10267(.O (I30480), .I (g23014));
INVX1 gate10268(.O (g23452), .I (I30480));
INVX1 gate10269(.O (I30483), .I (g23126));
INVX1 gate10270(.O (g23453), .I (I30483));
INVX1 gate10271(.O (I30486), .I (g23022));
INVX1 gate10272(.O (g23454), .I (I30486));
INVX1 gate10273(.O (I30489), .I (g22911));
INVX1 gate10274(.O (g23455), .I (I30489));
INVX1 gate10275(.O (I30493), .I (g23030));
INVX1 gate10276(.O (g23459), .I (I30493));
INVX1 gate10277(.O (I30496), .I (g23137));
INVX1 gate10278(.O (g23460), .I (I30496));
INVX1 gate10279(.O (I30501), .I (g23039));
INVX1 gate10280(.O (g23463), .I (I30501));
INVX1 gate10281(.O (I30504), .I (g22936));
INVX1 gate10282(.O (g23464), .I (I30504));
INVX1 gate10283(.O (I30508), .I (g23047));
INVX1 gate10284(.O (g23468), .I (I30508));
INVX1 gate10285(.O (I30511), .I (g21970));
INVX1 gate10286(.O (g23469), .I (I30511));
INVX1 gate10287(.O (g23470), .I (g22188));
INVX1 gate10288(.O (I30516), .I (g23058));
INVX1 gate10289(.O (g23472), .I (I30516));
INVX1 gate10290(.O (I30519), .I (g22942));
INVX1 gate10291(.O (g23473), .I (I30519));
INVX1 gate10292(.O (I30525), .I (g23067));
INVX1 gate10293(.O (g23481), .I (I30525));
INVX1 gate10294(.O (g23482), .I (g22197));
INVX1 gate10295(.O (I30531), .I (g23076));
INVX1 gate10296(.O (g23485), .I (I30531));
INVX1 gate10297(.O (I30536), .I (g23081));
INVX1 gate10298(.O (g23492), .I (I30536));
INVX1 gate10299(.O (g23493), .I (g22203));
INVX1 gate10300(.O (I30544), .I (g23092));
INVX1 gate10301(.O (g23500), .I (I30544));
INVX1 gate10302(.O (I30547), .I (g23093));
INVX1 gate10303(.O (g23501), .I (I30547));
INVX1 gate10304(.O (I30552), .I (g23097));
INVX1 gate10305(.O (g23508), .I (I30552));
INVX1 gate10306(.O (g23509), .I (g22209));
INVX1 gate10307(.O (I30560), .I (g23110));
INVX1 gate10308(.O (g23516), .I (I30560));
INVX1 gate10309(.O (I30563), .I (g23111));
INVX1 gate10310(.O (g23517), .I (I30563));
INVX1 gate10311(.O (I30568), .I (g23114));
INVX1 gate10312(.O (g23524), .I (I30568));
INVX1 gate10313(.O (I30575), .I (g23123));
INVX1 gate10314(.O (g23531), .I (I30575));
INVX1 gate10315(.O (I30578), .I (g23124));
INVX1 gate10316(.O (g23532), .I (I30578));
INVX1 gate10317(.O (I30586), .I (g23132));
INVX1 gate10318(.O (g23542), .I (I30586));
INVX1 gate10319(.O (I30589), .I (g23133));
INVX1 gate10320(.O (g23543), .I (I30589));
INVX1 gate10321(.O (I30594), .I (g22025));
INVX1 gate10322(.O (g23546), .I (I30594));
INVX1 gate10323(.O (I30598), .I (g22027));
INVX1 gate10324(.O (g23548), .I (I30598));
INVX1 gate10325(.O (I30601), .I (g22028));
INVX1 gate10326(.O (g23549), .I (I30601));
INVX1 gate10327(.O (I30607), .I (g22029));
INVX1 gate10328(.O (g23553), .I (I30607));
INVX1 gate10329(.O (I30611), .I (g22030));
INVX1 gate10330(.O (g23555), .I (I30611));
INVX1 gate10331(.O (I30614), .I (g22031));
INVX1 gate10332(.O (g23556), .I (I30614));
INVX1 gate10333(.O (I30617), .I (g22032));
INVX1 gate10334(.O (g23557), .I (I30617));
INVX1 gate10335(.O (I30623), .I (g22033));
INVX1 gate10336(.O (g23561), .I (I30623));
INVX1 gate10337(.O (I30626), .I (g22034));
INVX1 gate10338(.O (g23562), .I (I30626));
INVX1 gate10339(.O (I30632), .I (g22035));
INVX1 gate10340(.O (g23566), .I (I30632));
INVX1 gate10341(.O (I30636), .I (g22037));
INVX1 gate10342(.O (g23568), .I (I30636));
INVX1 gate10343(.O (I30639), .I (g22038));
INVX1 gate10344(.O (g23569), .I (I30639));
INVX1 gate10345(.O (I30642), .I (g22039));
INVX1 gate10346(.O (g23570), .I (I30642));
INVX1 gate10347(.O (I30648), .I (g22040));
INVX1 gate10348(.O (g23574), .I (I30648));
INVX1 gate10349(.O (I30651), .I (g22041));
INVX1 gate10350(.O (g23575), .I (I30651));
INVX1 gate10351(.O (I30654), .I (g22042));
INVX1 gate10352(.O (g23576), .I (I30654));
INVX1 gate10353(.O (I30660), .I (g22043));
INVX1 gate10354(.O (g23580), .I (I30660));
INVX1 gate10355(.O (I30663), .I (g22044));
INVX1 gate10356(.O (g23581), .I (I30663));
INVX1 gate10357(.O (I30669), .I (g22045));
INVX1 gate10358(.O (g23585), .I (I30669));
INVX1 gate10359(.O (I30673), .I (g22047));
INVX1 gate10360(.O (g23587), .I (I30673));
INVX1 gate10361(.O (I30676), .I (g22048));
INVX1 gate10362(.O (g23588), .I (I30676));
INVX1 gate10363(.O (I30679), .I (g22049));
INVX1 gate10364(.O (g23589), .I (I30679));
INVX1 gate10365(.O (I30686), .I (g23136));
INVX1 gate10366(.O (g23594), .I (I30686));
INVX1 gate10367(.O (I30689), .I (g22054));
INVX1 gate10368(.O (g23595), .I (I30689));
INVX1 gate10369(.O (I30692), .I (g22055));
INVX1 gate10370(.O (g23596), .I (I30692));
INVX1 gate10371(.O (I30695), .I (g22056));
INVX1 gate10372(.O (g23597), .I (I30695));
INVX1 gate10373(.O (I30701), .I (g22057));
INVX1 gate10374(.O (g23601), .I (I30701));
INVX1 gate10375(.O (I30704), .I (g22058));
INVX1 gate10376(.O (g23602), .I (I30704));
INVX1 gate10377(.O (I30707), .I (g22059));
INVX1 gate10378(.O (g23603), .I (I30707));
INVX1 gate10379(.O (I30713), .I (g22060));
INVX1 gate10380(.O (g23607), .I (I30713));
INVX1 gate10381(.O (I30716), .I (g22061));
INVX1 gate10382(.O (g23608), .I (I30716));
INVX1 gate10383(.O (I30722), .I (g22063));
INVX1 gate10384(.O (g23612), .I (I30722));
INVX1 gate10385(.O (I30725), .I (g22064));
INVX1 gate10386(.O (g23613), .I (I30725));
INVX1 gate10387(.O (I30728), .I (g22065));
INVX1 gate10388(.O (g23614), .I (I30728));
INVX1 gate10389(.O (I30735), .I (g22066));
INVX1 gate10390(.O (g23619), .I (I30735));
INVX1 gate10391(.O (I30738), .I (g22067));
INVX1 gate10392(.O (g23620), .I (I30738));
INVX1 gate10393(.O (I30741), .I (g22068));
INVX1 gate10394(.O (g23621), .I (I30741));
INVX1 gate10395(.O (I30748), .I (g21969));
INVX1 gate10396(.O (g23626), .I (I30748));
INVX1 gate10397(.O (I30751), .I (g22073));
INVX1 gate10398(.O (g23627), .I (I30751));
INVX1 gate10399(.O (I30754), .I (g22074));
INVX1 gate10400(.O (g23628), .I (I30754));
INVX1 gate10401(.O (I30757), .I (g22075));
INVX1 gate10402(.O (g23629), .I (I30757));
INVX1 gate10403(.O (I30763), .I (g22076));
INVX1 gate10404(.O (g23633), .I (I30763));
INVX1 gate10405(.O (I30766), .I (g22077));
INVX1 gate10406(.O (g23634), .I (I30766));
INVX1 gate10407(.O (I30769), .I (g22078));
INVX1 gate10408(.O (g23635), .I (I30769));
INVX1 gate10409(.O (I30776), .I (g22079));
INVX1 gate10410(.O (g23640), .I (I30776));
INVX1 gate10411(.O (I30779), .I (g22080));
INVX1 gate10412(.O (g23641), .I (I30779));
INVX1 gate10413(.O (I30782), .I (g22081));
INVX1 gate10414(.O (g23642), .I (I30782));
INVX1 gate10415(.O (I30786), .I (g22454));
INVX1 gate10416(.O (g23644), .I (I30786));
INVX1 gate10417(.O (I30797), .I (g22087));
INVX1 gate10418(.O (g23661), .I (I30797));
INVX1 gate10419(.O (I30800), .I (g22088));
INVX1 gate10420(.O (g23662), .I (I30800));
INVX1 gate10421(.O (I30803), .I (g22089));
INVX1 gate10422(.O (g23663), .I (I30803));
INVX1 gate10423(.O (I30810), .I (g22090));
INVX1 gate10424(.O (g23668), .I (I30810));
INVX1 gate10425(.O (I30813), .I (g22091));
INVX1 gate10426(.O (g23669), .I (I30813));
INVX1 gate10427(.O (I30816), .I (g22092));
INVX1 gate10428(.O (g23670), .I (I30816));
INVX1 gate10429(.O (I30823), .I (g21972));
INVX1 gate10430(.O (g23675), .I (I30823));
INVX1 gate10431(.O (I30826), .I (g22097));
INVX1 gate10432(.O (g23676), .I (I30826));
INVX1 gate10433(.O (I30829), .I (g22098));
INVX1 gate10434(.O (g23677), .I (I30829));
INVX1 gate10435(.O (I30832), .I (g22099));
INVX1 gate10436(.O (g23678), .I (I30832));
INVX1 gate10437(.O (I30838), .I (g22100));
INVX1 gate10438(.O (g23682), .I (I30838));
INVX1 gate10439(.O (I30841), .I (g22101));
INVX1 gate10440(.O (g23683), .I (I30841));
INVX1 gate10441(.O (I30844), .I (g22102));
INVX1 gate10442(.O (g23684), .I (I30844));
INVX1 gate10443(.O (I30847), .I (g22103));
INVX1 gate10444(.O (g23685), .I (I30847));
INVX1 gate10445(.O (I30854), .I (g22104));
INVX1 gate10446(.O (g23690), .I (I30854));
INVX1 gate10447(.O (I30857), .I (g22105));
INVX1 gate10448(.O (g23691), .I (I30857));
INVX1 gate10449(.O (I30860), .I (g22106));
INVX1 gate10450(.O (g23692), .I (I30860));
INVX1 gate10451(.O (I30864), .I (g22493));
INVX1 gate10452(.O (g23694), .I (I30864));
INVX1 gate10453(.O (I30875), .I (g22112));
INVX1 gate10454(.O (g23711), .I (I30875));
INVX1 gate10455(.O (I30878), .I (g22113));
INVX1 gate10456(.O (g23712), .I (I30878));
INVX1 gate10457(.O (I30881), .I (g22114));
INVX1 gate10458(.O (g23713), .I (I30881));
INVX1 gate10459(.O (I30888), .I (g22115));
INVX1 gate10460(.O (g23718), .I (I30888));
INVX1 gate10461(.O (I30891), .I (g22116));
INVX1 gate10462(.O (g23719), .I (I30891));
INVX1 gate10463(.O (I30894), .I (g22117));
INVX1 gate10464(.O (g23720), .I (I30894));
INVX1 gate10465(.O (I30901), .I (g21974));
INVX1 gate10466(.O (g23725), .I (I30901));
INVX1 gate10467(.O (I30905), .I (g22122));
INVX1 gate10468(.O (g23727), .I (I30905));
INVX1 gate10469(.O (I30908), .I (g22123));
INVX1 gate10470(.O (g23728), .I (I30908));
INVX1 gate10471(.O (I30911), .I (g22124));
INVX1 gate10472(.O (g23729), .I (I30911));
INVX1 gate10473(.O (I30914), .I (g22125));
INVX1 gate10474(.O (g23730), .I (I30914));
INVX1 gate10475(.O (I30917), .I (g22806));
INVX1 gate10476(.O (g23731), .I (I30917));
INVX1 gate10477(.O (I30922), .I (g22126));
INVX1 gate10478(.O (g23736), .I (I30922));
INVX1 gate10479(.O (I30925), .I (g22127));
INVX1 gate10480(.O (g23737), .I (I30925));
INVX1 gate10481(.O (I30928), .I (g22128));
INVX1 gate10482(.O (g23738), .I (I30928));
INVX1 gate10483(.O (I30931), .I (g22129));
INVX1 gate10484(.O (g23739), .I (I30931));
INVX1 gate10485(.O (I30938), .I (g22130));
INVX1 gate10486(.O (g23744), .I (I30938));
INVX1 gate10487(.O (I30941), .I (g22131));
INVX1 gate10488(.O (g23745), .I (I30941));
INVX1 gate10489(.O (I30944), .I (g22132));
INVX1 gate10490(.O (g23746), .I (I30944));
INVX1 gate10491(.O (I30948), .I (g22536));
INVX1 gate10492(.O (g23748), .I (I30948));
INVX1 gate10493(.O (I30959), .I (g22138));
INVX1 gate10494(.O (g23765), .I (I30959));
INVX1 gate10495(.O (I30962), .I (g22139));
INVX1 gate10496(.O (g23766), .I (I30962));
INVX1 gate10497(.O (I30965), .I (g22140));
INVX1 gate10498(.O (g23767), .I (I30965));
INVX1 gate10499(.O (I30973), .I (g22141));
INVX1 gate10500(.O (g23773), .I (I30973));
INVX1 gate10501(.O (I30976), .I (g22142));
INVX1 gate10502(.O (g23774), .I (I30976));
INVX1 gate10503(.O (I30979), .I (g22143));
INVX1 gate10504(.O (g23775), .I (I30979));
INVX1 gate10505(.O (I30985), .I (g22992));
INVX1 gate10506(.O (g23779), .I (I30985));
INVX1 gate10507(.O (I30988), .I (g22145));
INVX1 gate10508(.O (g23782), .I (I30988));
INVX1 gate10509(.O (I30991), .I (g22146));
INVX1 gate10510(.O (g23783), .I (I30991));
INVX1 gate10511(.O (I30994), .I (g22147));
INVX1 gate10512(.O (g23784), .I (I30994));
INVX1 gate10513(.O (I30997), .I (g22148));
INVX1 gate10514(.O (g23785), .I (I30997));
INVX1 gate10515(.O (I31000), .I (g22847));
INVX1 gate10516(.O (g23786), .I (I31000));
INVX1 gate10517(.O (I31005), .I (g22149));
INVX1 gate10518(.O (g23791), .I (I31005));
INVX1 gate10519(.O (I31008), .I (g22150));
INVX1 gate10520(.O (g23792), .I (I31008));
INVX1 gate10521(.O (I31011), .I (g22151));
INVX1 gate10522(.O (g23793), .I (I31011));
INVX1 gate10523(.O (I31014), .I (g22152));
INVX1 gate10524(.O (g23794), .I (I31014));
INVX1 gate10525(.O (I31021), .I (g22153));
INVX1 gate10526(.O (g23799), .I (I31021));
INVX1 gate10527(.O (I31024), .I (g22154));
INVX1 gate10528(.O (g23800), .I (I31024));
INVX1 gate10529(.O (I31027), .I (g22155));
INVX1 gate10530(.O (g23801), .I (I31027));
INVX1 gate10531(.O (I31031), .I (g22576));
INVX1 gate10532(.O (g23803), .I (I31031));
INVX1 gate10533(.O (I31043), .I (g22161));
INVX1 gate10534(.O (g23821), .I (I31043));
INVX1 gate10535(.O (I31050), .I (g22162));
INVX1 gate10536(.O (g23826), .I (I31050));
INVX1 gate10537(.O (I31053), .I (g22163));
INVX1 gate10538(.O (g23827), .I (I31053));
INVX1 gate10539(.O (I31056), .I (g22164));
INVX1 gate10540(.O (g23828), .I (I31056));
INVX1 gate10541(.O (I31062), .I (g23003));
INVX1 gate10542(.O (g23832), .I (I31062));
INVX1 gate10543(.O (I31065), .I (g22166));
INVX1 gate10544(.O (g23835), .I (I31065));
INVX1 gate10545(.O (I31068), .I (g22167));
INVX1 gate10546(.O (g23836), .I (I31068));
INVX1 gate10547(.O (I31071), .I (g22168));
INVX1 gate10548(.O (g23837), .I (I31071));
INVX1 gate10549(.O (I31074), .I (g22169));
INVX1 gate10550(.O (g23838), .I (I31074));
INVX1 gate10551(.O (I31077), .I (g22882));
INVX1 gate10552(.O (g23839), .I (I31077));
INVX1 gate10553(.O (I31082), .I (g22170));
INVX1 gate10554(.O (g23844), .I (I31082));
INVX1 gate10555(.O (I31085), .I (g22171));
INVX1 gate10556(.O (g23845), .I (I31085));
INVX1 gate10557(.O (I31088), .I (g22172));
INVX1 gate10558(.O (g23846), .I (I31088));
INVX1 gate10559(.O (I31091), .I (g22173));
INVX1 gate10560(.O (g23847), .I (I31091));
INVX1 gate10561(.O (g23853), .I (g22300));
INVX1 gate10562(.O (I31102), .I (g22177));
INVX1 gate10563(.O (g23856), .I (I31102));
INVX1 gate10564(.O (I31109), .I (g22178));
INVX1 gate10565(.O (g23861), .I (I31109));
INVX1 gate10566(.O (I31112), .I (g22179));
INVX1 gate10567(.O (g23862), .I (I31112));
INVX1 gate10568(.O (I31115), .I (g22180));
INVX1 gate10569(.O (g23863), .I (I31115));
INVX1 gate10570(.O (I31121), .I (g23017));
INVX1 gate10571(.O (g23867), .I (I31121));
INVX1 gate10572(.O (I31124), .I (g22182));
INVX1 gate10573(.O (g23870), .I (I31124));
INVX1 gate10574(.O (I31127), .I (g22183));
INVX1 gate10575(.O (g23871), .I (I31127));
INVX1 gate10576(.O (I31130), .I (g22184));
INVX1 gate10577(.O (g23872), .I (I31130));
INVX1 gate10578(.O (I31133), .I (g22185));
INVX1 gate10579(.O (g23873), .I (I31133));
INVX1 gate10580(.O (I31136), .I (g22917));
INVX1 gate10581(.O (g23874), .I (I31136));
INVX1 gate10582(.O (I31141), .I (g22777));
INVX1 gate10583(.O (g23879), .I (I31141));
INVX1 gate10584(.O (I31144), .I (g22935));
INVX1 gate10585(.O (g23882), .I (I31144));
INVX1 gate10586(.O (g23885), .I (g22062));
INVX1 gate10587(.O (g23887), .I (g22328));
INVX1 gate10588(.O (I31152), .I (g22191));
INVX1 gate10589(.O (g23890), .I (I31152));
INVX1 gate10590(.O (I31159), .I (g22192));
INVX1 gate10591(.O (g23895), .I (I31159));
INVX1 gate10592(.O (I31162), .I (g22193));
INVX1 gate10593(.O (g23896), .I (I31162));
INVX1 gate10594(.O (I31165), .I (g22194));
INVX1 gate10595(.O (g23897), .I (I31165));
INVX1 gate10596(.O (I31171), .I (g23033));
INVX1 gate10597(.O (g23901), .I (I31171));
INVX1 gate10598(.O (g23905), .I (g22046));
INVX1 gate10599(.O (g23908), .I (g22353));
INVX1 gate10600(.O (I31181), .I (g22200));
INVX1 gate10601(.O (g23911), .I (I31181));
INVX1 gate10602(.O (I31188), .I (g21989));
INVX1 gate10603(.O (g23916), .I (I31188));
INVX1 gate10604(.O (g23918), .I (g22036));
INVX1 gate10605(.O (I31195), .I (g22578));
INVX1 gate10606(.O (g23923), .I (I31195));
INVX1 gate10607(.O (g23940), .I (g22376));
INVX1 gate10608(.O (I31205), .I (g22002));
INVX1 gate10609(.O (g23943), .I (I31205));
INVX1 gate10610(.O (I31213), .I (g22615));
INVX1 gate10611(.O (g23955), .I (I31213));
INVX1 gate10612(.O (I31226), .I (g22651));
INVX1 gate10613(.O (g23984), .I (I31226));
INVX1 gate10614(.O (I31232), .I (g22026));
INVX1 gate10615(.O (g24000), .I (I31232));
INVX1 gate10616(.O (I31235), .I (g22218));
INVX1 gate10617(.O (g24001), .I (I31235));
INVX1 gate10618(.O (I31244), .I (g22687));
INVX1 gate10619(.O (g24014), .I (I31244));
INVX1 gate10620(.O (I31250), .I (g22953));
INVX1 gate10621(.O (g24030), .I (I31250));
INVX1 gate10622(.O (I31253), .I (g22231));
INVX1 gate10623(.O (g24033), .I (I31253));
INVX1 gate10624(.O (I31257), .I (g22234));
INVX1 gate10625(.O (g24035), .I (I31257));
INVX1 gate10626(.O (g24047), .I (g23023));
INVX1 gate10627(.O (I31266), .I (g22242));
INVX1 gate10628(.O (g24051), .I (I31266));
INVX1 gate10629(.O (I31270), .I (g22247));
INVX1 gate10630(.O (g24053), .I (I31270));
INVX1 gate10631(.O (I31274), .I (g22249));
INVX1 gate10632(.O (g24055), .I (I31274));
INVX1 gate10633(.O (g24060), .I (g23040));
INVX1 gate10634(.O (I31282), .I (g22263));
INVX1 gate10635(.O (g24064), .I (I31282));
INVX1 gate10636(.O (I31286), .I (g22267));
INVX1 gate10637(.O (g24066), .I (I31286));
INVX1 gate10638(.O (I31290), .I (g22269));
INVX1 gate10639(.O (g24068), .I (I31290));
INVX1 gate10640(.O (g24073), .I (g23059));
INVX1 gate10641(.O (I31298), .I (g22280));
INVX1 gate10642(.O (g24077), .I (I31298));
INVX1 gate10643(.O (I31302), .I (g22284));
INVX1 gate10644(.O (g24079), .I (I31302));
INVX1 gate10645(.O (g24084), .I (g23077));
INVX1 gate10646(.O (I31310), .I (g22299));
INVX1 gate10647(.O (g24088), .I (I31310));
INVX1 gate10648(.O (g24094), .I (g22339));
INVX1 gate10649(.O (g24095), .I (g22362));
INVX1 gate10650(.O (g24096), .I (g22405));
INVX1 gate10651(.O (g24097), .I (g22382));
INVX1 gate10652(.O (g24098), .I (g22409));
INVX1 gate10653(.O (g24099), .I (g22412));
INVX1 gate10654(.O (g24101), .I (g22415));
INVX1 gate10655(.O (g24102), .I (g22418));
INVX1 gate10656(.O (g24103), .I (g22397));
INVX1 gate10657(.O (g24104), .I (g22422));
INVX1 gate10658(.O (g24105), .I (g22425));
INVX1 gate10659(.O (g24106), .I (g22428));
INVX1 gate10660(.O (g24107), .I (g22431));
INVX1 gate10661(.O (g24108), .I (g22434));
INVX1 gate10662(.O (g24110), .I (g22437));
INVX1 gate10663(.O (g24111), .I (g22440));
INVX1 gate10664(.O (g24112), .I (g22445));
INVX1 gate10665(.O (g24113), .I (g22448));
INVX1 gate10666(.O (g24114), .I (g22451));
INVX1 gate10667(.O (g24115), .I (g22381));
INVX1 gate10668(.O (g24121), .I (g22455));
INVX1 gate10669(.O (g24122), .I (g22458));
INVX1 gate10670(.O (g24123), .I (g22461));
INVX1 gate10671(.O (g24124), .I (g22464));
INVX1 gate10672(.O (g24125), .I (g22467));
INVX1 gate10673(.O (g24127), .I (g22470));
INVX1 gate10674(.O (g24128), .I (g22473));
INVX1 gate10675(.O (g24129), .I (g22477));
INVX1 gate10676(.O (g24130), .I (g22480));
INVX1 gate10677(.O (g24131), .I (g22484));
INVX1 gate10678(.O (g24132), .I (g22487));
INVX1 gate10679(.O (g24133), .I (g22490));
INVX1 gate10680(.O (g24134), .I (g22396));
INVX1 gate10681(.O (g24140), .I (g22494));
INVX1 gate10682(.O (g24141), .I (g22497));
INVX1 gate10683(.O (g24142), .I (g22500));
INVX1 gate10684(.O (g24143), .I (g22503));
INVX1 gate10685(.O (g24144), .I (g22506));
INVX1 gate10686(.O (g24146), .I (g22509));
INVX1 gate10687(.O (g24147), .I (g22512));
INVX1 gate10688(.O (g24148), .I (g22520));
INVX1 gate10689(.O (g24149), .I (g22523));
INVX1 gate10690(.O (g24150), .I (g22527));
INVX1 gate10691(.O (g24151), .I (g22530));
INVX1 gate10692(.O (g24152), .I (g22533));
INVX1 gate10693(.O (g24153), .I (g22399));
INVX1 gate10694(.O (g24159), .I (g22537));
INVX1 gate10695(.O (g24160), .I (g22540));
INVX1 gate10696(.O (g24161), .I (g22543));
INVX1 gate10697(.O (g24162), .I (g22552));
INVX1 gate10698(.O (g24163), .I (g22560));
INVX1 gate10699(.O (g24164), .I (g22563));
INVX1 gate10700(.O (g24165), .I (g22567));
INVX1 gate10701(.O (g24166), .I (g22570));
INVX1 gate10702(.O (g24167), .I (g22573));
INVX1 gate10703(.O (g24168), .I (g22400));
INVX1 gate10704(.O (g24175), .I (g22592));
INVX1 gate10705(.O (g24176), .I (g22600));
INVX1 gate10706(.O (g24177), .I (g22603));
INVX1 gate10707(.O (g24180), .I (g22629));
INVX1 gate10708(.O (I31387), .I (g22811));
INVX1 gate10709(.O (g24183), .I (I31387));
INVX1 gate10710(.O (g24210), .I (g22696));
INVX1 gate10711(.O (g24220), .I (g22750));
INVX1 gate10712(.O (I31417), .I (g22578));
INVX1 gate10713(.O (g24233), .I (I31417));
INVX1 gate10714(.O (I31426), .I (g22615));
INVX1 gate10715(.O (g24240), .I (I31426));
INVX1 gate10716(.O (I31436), .I (g22651));
INVX1 gate10717(.O (g24248), .I (I31436));
INVX1 gate10718(.O (g24251), .I (g22903));
INVX1 gate10719(.O (I31445), .I (g22687));
INVX1 gate10720(.O (g24255), .I (I31445));
INVX1 gate10721(.O (I31451), .I (g23682));
INVX1 gate10722(.O (g24259), .I (I31451));
INVX1 gate10723(.O (I31454), .I (g23727));
INVX1 gate10724(.O (g24260), .I (I31454));
INVX1 gate10725(.O (I31457), .I (g23773));
INVX1 gate10726(.O (g24261), .I (I31457));
INVX1 gate10727(.O (I31460), .I (g23728));
INVX1 gate10728(.O (g24262), .I (I31460));
INVX1 gate10729(.O (I31463), .I (g23774));
INVX1 gate10730(.O (g24263), .I (I31463));
INVX1 gate10731(.O (I31466), .I (g23821));
INVX1 gate10732(.O (g24264), .I (I31466));
INVX1 gate10733(.O (I31469), .I (g23546));
INVX1 gate10734(.O (g24265), .I (I31469));
INVX1 gate10735(.O (I31472), .I (g23548));
INVX1 gate10736(.O (g24266), .I (I31472));
INVX1 gate10737(.O (I31475), .I (g23555));
INVX1 gate10738(.O (g24267), .I (I31475));
INVX1 gate10739(.O (I31478), .I (g23549));
INVX1 gate10740(.O (g24268), .I (I31478));
INVX1 gate10741(.O (I31481), .I (g23556));
INVX1 gate10742(.O (g24269), .I (I31481));
INVX1 gate10743(.O (I31484), .I (g23568));
INVX1 gate10744(.O (g24270), .I (I31484));
INVX1 gate10745(.O (I31487), .I (g23557));
INVX1 gate10746(.O (g24271), .I (I31487));
INVX1 gate10747(.O (I31490), .I (g23569));
INVX1 gate10748(.O (g24272), .I (I31490));
INVX1 gate10749(.O (I31493), .I (g23587));
INVX1 gate10750(.O (g24273), .I (I31493));
INVX1 gate10751(.O (I31496), .I (g23570));
INVX1 gate10752(.O (g24274), .I (I31496));
INVX1 gate10753(.O (I31499), .I (g23588));
INVX1 gate10754(.O (g24275), .I (I31499));
INVX1 gate10755(.O (I31502), .I (g23612));
INVX1 gate10756(.O (g24276), .I (I31502));
INVX1 gate10757(.O (I31505), .I (g23589));
INVX1 gate10758(.O (g24277), .I (I31505));
INVX1 gate10759(.O (I31508), .I (g23613));
INVX1 gate10760(.O (g24278), .I (I31508));
INVX1 gate10761(.O (I31511), .I (g23640));
INVX1 gate10762(.O (g24279), .I (I31511));
INVX1 gate10763(.O (I31514), .I (g23614));
INVX1 gate10764(.O (g24280), .I (I31514));
INVX1 gate10765(.O (I31517), .I (g23641));
INVX1 gate10766(.O (g24281), .I (I31517));
INVX1 gate10767(.O (I31520), .I (g23683));
INVX1 gate10768(.O (g24282), .I (I31520));
INVX1 gate10769(.O (I31523), .I (g23642));
INVX1 gate10770(.O (g24283), .I (I31523));
INVX1 gate10771(.O (I31526), .I (g23684));
INVX1 gate10772(.O (g24284), .I (I31526));
INVX1 gate10773(.O (I31529), .I (g23729));
INVX1 gate10774(.O (g24285), .I (I31529));
INVX1 gate10775(.O (I31532), .I (g23685));
INVX1 gate10776(.O (g24286), .I (I31532));
INVX1 gate10777(.O (I31535), .I (g23730));
INVX1 gate10778(.O (g24287), .I (I31535));
INVX1 gate10779(.O (I31538), .I (g23775));
INVX1 gate10780(.O (g24288), .I (I31538));
INVX1 gate10781(.O (I31541), .I (g23500));
INVX1 gate10782(.O (g24289), .I (I31541));
INVX1 gate10783(.O (I31544), .I (g23438));
INVX1 gate10784(.O (g24290), .I (I31544));
INVX1 gate10785(.O (I31547), .I (g23454));
INVX1 gate10786(.O (g24291), .I (I31547));
INVX1 gate10787(.O (I31550), .I (g23481));
INVX1 gate10788(.O (g24292), .I (I31550));
INVX1 gate10789(.O (I31553), .I (g23501));
INVX1 gate10790(.O (g24293), .I (I31553));
INVX1 gate10791(.O (I31556), .I (g23439));
INVX1 gate10792(.O (g24294), .I (I31556));
INVX1 gate10793(.O (I31559), .I (g24233));
INVX1 gate10794(.O (g24295), .I (I31559));
INVX1 gate10795(.O (I31562), .I (g23594));
INVX1 gate10796(.O (g24296), .I (I31562));
INVX1 gate10797(.O (I31565), .I (g24001));
INVX1 gate10798(.O (g24297), .I (I31565));
INVX1 gate10799(.O (I31568), .I (g24033));
INVX1 gate10800(.O (g24298), .I (I31568));
INVX1 gate10801(.O (I31571), .I (g24051));
INVX1 gate10802(.O (g24299), .I (I31571));
INVX1 gate10803(.O (I31574), .I (g23736));
INVX1 gate10804(.O (g24300), .I (I31574));
INVX1 gate10805(.O (I31577), .I (g23782));
INVX1 gate10806(.O (g24301), .I (I31577));
INVX1 gate10807(.O (I31580), .I (g23826));
INVX1 gate10808(.O (g24302), .I (I31580));
INVX1 gate10809(.O (I31583), .I (g23783));
INVX1 gate10810(.O (g24303), .I (I31583));
INVX1 gate10811(.O (I31586), .I (g23827));
INVX1 gate10812(.O (g24304), .I (I31586));
INVX1 gate10813(.O (I31589), .I (g23856));
INVX1 gate10814(.O (g24305), .I (I31589));
INVX1 gate10815(.O (I31592), .I (g23553));
INVX1 gate10816(.O (g24306), .I (I31592));
INVX1 gate10817(.O (I31595), .I (g23561));
INVX1 gate10818(.O (g24307), .I (I31595));
INVX1 gate10819(.O (I31598), .I (g23574));
INVX1 gate10820(.O (g24308), .I (I31598));
INVX1 gate10821(.O (I31601), .I (g23562));
INVX1 gate10822(.O (g24309), .I (I31601));
INVX1 gate10823(.O (I31604), .I (g23575));
INVX1 gate10824(.O (g24310), .I (I31604));
INVX1 gate10825(.O (I31607), .I (g23595));
INVX1 gate10826(.O (g24311), .I (I31607));
INVX1 gate10827(.O (I31610), .I (g23576));
INVX1 gate10828(.O (g24312), .I (I31610));
INVX1 gate10829(.O (I31613), .I (g23596));
INVX1 gate10830(.O (g24313), .I (I31613));
INVX1 gate10831(.O (I31616), .I (g23619));
INVX1 gate10832(.O (g24314), .I (I31616));
INVX1 gate10833(.O (I31619), .I (g23597));
INVX1 gate10834(.O (g24315), .I (I31619));
INVX1 gate10835(.O (I31622), .I (g23620));
INVX1 gate10836(.O (g24316), .I (I31622));
INVX1 gate10837(.O (I31625), .I (g23661));
INVX1 gate10838(.O (g24317), .I (I31625));
INVX1 gate10839(.O (I31628), .I (g23621));
INVX1 gate10840(.O (g24318), .I (I31628));
INVX1 gate10841(.O (I31631), .I (g23662));
INVX1 gate10842(.O (g24319), .I (I31631));
INVX1 gate10843(.O (I31634), .I (g23690));
INVX1 gate10844(.O (g24320), .I (I31634));
INVX1 gate10845(.O (I31637), .I (g23663));
INVX1 gate10846(.O (g24321), .I (I31637));
INVX1 gate10847(.O (I31640), .I (g23691));
INVX1 gate10848(.O (g24322), .I (I31640));
INVX1 gate10849(.O (I31643), .I (g23737));
INVX1 gate10850(.O (g24323), .I (I31643));
INVX1 gate10851(.O (I31646), .I (g23692));
INVX1 gate10852(.O (g24324), .I (I31646));
INVX1 gate10853(.O (I31649), .I (g23738));
INVX1 gate10854(.O (g24325), .I (I31649));
INVX1 gate10855(.O (I31652), .I (g23784));
INVX1 gate10856(.O (g24326), .I (I31652));
INVX1 gate10857(.O (I31655), .I (g23739));
INVX1 gate10858(.O (g24327), .I (I31655));
INVX1 gate10859(.O (I31658), .I (g23785));
INVX1 gate10860(.O (g24328), .I (I31658));
INVX1 gate10861(.O (I31661), .I (g23828));
INVX1 gate10862(.O (g24329), .I (I31661));
INVX1 gate10863(.O (I31664), .I (g23516));
INVX1 gate10864(.O (g24330), .I (I31664));
INVX1 gate10865(.O (I31667), .I (g23452));
INVX1 gate10866(.O (g24331), .I (I31667));
INVX1 gate10867(.O (I31670), .I (g23463));
INVX1 gate10868(.O (g24332), .I (I31670));
INVX1 gate10869(.O (I31673), .I (g23492));
INVX1 gate10870(.O (g24333), .I (I31673));
INVX1 gate10871(.O (I31676), .I (g23517));
INVX1 gate10872(.O (g24334), .I (I31676));
INVX1 gate10873(.O (I31679), .I (g23453));
INVX1 gate10874(.O (g24335), .I (I31679));
INVX1 gate10875(.O (I31682), .I (g24240));
INVX1 gate10876(.O (g24336), .I (I31682));
INVX1 gate10877(.O (I31685), .I (g23626));
INVX1 gate10878(.O (g24337), .I (I31685));
INVX1 gate10879(.O (I31688), .I (g24035));
INVX1 gate10880(.O (g24338), .I (I31688));
INVX1 gate10881(.O (I31691), .I (g24053));
INVX1 gate10882(.O (g24339), .I (I31691));
INVX1 gate10883(.O (I31694), .I (g24064));
INVX1 gate10884(.O (g24340), .I (I31694));
INVX1 gate10885(.O (I31697), .I (g23791));
INVX1 gate10886(.O (g24341), .I (I31697));
INVX1 gate10887(.O (I31700), .I (g23835));
INVX1 gate10888(.O (g24342), .I (I31700));
INVX1 gate10889(.O (I31703), .I (g23861));
INVX1 gate10890(.O (g24343), .I (I31703));
INVX1 gate10891(.O (I31706), .I (g23836));
INVX1 gate10892(.O (g24344), .I (I31706));
INVX1 gate10893(.O (I31709), .I (g23862));
INVX1 gate10894(.O (g24345), .I (I31709));
INVX1 gate10895(.O (I31712), .I (g23890));
INVX1 gate10896(.O (g24346), .I (I31712));
INVX1 gate10897(.O (I31715), .I (g23566));
INVX1 gate10898(.O (g24347), .I (I31715));
INVX1 gate10899(.O (I31718), .I (g23580));
INVX1 gate10900(.O (g24348), .I (I31718));
INVX1 gate10901(.O (I31721), .I (g23601));
INVX1 gate10902(.O (g24349), .I (I31721));
INVX1 gate10903(.O (I31724), .I (g23581));
INVX1 gate10904(.O (g24350), .I (I31724));
INVX1 gate10905(.O (I31727), .I (g23602));
INVX1 gate10906(.O (g24351), .I (I31727));
INVX1 gate10907(.O (I31730), .I (g23627));
INVX1 gate10908(.O (g24352), .I (I31730));
INVX1 gate10909(.O (I31733), .I (g23603));
INVX1 gate10910(.O (g24353), .I (I31733));
INVX1 gate10911(.O (I31736), .I (g23628));
INVX1 gate10912(.O (g24354), .I (I31736));
INVX1 gate10913(.O (I31739), .I (g23668));
INVX1 gate10914(.O (g24355), .I (I31739));
INVX1 gate10915(.O (I31742), .I (g23629));
INVX1 gate10916(.O (g24356), .I (I31742));
INVX1 gate10917(.O (I31745), .I (g23669));
INVX1 gate10918(.O (g24357), .I (I31745));
INVX1 gate10919(.O (I31748), .I (g23711));
INVX1 gate10920(.O (g24358), .I (I31748));
INVX1 gate10921(.O (I31751), .I (g23670));
INVX1 gate10922(.O (g24359), .I (I31751));
INVX1 gate10923(.O (I31754), .I (g23712));
INVX1 gate10924(.O (g24360), .I (I31754));
INVX1 gate10925(.O (I31757), .I (g23744));
INVX1 gate10926(.O (g24361), .I (I31757));
INVX1 gate10927(.O (I31760), .I (g23713));
INVX1 gate10928(.O (g24362), .I (I31760));
INVX1 gate10929(.O (I31763), .I (g23745));
INVX1 gate10930(.O (g24363), .I (I31763));
INVX1 gate10931(.O (I31766), .I (g23792));
INVX1 gate10932(.O (g24364), .I (I31766));
INVX1 gate10933(.O (I31769), .I (g23746));
INVX1 gate10934(.O (g24365), .I (I31769));
INVX1 gate10935(.O (I31772), .I (g23793));
INVX1 gate10936(.O (g24366), .I (I31772));
INVX1 gate10937(.O (I31775), .I (g23837));
INVX1 gate10938(.O (g24367), .I (I31775));
INVX1 gate10939(.O (I31778), .I (g23794));
INVX1 gate10940(.O (g24368), .I (I31778));
INVX1 gate10941(.O (I31781), .I (g23838));
INVX1 gate10942(.O (g24369), .I (I31781));
INVX1 gate10943(.O (I31784), .I (g23863));
INVX1 gate10944(.O (g24370), .I (I31784));
INVX1 gate10945(.O (I31787), .I (g23531));
INVX1 gate10946(.O (g24371), .I (I31787));
INVX1 gate10947(.O (I31790), .I (g23459));
INVX1 gate10948(.O (g24372), .I (I31790));
INVX1 gate10949(.O (I31793), .I (g23472));
INVX1 gate10950(.O (g24373), .I (I31793));
INVX1 gate10951(.O (I31796), .I (g23508));
INVX1 gate10952(.O (g24374), .I (I31796));
INVX1 gate10953(.O (I31799), .I (g23532));
INVX1 gate10954(.O (g24375), .I (I31799));
INVX1 gate10955(.O (I31802), .I (g23460));
INVX1 gate10956(.O (g24376), .I (I31802));
INVX1 gate10957(.O (I31805), .I (g24248));
INVX1 gate10958(.O (g24377), .I (I31805));
INVX1 gate10959(.O (I31808), .I (g23675));
INVX1 gate10960(.O (g24378), .I (I31808));
INVX1 gate10961(.O (I31811), .I (g24055));
INVX1 gate10962(.O (g24379), .I (I31811));
INVX1 gate10963(.O (I31814), .I (g24066));
INVX1 gate10964(.O (g24380), .I (I31814));
INVX1 gate10965(.O (I31817), .I (g24077));
INVX1 gate10966(.O (g24381), .I (I31817));
INVX1 gate10967(.O (I31820), .I (g23844));
INVX1 gate10968(.O (g24382), .I (I31820));
INVX1 gate10969(.O (I31823), .I (g23870));
INVX1 gate10970(.O (g24383), .I (I31823));
INVX1 gate10971(.O (I31826), .I (g23895));
INVX1 gate10972(.O (g24384), .I (I31826));
INVX1 gate10973(.O (I31829), .I (g23871));
INVX1 gate10974(.O (g24385), .I (I31829));
INVX1 gate10975(.O (I31832), .I (g23896));
INVX1 gate10976(.O (g24386), .I (I31832));
INVX1 gate10977(.O (I31835), .I (g23911));
INVX1 gate10978(.O (g24387), .I (I31835));
INVX1 gate10979(.O (I31838), .I (g23585));
INVX1 gate10980(.O (g24388), .I (I31838));
INVX1 gate10981(.O (I31841), .I (g23607));
INVX1 gate10982(.O (g24389), .I (I31841));
INVX1 gate10983(.O (I31844), .I (g23633));
INVX1 gate10984(.O (g24390), .I (I31844));
INVX1 gate10985(.O (I31847), .I (g23608));
INVX1 gate10986(.O (g24391), .I (I31847));
INVX1 gate10987(.O (I31850), .I (g23634));
INVX1 gate10988(.O (g24392), .I (I31850));
INVX1 gate10989(.O (I31853), .I (g23676));
INVX1 gate10990(.O (g24393), .I (I31853));
INVX1 gate10991(.O (I31856), .I (g23635));
INVX1 gate10992(.O (g24394), .I (I31856));
INVX1 gate10993(.O (I31859), .I (g23677));
INVX1 gate10994(.O (g24395), .I (I31859));
INVX1 gate10995(.O (I31862), .I (g23718));
INVX1 gate10996(.O (g24396), .I (I31862));
INVX1 gate10997(.O (I31865), .I (g23678));
INVX1 gate10998(.O (g24397), .I (I31865));
INVX1 gate10999(.O (I31868), .I (g23719));
INVX1 gate11000(.O (g24398), .I (I31868));
INVX1 gate11001(.O (I31871), .I (g23765));
INVX1 gate11002(.O (g24399), .I (I31871));
INVX1 gate11003(.O (I31874), .I (g23720));
INVX1 gate11004(.O (g24400), .I (I31874));
INVX1 gate11005(.O (I31877), .I (g23766));
INVX1 gate11006(.O (g24401), .I (I31877));
INVX1 gate11007(.O (I31880), .I (g23799));
INVX1 gate11008(.O (g24402), .I (I31880));
INVX1 gate11009(.O (I31883), .I (g23767));
INVX1 gate11010(.O (g24403), .I (I31883));
INVX1 gate11011(.O (I31886), .I (g23800));
INVX1 gate11012(.O (g24404), .I (I31886));
INVX1 gate11013(.O (I31889), .I (g23845));
INVX1 gate11014(.O (g24405), .I (I31889));
INVX1 gate11015(.O (I31892), .I (g23801));
INVX1 gate11016(.O (g24406), .I (I31892));
INVX1 gate11017(.O (I31895), .I (g23846));
INVX1 gate11018(.O (g24407), .I (I31895));
INVX1 gate11019(.O (I31898), .I (g23872));
INVX1 gate11020(.O (g24408), .I (I31898));
INVX1 gate11021(.O (I31901), .I (g23847));
INVX1 gate11022(.O (g24409), .I (I31901));
INVX1 gate11023(.O (I31904), .I (g23873));
INVX1 gate11024(.O (g24410), .I (I31904));
INVX1 gate11025(.O (I31907), .I (g23897));
INVX1 gate11026(.O (g24411), .I (I31907));
INVX1 gate11027(.O (I31910), .I (g23542));
INVX1 gate11028(.O (g24412), .I (I31910));
INVX1 gate11029(.O (I31913), .I (g23468));
INVX1 gate11030(.O (g24413), .I (I31913));
INVX1 gate11031(.O (I31916), .I (g23485));
INVX1 gate11032(.O (g24414), .I (I31916));
INVX1 gate11033(.O (I31919), .I (g23524));
INVX1 gate11034(.O (g24415), .I (I31919));
INVX1 gate11035(.O (I31922), .I (g23543));
INVX1 gate11036(.O (g24416), .I (I31922));
INVX1 gate11037(.O (I31925), .I (g23469));
INVX1 gate11038(.O (g24417), .I (I31925));
INVX1 gate11039(.O (I31928), .I (g24255));
INVX1 gate11040(.O (g24418), .I (I31928));
INVX1 gate11041(.O (I31931), .I (g23725));
INVX1 gate11042(.O (g24419), .I (I31931));
INVX1 gate11043(.O (I31934), .I (g24068));
INVX1 gate11044(.O (g24420), .I (I31934));
INVX1 gate11045(.O (I31937), .I (g24079));
INVX1 gate11046(.O (g24421), .I (I31937));
INVX1 gate11047(.O (I31940), .I (g24088));
INVX1 gate11048(.O (g24422), .I (I31940));
INVX1 gate11049(.O (I31943), .I (g24000));
INVX1 gate11050(.O (g24423), .I (I31943));
INVX1 gate11051(.O (I31946), .I (g23916));
INVX1 gate11052(.O (g24424), .I (I31946));
INVX1 gate11053(.O (I31949), .I (g23943));
INVX1 gate11054(.O (g24425), .I (I31949));
INVX1 gate11055(.O (g24482), .I (g24183));
INVX1 gate11056(.O (I32042), .I (g23399));
INVX1 gate11057(.O (g24518), .I (I32042));
INVX1 gate11058(.O (I32057), .I (g23406));
INVX1 gate11059(.O (g24531), .I (I32057));
INVX1 gate11060(.O (I32067), .I (g24174));
INVX1 gate11061(.O (g24539), .I (I32067));
INVX1 gate11062(.O (I32074), .I (g23413));
INVX1 gate11063(.O (g24544), .I (I32074));
INVX1 gate11064(.O (I32081), .I (g24178));
INVX1 gate11065(.O (g24549), .I (I32081));
INVX1 gate11066(.O (I32085), .I (g24179));
INVX1 gate11067(.O (g24551), .I (I32085));
INVX1 gate11068(.O (I32092), .I (g23418));
INVX1 gate11069(.O (g24556), .I (I32092));
INVX1 gate11070(.O (I32098), .I (g24181));
INVX1 gate11071(.O (g24560), .I (I32098));
INVX1 gate11072(.O (I32102), .I (g24182));
INVX1 gate11073(.O (g24562), .I (I32102));
INVX1 gate11074(.O (I32109), .I (g24206));
INVX1 gate11075(.O (g24567), .I (I32109));
INVX1 gate11076(.O (I32112), .I (g24207));
INVX1 gate11077(.O (g24568), .I (I32112));
INVX1 gate11078(.O (I32116), .I (g24208));
INVX1 gate11079(.O (g24570), .I (I32116));
INVX1 gate11080(.O (I32120), .I (g24209));
INVX1 gate11081(.O (g24572), .I (I32120));
INVX1 gate11082(.O (I32126), .I (g24212));
INVX1 gate11083(.O (g24576), .I (I32126));
INVX1 gate11084(.O (I32129), .I (g24213));
INVX1 gate11085(.O (g24577), .I (I32129));
INVX1 gate11086(.O (I32133), .I (g24214));
INVX1 gate11087(.O (g24579), .I (I32133));
INVX1 gate11088(.O (I32137), .I (g24215));
INVX1 gate11089(.O (g24581), .I (I32137));
INVX1 gate11090(.O (I32140), .I (g24216));
INVX1 gate11091(.O (g24582), .I (I32140));
INVX1 gate11092(.O (I32143), .I (g24218));
INVX1 gate11093(.O (g24583), .I (I32143));
INVX1 gate11094(.O (I32146), .I (g24219));
INVX1 gate11095(.O (g24584), .I (I32146));
INVX1 gate11096(.O (I32150), .I (g24222));
INVX1 gate11097(.O (g24586), .I (I32150));
INVX1 gate11098(.O (I32153), .I (g24223));
INVX1 gate11099(.O (g24587), .I (I32153));
INVX1 gate11100(.O (I32156), .I (g24225));
INVX1 gate11101(.O (g24588), .I (I32156));
INVX1 gate11102(.O (I32159), .I (g24226));
INVX1 gate11103(.O (g24589), .I (I32159));
INVX1 gate11104(.O (I32164), .I (g24228));
INVX1 gate11105(.O (g24592), .I (I32164));
INVX1 gate11106(.O (I32167), .I (g24230));
INVX1 gate11107(.O (g24593), .I (I32167));
INVX1 gate11108(.O (I32170), .I (g24231));
INVX1 gate11109(.O (g24594), .I (I32170));
INVX1 gate11110(.O (I32175), .I (g24235));
INVX1 gate11111(.O (g24597), .I (I32175));
INVX1 gate11112(.O (I32178), .I (g24237));
INVX1 gate11113(.O (g24598), .I (I32178));
INVX1 gate11114(.O (I32181), .I (g24238));
INVX1 gate11115(.O (g24599), .I (I32181));
INVX1 gate11116(.O (I32184), .I (g23497));
INVX1 gate11117(.O (g24600), .I (I32184));
INVX1 gate11118(.O (I32189), .I (g24243));
INVX1 gate11119(.O (g24605), .I (I32189));
INVX1 gate11120(.O (I32193), .I (g23513));
INVX1 gate11121(.O (g24607), .I (I32193));
INVX1 gate11122(.O (I32198), .I (g24250));
INVX1 gate11123(.O (g24612), .I (I32198));
INVX1 gate11124(.O (I32203), .I (g23528));
INVX1 gate11125(.O (g24619), .I (I32203));
INVX1 gate11126(.O (I32210), .I (g23539));
INVX1 gate11127(.O (g24630), .I (I32210));
INVX1 gate11128(.O (g24648), .I (g23470));
INVX1 gate11129(.O (g24668), .I (g23482));
INVX1 gate11130(.O (g24687), .I (g23493));
INVX1 gate11131(.O (g24704), .I (g23509));
INVX1 gate11132(.O (I32248), .I (g23919));
INVX1 gate11133(.O (g24734), .I (I32248));
INVX1 gate11134(.O (I32251), .I (g23919));
INVX1 gate11135(.O (g24735), .I (I32251));
INVX1 gate11136(.O (I32281), .I (g23950));
INVX1 gate11137(.O (g24763), .I (I32281));
INVX1 gate11138(.O (I32320), .I (g23979));
INVX1 gate11139(.O (g24784), .I (I32320));
INVX1 gate11140(.O (I32365), .I (g24009));
INVX1 gate11141(.O (g24805), .I (I32365));
INVX1 gate11142(.O (g24815), .I (g23448));
INVX1 gate11143(.O (I32388), .I (g23385));
INVX1 gate11144(.O (g24816), .I (I32388));
INVX1 gate11145(.O (I32419), .I (g24043));
INVX1 gate11146(.O (g24827), .I (I32419));
INVX1 gate11147(.O (g24834), .I (g23455));
INVX1 gate11148(.O (I32439), .I (g23392));
INVX1 gate11149(.O (g24835), .I (I32439));
INVX1 gate11150(.O (g24850), .I (g23464));
INVX1 gate11151(.O (I32487), .I (g23400));
INVX1 gate11152(.O (g24851), .I (I32487));
INVX1 gate11153(.O (I32506), .I (g23324));
INVX1 gate11154(.O (g24856), .I (I32506));
INVX1 gate11155(.O (g24864), .I (g23473));
INVX1 gate11156(.O (I32535), .I (g23407));
INVX1 gate11157(.O (g24865), .I (I32535));
INVX1 gate11158(.O (I32556), .I (g23329));
INVX1 gate11159(.O (g24872), .I (I32556));
INVX1 gate11160(.O (I32583), .I (g23330));
INVX1 gate11161(.O (g24879), .I (I32583));
INVX1 gate11162(.O (I32604), .I (g23339));
INVX1 gate11163(.O (g24886), .I (I32604));
INVX1 gate11164(.O (g24893), .I (g23486));
INVX1 gate11165(.O (I32642), .I (g23348));
INVX1 gate11166(.O (g24903), .I (I32642));
INVX1 gate11167(.O (g24912), .I (g23495));
INVX1 gate11168(.O (g24916), .I (g23502));
INVX1 gate11169(.O (g24929), .I (g23511));
INVX1 gate11170(.O (g24933), .I (g23518));
INVX1 gate11171(.O (g24939), .I (g23660));
INVX1 gate11172(.O (g24941), .I (g23526));
INVX1 gate11173(.O (g24945), .I (g23533));
INVX1 gate11174(.O (I32704), .I (g23357));
INVX1 gate11175(.O (g24949), .I (I32704));
INVX1 gate11176(.O (g24950), .I (g23710));
INVX1 gate11177(.O (g24952), .I (g23537));
INVX1 gate11178(.O (I32716), .I (g23358));
INVX1 gate11179(.O (g24956), .I (I32716));
INVX1 gate11180(.O (I32719), .I (g23359));
INVX1 gate11181(.O (g24957), .I (I32719));
INVX1 gate11182(.O (g24958), .I (g23478));
INVX1 gate11183(.O (g24962), .I (g23764));
INVX1 gate11184(.O (g24969), .I (g23489));
INVX1 gate11185(.O (g24973), .I (g23819));
INVX1 gate11186(.O (g24982), .I (g23505));
INVX1 gate11187(.O (g24993), .I (g23521));
INVX1 gate11188(.O (g25087), .I (g23731));
INVX1 gate11189(.O (g25094), .I (g23779));
INVX1 gate11190(.O (g25095), .I (g23786));
INVX1 gate11191(.O (I32829), .I (g24059));
INVX1 gate11192(.O (g25103), .I (I32829));
INVX1 gate11193(.O (g25104), .I (g23832));
INVX1 gate11194(.O (g25105), .I (g23839));
INVX1 gate11195(.O (I32835), .I (g24072));
INVX1 gate11196(.O (g25109), .I (I32835));
INVX1 gate11197(.O (g25110), .I (g23867));
INVX1 gate11198(.O (g25111), .I (g23874));
INVX1 gate11199(.O (g25115), .I (g23879));
INVX1 gate11200(.O (g25116), .I (g23882));
INVX1 gate11201(.O (I32844), .I (g23644));
INVX1 gate11202(.O (g25118), .I (I32844));
INVX1 gate11203(.O (I32847), .I (g24083));
INVX1 gate11204(.O (g25119), .I (I32847));
INVX1 gate11205(.O (g25120), .I (g23901));
INVX1 gate11206(.O (I32851), .I (g23694));
INVX1 gate11207(.O (g25121), .I (I32851));
INVX1 gate11208(.O (I32854), .I (g24092));
INVX1 gate11209(.O (g25122), .I (I32854));
INVX1 gate11210(.O (I32857), .I (g23748));
INVX1 gate11211(.O (g25123), .I (I32857));
INVX1 gate11212(.O (I32860), .I (g23803));
INVX1 gate11213(.O (g25124), .I (I32860));
INVX1 gate11214(.O (g25126), .I (g24030));
INVX1 gate11215(.O (I32868), .I (g25118));
INVX1 gate11216(.O (g25130), .I (I32868));
INVX1 gate11217(.O (I32871), .I (g24518));
INVX1 gate11218(.O (g25131), .I (I32871));
INVX1 gate11219(.O (I32874), .I (g24539));
INVX1 gate11220(.O (g25132), .I (I32874));
INVX1 gate11221(.O (I32877), .I (g24567));
INVX1 gate11222(.O (g25133), .I (I32877));
INVX1 gate11223(.O (I32880), .I (g24581));
INVX1 gate11224(.O (g25134), .I (I32880));
INVX1 gate11225(.O (I32883), .I (g24592));
INVX1 gate11226(.O (g25135), .I (I32883));
INVX1 gate11227(.O (I32886), .I (g24549));
INVX1 gate11228(.O (g25136), .I (I32886));
INVX1 gate11229(.O (I32889), .I (g24568));
INVX1 gate11230(.O (g25137), .I (I32889));
INVX1 gate11231(.O (I32892), .I (g24582));
INVX1 gate11232(.O (g25138), .I (I32892));
INVX1 gate11233(.O (I32895), .I (g24816));
INVX1 gate11234(.O (g25139), .I (I32895));
INVX1 gate11235(.O (I32898), .I (g24856));
INVX1 gate11236(.O (g25140), .I (I32898));
INVX1 gate11237(.O (I32901), .I (g25121));
INVX1 gate11238(.O (g25141), .I (I32901));
INVX1 gate11239(.O (I32904), .I (g24531));
INVX1 gate11240(.O (g25142), .I (I32904));
INVX1 gate11241(.O (I32907), .I (g24551));
INVX1 gate11242(.O (g25143), .I (I32907));
INVX1 gate11243(.O (I32910), .I (g24576));
INVX1 gate11244(.O (g25144), .I (I32910));
INVX1 gate11245(.O (I32913), .I (g24586));
INVX1 gate11246(.O (g25145), .I (I32913));
INVX1 gate11247(.O (I32916), .I (g24597));
INVX1 gate11248(.O (g25146), .I (I32916));
INVX1 gate11249(.O (I32919), .I (g24560));
INVX1 gate11250(.O (g25147), .I (I32919));
INVX1 gate11251(.O (I32922), .I (g24577));
INVX1 gate11252(.O (g25148), .I (I32922));
INVX1 gate11253(.O (I32925), .I (g24587));
INVX1 gate11254(.O (g25149), .I (I32925));
INVX1 gate11255(.O (I32928), .I (g24835));
INVX1 gate11256(.O (g25150), .I (I32928));
INVX1 gate11257(.O (I32931), .I (g24872));
INVX1 gate11258(.O (g25151), .I (I32931));
INVX1 gate11259(.O (I32934), .I (g25123));
INVX1 gate11260(.O (g25152), .I (I32934));
INVX1 gate11261(.O (I32937), .I (g24544));
INVX1 gate11262(.O (g25153), .I (I32937));
INVX1 gate11263(.O (I32940), .I (g24562));
INVX1 gate11264(.O (g25154), .I (I32940));
INVX1 gate11265(.O (I32943), .I (g24583));
INVX1 gate11266(.O (g25155), .I (I32943));
INVX1 gate11267(.O (I32946), .I (g24593));
INVX1 gate11268(.O (g25156), .I (I32946));
INVX1 gate11269(.O (I32949), .I (g24605));
INVX1 gate11270(.O (g25157), .I (I32949));
INVX1 gate11271(.O (I32952), .I (g24570));
INVX1 gate11272(.O (g25158), .I (I32952));
INVX1 gate11273(.O (I32955), .I (g24584));
INVX1 gate11274(.O (g25159), .I (I32955));
INVX1 gate11275(.O (I32958), .I (g24594));
INVX1 gate11276(.O (g25160), .I (I32958));
INVX1 gate11277(.O (I32961), .I (g24851));
INVX1 gate11278(.O (g25161), .I (I32961));
INVX1 gate11279(.O (I32964), .I (g24886));
INVX1 gate11280(.O (g25162), .I (I32964));
INVX1 gate11281(.O (I32967), .I (g25124));
INVX1 gate11282(.O (g25163), .I (I32967));
INVX1 gate11283(.O (I32970), .I (g24556));
INVX1 gate11284(.O (g25164), .I (I32970));
INVX1 gate11285(.O (I32973), .I (g24572));
INVX1 gate11286(.O (g25165), .I (I32973));
INVX1 gate11287(.O (I32976), .I (g24588));
INVX1 gate11288(.O (g25166), .I (I32976));
INVX1 gate11289(.O (I32979), .I (g24598));
INVX1 gate11290(.O (g25167), .I (I32979));
INVX1 gate11291(.O (I32982), .I (g24612));
INVX1 gate11292(.O (g25168), .I (I32982));
INVX1 gate11293(.O (I32985), .I (g24579));
INVX1 gate11294(.O (g25169), .I (I32985));
INVX1 gate11295(.O (I32988), .I (g24589));
INVX1 gate11296(.O (g25170), .I (I32988));
INVX1 gate11297(.O (I32991), .I (g24599));
INVX1 gate11298(.O (g25171), .I (I32991));
INVX1 gate11299(.O (I32994), .I (g24865));
INVX1 gate11300(.O (g25172), .I (I32994));
INVX1 gate11301(.O (I32997), .I (g24903));
INVX1 gate11302(.O (g25173), .I (I32997));
INVX1 gate11303(.O (I33000), .I (g24949));
INVX1 gate11304(.O (g25174), .I (I33000));
INVX1 gate11305(.O (I33003), .I (g24956));
INVX1 gate11306(.O (g25175), .I (I33003));
INVX1 gate11307(.O (I33006), .I (g24957));
INVX1 gate11308(.O (g25176), .I (I33006));
INVX1 gate11309(.O (I33009), .I (g24879));
INVX1 gate11310(.O (g25177), .I (I33009));
INVX1 gate11311(.O (I33013), .I (g25119));
INVX1 gate11312(.O (g25179), .I (I33013));
INVX1 gate11313(.O (I33016), .I (g25122));
INVX1 gate11314(.O (g25180), .I (I33016));
INVX1 gate11315(.O (g25274), .I (g24912));
INVX1 gate11316(.O (g25283), .I (g24929));
INVX1 gate11317(.O (g25291), .I (g24941));
INVX1 gate11318(.O (I33128), .I (g24975));
INVX1 gate11319(.O (g25296), .I (I33128));
INVX1 gate11320(.O (g25301), .I (g24952));
INVX1 gate11321(.O (g25305), .I (g24880));
INVX1 gate11322(.O (I33136), .I (g24986));
INVX1 gate11323(.O (g25306), .I (I33136));
INVX1 gate11324(.O (g25313), .I (g24868));
INVX1 gate11325(.O (g25314), .I (g24897));
INVX1 gate11326(.O (I33145), .I (g24997));
INVX1 gate11327(.O (g25315), .I (I33145));
INVX1 gate11328(.O (g25319), .I (g24857));
INVX1 gate11329(.O (g25322), .I (g24883));
INVX1 gate11330(.O (g25323), .I (g24920));
INVX1 gate11331(.O (I33154), .I (g25005));
INVX1 gate11332(.O (g25324), .I (I33154));
INVX1 gate11333(.O (I33157), .I (g25027));
INVX1 gate11334(.O (g25327), .I (I33157));
INVX1 gate11335(.O (g25329), .I (g24844));
INVX1 gate11336(.O (g25330), .I (g24873));
INVX1 gate11337(.O (g25332), .I (g24900));
INVX1 gate11338(.O (g25333), .I (g24937));
INVX1 gate11339(.O (g25335), .I (g24832));
INVX1 gate11340(.O (I33168), .I (g25042));
INVX1 gate11341(.O (g25336), .I (I33168));
INVX1 gate11342(.O (g25338), .I (g24860));
INVX1 gate11343(.O (g25339), .I (g24887));
INVX1 gate11344(.O (g25341), .I (g24923));
INVX1 gate11345(.O (g25347), .I (g24817));
INVX1 gate11346(.O (g25349), .I (g24848));
INVX1 gate11347(.O (I33182), .I (g25056));
INVX1 gate11348(.O (g25350), .I (I33182));
INVX1 gate11349(.O (g25352), .I (g24875));
INVX1 gate11350(.O (g25353), .I (g24904));
INVX1 gate11351(.O (I33188), .I (g24814));
INVX1 gate11352(.O (g25354), .I (I33188));
INVX1 gate11353(.O (g25355), .I (g24797));
INVX1 gate11354(.O (g25361), .I (g24837));
INVX1 gate11355(.O (g25363), .I (g24862));
INVX1 gate11356(.O (I33198), .I (g25067));
INVX1 gate11357(.O (g25364), .I (I33198));
INVX1 gate11358(.O (g25366), .I (g24889));
INVX1 gate11359(.O (g25367), .I (g24676));
INVX1 gate11360(.O (g25368), .I (g24778));
INVX1 gate11361(.O (I33205), .I (g24833));
INVX1 gate11362(.O (g25369), .I (I33205));
INVX1 gate11363(.O (g25370), .I (g24820));
INVX1 gate11364(.O (g25376), .I (g24852));
INVX1 gate11365(.O (g25378), .I (g24877));
INVX1 gate11366(.O (g25379), .I (g24893));
INVX1 gate11367(.O (g25383), .I (g24766));
INVX1 gate11368(.O (g25384), .I (g24695));
INVX1 gate11369(.O (g25385), .I (g24801));
INVX1 gate11370(.O (I33219), .I (g24849));
INVX1 gate11371(.O (g25386), .I (I33219));
INVX1 gate11372(.O (g25387), .I (g24839));
INVX1 gate11373(.O (g25393), .I (g24866));
INVX1 gate11374(.O (g25394), .I (g24753));
INVX1 gate11375(.O (g25395), .I (g24916));
INVX1 gate11376(.O (g25399), .I (g24787));
INVX1 gate11377(.O (g25400), .I (g24712));
INVX1 gate11378(.O (g25401), .I (g24823));
INVX1 gate11379(.O (I33232), .I (g24863));
INVX1 gate11380(.O (g25402), .I (I33232));
INVX1 gate11381(.O (g25403), .I (g24854));
INVX1 gate11382(.O (g25404), .I (g24771));
INVX1 gate11383(.O (g25405), .I (g24933));
INVX1 gate11384(.O (g25409), .I (g24808));
INVX1 gate11385(.O (g25410), .I (g24723));
INVX1 gate11386(.O (g25411), .I (g24842));
INVX1 gate11387(.O (g25412), .I (g24791));
INVX1 gate11388(.O (g25413), .I (g24945));
INVX1 gate11389(.O (g25417), .I (g24830));
INVX1 gate11390(.O (g25419), .I (g24812));
INVX1 gate11391(.O (I33246), .I (g24890));
INVX1 gate11392(.O (g25420), .I (I33246));
INVX1 gate11393(.O (I33249), .I (g24890));
INVX1 gate11394(.O (g25421), .I (I33249));
INVX1 gate11395(.O (g25422), .I (g24958));
INVX1 gate11396(.O (g25430), .I (g24616));
INVX1 gate11397(.O (g25431), .I (g24969));
INVX1 gate11398(.O (I33257), .I (g24909));
INVX1 gate11399(.O (g25435), .I (I33257));
INVX1 gate11400(.O (I33260), .I (g24909));
INVX1 gate11401(.O (g25436), .I (I33260));
INVX1 gate11402(.O (g25437), .I (g24627));
INVX1 gate11403(.O (g25438), .I (g24982));
INVX1 gate11404(.O (I33265), .I (g24925));
INVX1 gate11405(.O (g25442), .I (I33265));
INVX1 gate11406(.O (I33268), .I (g24925));
INVX1 gate11407(.O (g25443), .I (I33268));
INVX1 gate11408(.O (g25444), .I (g24641));
INVX1 gate11409(.O (g25445), .I (g24993));
INVX1 gate11410(.O (g25449), .I (g24660));
INVX1 gate11411(.O (I33278), .I (g25088));
INVX1 gate11412(.O (g25454), .I (I33278));
INVX1 gate11413(.O (I33282), .I (g25096));
INVX1 gate11414(.O (g25458), .I (I33282));
INVX1 gate11415(.O (I33286), .I (g24426));
INVX1 gate11416(.O (g25462), .I (I33286));
INVX1 gate11417(.O (I33289), .I (g25106));
INVX1 gate11418(.O (g25463), .I (I33289));
INVX1 gate11419(.O (I33293), .I (g25008));
INVX1 gate11420(.O (g25467), .I (I33293));
INVX1 gate11421(.O (I33297), .I (g24430));
INVX1 gate11422(.O (g25471), .I (I33297));
INVX1 gate11423(.O (I33300), .I (g25112));
INVX1 gate11424(.O (g25472), .I (I33300));
INVX1 gate11425(.O (I33304), .I (g25004));
INVX1 gate11426(.O (g25476), .I (I33304));
INVX1 gate11427(.O (I33307), .I (g25011));
INVX1 gate11428(.O (g25479), .I (I33307));
INVX1 gate11429(.O (I33312), .I (g25014));
INVX1 gate11430(.O (g25484), .I (I33312));
INVX1 gate11431(.O (I33316), .I (g24434));
INVX1 gate11432(.O (g25488), .I (I33316));
INVX1 gate11433(.O (I33321), .I (g24442));
INVX1 gate11434(.O (g25493), .I (I33321));
INVX1 gate11435(.O (I33324), .I (g25009));
INVX1 gate11436(.O (g25496), .I (I33324));
INVX1 gate11437(.O (I33327), .I (g25017));
INVX1 gate11438(.O (g25499), .I (I33327));
INVX1 gate11439(.O (I33330), .I (g25019));
INVX1 gate11440(.O (g25502), .I (I33330));
INVX1 gate11441(.O (I33335), .I (g25010));
INVX1 gate11442(.O (g25507), .I (I33335));
INVX1 gate11443(.O (I33338), .I (g25021));
INVX1 gate11444(.O (g25510), .I (I33338));
INVX1 gate11445(.O (I33343), .I (g25024));
INVX1 gate11446(.O (g25515), .I (I33343));
INVX1 gate11447(.O (I33347), .I (g24438));
INVX1 gate11448(.O (g25519), .I (I33347));
INVX1 gate11449(.O (I33352), .I (g24443));
INVX1 gate11450(.O (g25524), .I (I33352));
INVX1 gate11451(.O (I33355), .I (g25012));
INVX1 gate11452(.O (g25527), .I (I33355));
INVX1 gate11453(.O (I33358), .I (g25028));
INVX1 gate11454(.O (g25530), .I (I33358));
INVX1 gate11455(.O (I33361), .I (g25013));
INVX1 gate11456(.O (g25533), .I (I33361));
INVX1 gate11457(.O (I33364), .I (g25029));
INVX1 gate11458(.O (g25536), .I (I33364));
INVX1 gate11459(.O (I33368), .I (g24444));
INVX1 gate11460(.O (g25540), .I (I33368));
INVX1 gate11461(.O (I33371), .I (g25015));
INVX1 gate11462(.O (g25543), .I (I33371));
INVX1 gate11463(.O (I33374), .I (g25031));
INVX1 gate11464(.O (g25546), .I (I33374));
INVX1 gate11465(.O (I33377), .I (g25033));
INVX1 gate11466(.O (g25549), .I (I33377));
INVX1 gate11467(.O (I33382), .I (g25016));
INVX1 gate11468(.O (g25554), .I (I33382));
INVX1 gate11469(.O (I33385), .I (g25035));
INVX1 gate11470(.O (g25557), .I (I33385));
INVX1 gate11471(.O (I33390), .I (g25038));
INVX1 gate11472(.O (g25562), .I (I33390));
INVX1 gate11473(.O (I33396), .I (g24447));
INVX1 gate11474(.O (g25573), .I (I33396));
INVX1 gate11475(.O (I33399), .I (g25018));
INVX1 gate11476(.O (g25576), .I (I33399));
INVX1 gate11477(.O (I33402), .I (g24448));
INVX1 gate11478(.O (g25579), .I (I33402));
INVX1 gate11479(.O (I33405), .I (g25020));
INVX1 gate11480(.O (g25582), .I (I33405));
INVX1 gate11481(.O (I33408), .I (g25040));
INVX1 gate11482(.O (g25585), .I (I33408));
INVX1 gate11483(.O (I33411), .I (g24491));
INVX1 gate11484(.O (g25588), .I (I33411));
INVX1 gate11485(.O (I33415), .I (g24449));
INVX1 gate11486(.O (g25590), .I (I33415));
INVX1 gate11487(.O (I33418), .I (g25022));
INVX1 gate11488(.O (g25593), .I (I33418));
INVX1 gate11489(.O (I33421), .I (g25043));
INVX1 gate11490(.O (g25596), .I (I33421));
INVX1 gate11491(.O (I33424), .I (g25023));
INVX1 gate11492(.O (g25599), .I (I33424));
INVX1 gate11493(.O (I33427), .I (g25044));
INVX1 gate11494(.O (g25602), .I (I33427));
INVX1 gate11495(.O (I33431), .I (g24450));
INVX1 gate11496(.O (g25606), .I (I33431));
INVX1 gate11497(.O (I33434), .I (g25025));
INVX1 gate11498(.O (g25609), .I (I33434));
INVX1 gate11499(.O (I33437), .I (g25046));
INVX1 gate11500(.O (g25612), .I (I33437));
INVX1 gate11501(.O (I33440), .I (g25048));
INVX1 gate11502(.O (g25615), .I (I33440));
INVX1 gate11503(.O (I33445), .I (g25026));
INVX1 gate11504(.O (g25620), .I (I33445));
INVX1 gate11505(.O (I33448), .I (g25050));
INVX1 gate11506(.O (g25623), .I (I33448));
INVX1 gate11507(.O (g25630), .I (g24478));
INVX1 gate11508(.O (I33457), .I (g24451));
INVX1 gate11509(.O (g25634), .I (I33457));
INVX1 gate11510(.O (I33460), .I (g24452));
INVX1 gate11511(.O (g25637), .I (I33460));
INVX1 gate11512(.O (I33463), .I (g25030));
INVX1 gate11513(.O (g25640), .I (I33463));
INVX1 gate11514(.O (I33466), .I (g25053));
INVX1 gate11515(.O (g25643), .I (I33466));
INVX1 gate11516(.O (I33469), .I (g24498));
INVX1 gate11517(.O (g25646), .I (I33469));
INVX1 gate11518(.O (I33472), .I (g24499));
INVX1 gate11519(.O (g25647), .I (I33472));
INVX1 gate11520(.O (I33476), .I (g24453));
INVX1 gate11521(.O (g25652), .I (I33476));
INVX1 gate11522(.O (I33479), .I (g25032));
INVX1 gate11523(.O (g25655), .I (I33479));
INVX1 gate11524(.O (I33482), .I (g24454));
INVX1 gate11525(.O (g25658), .I (I33482));
INVX1 gate11526(.O (I33485), .I (g25034));
INVX1 gate11527(.O (g25661), .I (I33485));
INVX1 gate11528(.O (I33488), .I (g25054));
INVX1 gate11529(.O (g25664), .I (I33488));
INVX1 gate11530(.O (I33491), .I (g24501));
INVX1 gate11531(.O (g25667), .I (I33491));
INVX1 gate11532(.O (I33495), .I (g24455));
INVX1 gate11533(.O (g25669), .I (I33495));
INVX1 gate11534(.O (I33498), .I (g25036));
INVX1 gate11535(.O (g25672), .I (I33498));
INVX1 gate11536(.O (I33501), .I (g25057));
INVX1 gate11537(.O (g25675), .I (I33501));
INVX1 gate11538(.O (I33504), .I (g25037));
INVX1 gate11539(.O (g25678), .I (I33504));
INVX1 gate11540(.O (I33507), .I (g25058));
INVX1 gate11541(.O (g25681), .I (I33507));
INVX1 gate11542(.O (I33511), .I (g24456));
INVX1 gate11543(.O (g25685), .I (I33511));
INVX1 gate11544(.O (I33514), .I (g25039));
INVX1 gate11545(.O (g25688), .I (I33514));
INVX1 gate11546(.O (I33517), .I (g25060));
INVX1 gate11547(.O (g25691), .I (I33517));
INVX1 gate11548(.O (I33520), .I (g25062));
INVX1 gate11549(.O (g25694), .I (I33520));
INVX1 gate11550(.O (g25698), .I (g24600));
INVX1 gate11551(.O (I33526), .I (g24457));
INVX1 gate11552(.O (g25700), .I (I33526));
INVX1 gate11553(.O (I33529), .I (g25041));
INVX1 gate11554(.O (g25703), .I (I33529));
INVX1 gate11555(.O (I33532), .I (g24507));
INVX1 gate11556(.O (g25706), .I (I33532));
INVX1 gate11557(.O (I33535), .I (g24508));
INVX1 gate11558(.O (g25707), .I (I33535));
INVX1 gate11559(.O (I33539), .I (g24458));
INVX1 gate11560(.O (g25711), .I (I33539));
INVX1 gate11561(.O (I33542), .I (g24459));
INVX1 gate11562(.O (g25714), .I (I33542));
INVX1 gate11563(.O (I33545), .I (g25045));
INVX1 gate11564(.O (g25717), .I (I33545));
INVX1 gate11565(.O (I33548), .I (g25064));
INVX1 gate11566(.O (g25720), .I (I33548));
INVX1 gate11567(.O (I33551), .I (g24510));
INVX1 gate11568(.O (g25723), .I (I33551));
INVX1 gate11569(.O (I33554), .I (g24511));
INVX1 gate11570(.O (g25724), .I (I33554));
INVX1 gate11571(.O (I33558), .I (g24460));
INVX1 gate11572(.O (g25729), .I (I33558));
INVX1 gate11573(.O (I33561), .I (g25047));
INVX1 gate11574(.O (g25732), .I (I33561));
INVX1 gate11575(.O (I33564), .I (g24461));
INVX1 gate11576(.O (g25735), .I (I33564));
INVX1 gate11577(.O (I33567), .I (g25049));
INVX1 gate11578(.O (g25738), .I (I33567));
INVX1 gate11579(.O (I33570), .I (g25065));
INVX1 gate11580(.O (g25741), .I (I33570));
INVX1 gate11581(.O (I33573), .I (g24513));
INVX1 gate11582(.O (g25744), .I (I33573));
INVX1 gate11583(.O (I33577), .I (g24462));
INVX1 gate11584(.O (g25746), .I (I33577));
INVX1 gate11585(.O (I33580), .I (g25051));
INVX1 gate11586(.O (g25749), .I (I33580));
INVX1 gate11587(.O (I33583), .I (g25068));
INVX1 gate11588(.O (g25752), .I (I33583));
INVX1 gate11589(.O (I33586), .I (g25052));
INVX1 gate11590(.O (g25755), .I (I33586));
INVX1 gate11591(.O (I33589), .I (g25069));
INVX1 gate11592(.O (g25758), .I (I33589));
INVX1 gate11593(.O (I33593), .I (g24445));
INVX1 gate11594(.O (g25762), .I (I33593));
INVX1 gate11595(.O (I33596), .I (g24446));
INVX1 gate11596(.O (g25763), .I (I33596));
INVX1 gate11597(.O (I33600), .I (g24463));
INVX1 gate11598(.O (g25767), .I (I33600));
INVX1 gate11599(.O (I33603), .I (g24519));
INVX1 gate11600(.O (g25770), .I (I33603));
INVX1 gate11601(.O (g25771), .I (g24607));
INVX1 gate11602(.O (I33608), .I (g24464));
INVX1 gate11603(.O (g25773), .I (I33608));
INVX1 gate11604(.O (I33611), .I (g25055));
INVX1 gate11605(.O (g25776), .I (I33611));
INVX1 gate11606(.O (I33614), .I (g24521));
INVX1 gate11607(.O (g25779), .I (I33614));
INVX1 gate11608(.O (I33617), .I (g24522));
INVX1 gate11609(.O (g25780), .I (I33617));
INVX1 gate11610(.O (I33621), .I (g24465));
INVX1 gate11611(.O (g25784), .I (I33621));
INVX1 gate11612(.O (I33624), .I (g24466));
INVX1 gate11613(.O (g25787), .I (I33624));
INVX1 gate11614(.O (I33627), .I (g25059));
INVX1 gate11615(.O (g25790), .I (I33627));
INVX1 gate11616(.O (I33630), .I (g25071));
INVX1 gate11617(.O (g25793), .I (I33630));
INVX1 gate11618(.O (I33633), .I (g24524));
INVX1 gate11619(.O (g25796), .I (I33633));
INVX1 gate11620(.O (I33636), .I (g24525));
INVX1 gate11621(.O (g25797), .I (I33636));
INVX1 gate11622(.O (I33640), .I (g24467));
INVX1 gate11623(.O (g25802), .I (I33640));
INVX1 gate11624(.O (I33643), .I (g25061));
INVX1 gate11625(.O (g25805), .I (I33643));
INVX1 gate11626(.O (I33646), .I (g24468));
INVX1 gate11627(.O (g25808), .I (I33646));
INVX1 gate11628(.O (I33649), .I (g25063));
INVX1 gate11629(.O (g25811), .I (I33649));
INVX1 gate11630(.O (I33652), .I (g25072));
INVX1 gate11631(.O (g25814), .I (I33652));
INVX1 gate11632(.O (I33655), .I (g24527));
INVX1 gate11633(.O (g25817), .I (I33655));
INVX1 gate11634(.O (I33659), .I (g24469));
INVX1 gate11635(.O (g25821), .I (I33659));
INVX1 gate11636(.O (I33662), .I (g24532));
INVX1 gate11637(.O (g25824), .I (I33662));
INVX1 gate11638(.O (g25825), .I (g24619));
INVX1 gate11639(.O (I33667), .I (g24470));
INVX1 gate11640(.O (g25827), .I (I33667));
INVX1 gate11641(.O (I33670), .I (g25066));
INVX1 gate11642(.O (g25830), .I (I33670));
INVX1 gate11643(.O (I33673), .I (g24534));
INVX1 gate11644(.O (g25833), .I (I33673));
INVX1 gate11645(.O (I33676), .I (g24535));
INVX1 gate11646(.O (g25834), .I (I33676));
INVX1 gate11647(.O (I33680), .I (g24471));
INVX1 gate11648(.O (g25838), .I (I33680));
INVX1 gate11649(.O (I33683), .I (g24472));
INVX1 gate11650(.O (g25841), .I (I33683));
INVX1 gate11651(.O (I33686), .I (g25070));
INVX1 gate11652(.O (g25844), .I (I33686));
INVX1 gate11653(.O (I33689), .I (g25074));
INVX1 gate11654(.O (g25847), .I (I33689));
INVX1 gate11655(.O (I33692), .I (g24537));
INVX1 gate11656(.O (g25850), .I (I33692));
INVX1 gate11657(.O (I33695), .I (g24538));
INVX1 gate11658(.O (g25851), .I (I33695));
INVX1 gate11659(.O (I33700), .I (g24474));
INVX1 gate11660(.O (g25856), .I (I33700));
INVX1 gate11661(.O (I33703), .I (g24545));
INVX1 gate11662(.O (g25859), .I (I33703));
INVX1 gate11663(.O (g25860), .I (g24630));
INVX1 gate11664(.O (I33708), .I (g24475));
INVX1 gate11665(.O (g25862), .I (I33708));
INVX1 gate11666(.O (I33711), .I (g25073));
INVX1 gate11667(.O (g25865), .I (I33711));
INVX1 gate11668(.O (I33714), .I (g24547));
INVX1 gate11669(.O (g25868), .I (I33714));
INVX1 gate11670(.O (I33717), .I (g24548));
INVX1 gate11671(.O (g25869), .I (I33717));
INVX1 gate11672(.O (I33723), .I (g24477));
INVX1 gate11673(.O (g25877), .I (I33723));
INVX1 gate11674(.O (I33726), .I (g24557));
INVX1 gate11675(.O (g25880), .I (I33726));
INVX1 gate11676(.O (I33732), .I (g24473));
INVX1 gate11677(.O (g25886), .I (I33732));
INVX1 gate11678(.O (I33737), .I (g24476));
INVX1 gate11679(.O (g25891), .I (I33737));
INVX1 gate11680(.O (g25895), .I (g24939));
INVX1 gate11681(.O (g25899), .I (g24928));
INVX1 gate11682(.O (g25903), .I (g24950));
INVX1 gate11683(.O (g25907), .I (g24940));
INVX1 gate11684(.O (g25911), .I (g24962));
INVX1 gate11685(.O (g25915), .I (g24951));
INVX1 gate11686(.O (g25919), .I (g24973));
INVX1 gate11687(.O (g25923), .I (g24963));
INVX1 gate11688(.O (g25937), .I (g24763));
INVX1 gate11689(.O (g25939), .I (g24784));
INVX1 gate11690(.O (g25942), .I (g24805));
INVX1 gate11691(.O (g25945), .I (g24827));
INVX1 gate11692(.O (g25952), .I (g24735));
INVX1 gate11693(.O (I33790), .I (g25103));
INVX1 gate11694(.O (g25976), .I (I33790));
INVX1 gate11695(.O (I33798), .I (g25109));
INVX1 gate11696(.O (g25982), .I (I33798));
INVX1 gate11697(.O (I33801), .I (g25327));
INVX1 gate11698(.O (g25983), .I (I33801));
INVX1 gate11699(.O (I33804), .I (g25976));
INVX1 gate11700(.O (g25984), .I (I33804));
INVX1 gate11701(.O (I33807), .I (g25588));
INVX1 gate11702(.O (g25985), .I (I33807));
INVX1 gate11703(.O (I33810), .I (g25646));
INVX1 gate11704(.O (g25986), .I (I33810));
INVX1 gate11705(.O (I33813), .I (g25706));
INVX1 gate11706(.O (g25987), .I (I33813));
INVX1 gate11707(.O (I33816), .I (g25647));
INVX1 gate11708(.O (g25988), .I (I33816));
INVX1 gate11709(.O (I33819), .I (g25707));
INVX1 gate11710(.O (g25989), .I (I33819));
INVX1 gate11711(.O (I33822), .I (g25770));
INVX1 gate11712(.O (g25990), .I (I33822));
INVX1 gate11713(.O (I33825), .I (g25462));
INVX1 gate11714(.O (g25991), .I (I33825));
INVX1 gate11715(.O (I33828), .I (g25336));
INVX1 gate11716(.O (g25992), .I (I33828));
INVX1 gate11717(.O (I33831), .I (g25982));
INVX1 gate11718(.O (g25993), .I (I33831));
INVX1 gate11719(.O (I33834), .I (g25667));
INVX1 gate11720(.O (g25994), .I (I33834));
INVX1 gate11721(.O (I33837), .I (g25723));
INVX1 gate11722(.O (g25995), .I (I33837));
INVX1 gate11723(.O (I33840), .I (g25779));
INVX1 gate11724(.O (g25996), .I (I33840));
INVX1 gate11725(.O (I33843), .I (g25724));
INVX1 gate11726(.O (g25997), .I (I33843));
INVX1 gate11727(.O (I33846), .I (g25780));
INVX1 gate11728(.O (g25998), .I (I33846));
INVX1 gate11729(.O (I33849), .I (g25824));
INVX1 gate11730(.O (g25999), .I (I33849));
INVX1 gate11731(.O (I33852), .I (g25471));
INVX1 gate11732(.O (g26000), .I (I33852));
INVX1 gate11733(.O (I33855), .I (g25350));
INVX1 gate11734(.O (g26001), .I (I33855));
INVX1 gate11735(.O (I33858), .I (g25179));
INVX1 gate11736(.O (g26002), .I (I33858));
INVX1 gate11737(.O (I33861), .I (g25744));
INVX1 gate11738(.O (g26003), .I (I33861));
INVX1 gate11739(.O (I33864), .I (g25796));
INVX1 gate11740(.O (g26004), .I (I33864));
INVX1 gate11741(.O (I33867), .I (g25833));
INVX1 gate11742(.O (g26005), .I (I33867));
INVX1 gate11743(.O (I33870), .I (g25797));
INVX1 gate11744(.O (g26006), .I (I33870));
INVX1 gate11745(.O (I33873), .I (g25834));
INVX1 gate11746(.O (g26007), .I (I33873));
INVX1 gate11747(.O (I33876), .I (g25859));
INVX1 gate11748(.O (g26008), .I (I33876));
INVX1 gate11749(.O (I33879), .I (g25488));
INVX1 gate11750(.O (g26009), .I (I33879));
INVX1 gate11751(.O (I33882), .I (g25364));
INVX1 gate11752(.O (g26010), .I (I33882));
INVX1 gate11753(.O (I33885), .I (g25180));
INVX1 gate11754(.O (g26011), .I (I33885));
INVX1 gate11755(.O (I33888), .I (g25817));
INVX1 gate11756(.O (g26012), .I (I33888));
INVX1 gate11757(.O (I33891), .I (g25850));
INVX1 gate11758(.O (g26013), .I (I33891));
INVX1 gate11759(.O (I33894), .I (g25868));
INVX1 gate11760(.O (g26014), .I (I33894));
INVX1 gate11761(.O (I33897), .I (g25851));
INVX1 gate11762(.O (g26015), .I (I33897));
INVX1 gate11763(.O (I33900), .I (g25869));
INVX1 gate11764(.O (g26016), .I (I33900));
INVX1 gate11765(.O (I33903), .I (g25880));
INVX1 gate11766(.O (g26017), .I (I33903));
INVX1 gate11767(.O (I33906), .I (g25519));
INVX1 gate11768(.O (g26018), .I (I33906));
INVX1 gate11769(.O (I33909), .I (g25886));
INVX1 gate11770(.O (g26019), .I (I33909));
INVX1 gate11771(.O (I33912), .I (g25891));
INVX1 gate11772(.O (g26020), .I (I33912));
INVX1 gate11773(.O (I33915), .I (g25762));
INVX1 gate11774(.O (g26021), .I (I33915));
INVX1 gate11775(.O (I33918), .I (g25763));
INVX1 gate11776(.O (g26022), .I (I33918));
INVX1 gate11777(.O (I33954), .I (g25343));
INVX1 gate11778(.O (g26056), .I (I33954));
INVX1 gate11779(.O (I33961), .I (g25357));
INVX1 gate11780(.O (g26063), .I (I33961));
INVX1 gate11781(.O (I33968), .I (g25372));
INVX1 gate11782(.O (g26070), .I (I33968));
INVX1 gate11783(.O (I33974), .I (g25389));
INVX1 gate11784(.O (g26076), .I (I33974));
INVX1 gate11785(.O (I33984), .I (g25932));
INVX1 gate11786(.O (g26086), .I (I33984));
INVX1 gate11787(.O (I33990), .I (g25870));
INVX1 gate11788(.O (g26092), .I (I33990));
INVX1 gate11789(.O (I33995), .I (g25935));
INVX1 gate11790(.O (g26102), .I (I33995));
INVX1 gate11791(.O (I33999), .I (g25490));
INVX1 gate11792(.O (g26104), .I (I33999));
INVX1 gate11793(.O (I34002), .I (g25490));
INVX1 gate11794(.O (g26105), .I (I34002));
INVX1 gate11795(.O (I34009), .I (g25882));
INVX1 gate11796(.O (g26114), .I (I34009));
INVX1 gate11797(.O (I34012), .I (g25938));
INVX1 gate11798(.O (g26118), .I (I34012));
INVX1 gate11799(.O (I34017), .I (g25887));
INVX1 gate11800(.O (g26121), .I (I34017));
INVX1 gate11801(.O (I34020), .I (g25940));
INVX1 gate11802(.O (g26125), .I (I34020));
INVX1 gate11803(.O (I34026), .I (g25892));
INVX1 gate11804(.O (g26131), .I (I34026));
INVX1 gate11805(.O (I34029), .I (g25520));
INVX1 gate11806(.O (g26135), .I (I34029));
INVX1 gate11807(.O (I34032), .I (g25520));
INVX1 gate11808(.O (g26136), .I (I34032));
INVX1 gate11809(.O (I34041), .I (g25566));
INVX1 gate11810(.O (g26149), .I (I34041));
INVX1 gate11811(.O (I34044), .I (g25566));
INVX1 gate11812(.O (g26150), .I (I34044));
INVX1 gate11813(.O (I34051), .I (g25204));
INVX1 gate11814(.O (g26159), .I (I34051));
INVX1 gate11815(.O (I34056), .I (g25206));
INVX1 gate11816(.O (g26164), .I (I34056));
INVX1 gate11817(.O (I34059), .I (g25207));
INVX1 gate11818(.O (g26165), .I (I34059));
INVX1 gate11819(.O (I34063), .I (g25209));
INVX1 gate11820(.O (g26167), .I (I34063));
INVX1 gate11821(.O (I34068), .I (g25211));
INVX1 gate11822(.O (g26172), .I (I34068));
INVX1 gate11823(.O (I34071), .I (g25212));
INVX1 gate11824(.O (g26173), .I (I34071));
INVX1 gate11825(.O (I34074), .I (g25213));
INVX1 gate11826(.O (g26174), .I (I34074));
INVX1 gate11827(.O (I34077), .I (g25954));
INVX1 gate11828(.O (g26175), .I (I34077));
INVX1 gate11829(.O (I34080), .I (g25539));
INVX1 gate11830(.O (g26178), .I (I34080));
INVX1 gate11831(.O (I34083), .I (g25214));
INVX1 gate11832(.O (g26181), .I (I34083));
INVX1 gate11833(.O (I34086), .I (g25215));
INVX1 gate11834(.O (g26182), .I (I34086));
INVX1 gate11835(.O (I34091), .I (g25217));
INVX1 gate11836(.O (g26187), .I (I34091));
INVX1 gate11837(.O (g26189), .I (g25952));
INVX1 gate11838(.O (I34096), .I (g25218));
INVX1 gate11839(.O (g26190), .I (I34096));
INVX1 gate11840(.O (I34099), .I (g25219));
INVX1 gate11841(.O (g26191), .I (I34099));
INVX1 gate11842(.O (I34102), .I (g25220));
INVX1 gate11843(.O (g26192), .I (I34102));
INVX1 gate11844(.O (I34105), .I (g25221));
INVX1 gate11845(.O (g26193), .I (I34105));
INVX1 gate11846(.O (I34108), .I (g25222));
INVX1 gate11847(.O (g26194), .I (I34108));
INVX1 gate11848(.O (I34111), .I (g25223));
INVX1 gate11849(.O (g26195), .I (I34111));
INVX1 gate11850(.O (I34114), .I (g25958));
INVX1 gate11851(.O (g26196), .I (I34114));
INVX1 gate11852(.O (I34118), .I (g25605));
INVX1 gate11853(.O (g26202), .I (I34118));
INVX1 gate11854(.O (I34121), .I (g25224));
INVX1 gate11855(.O (g26205), .I (I34121));
INVX1 gate11856(.O (I34124), .I (g25225));
INVX1 gate11857(.O (g26206), .I (I34124));
INVX1 gate11858(.O (I34128), .I (g25227));
INVX1 gate11859(.O (g26208), .I (I34128));
INVX1 gate11860(.O (g26209), .I (g25296));
INVX1 gate11861(.O (I34132), .I (g25228));
INVX1 gate11862(.O (g26210), .I (I34132));
INVX1 gate11863(.O (I34135), .I (g25229));
INVX1 gate11864(.O (g26211), .I (I34135));
INVX1 gate11865(.O (I34140), .I (g25230));
INVX1 gate11866(.O (g26214), .I (I34140));
INVX1 gate11867(.O (I34143), .I (g25231));
INVX1 gate11868(.O (g26215), .I (I34143));
INVX1 gate11869(.O (I34146), .I (g25232));
INVX1 gate11870(.O (g26216), .I (I34146));
INVX1 gate11871(.O (I34150), .I (g25233));
INVX1 gate11872(.O (g26220), .I (I34150));
INVX1 gate11873(.O (I34153), .I (g25234));
INVX1 gate11874(.O (g26221), .I (I34153));
INVX1 gate11875(.O (I34156), .I (g25235));
INVX1 gate11876(.O (g26222), .I (I34156));
INVX1 gate11877(.O (I34159), .I (g25964));
INVX1 gate11878(.O (g26223), .I (I34159));
INVX1 gate11879(.O (I34162), .I (g25684));
INVX1 gate11880(.O (g26226), .I (I34162));
INVX1 gate11881(.O (I34165), .I (g25236));
INVX1 gate11882(.O (g26229), .I (I34165));
INVX1 gate11883(.O (I34168), .I (g25237));
INVX1 gate11884(.O (g26230), .I (I34168));
INVX1 gate11885(.O (I34172), .I (g25239));
INVX1 gate11886(.O (g26232), .I (I34172));
INVX1 gate11887(.O (g26237), .I (g25306));
INVX1 gate11888(.O (I34180), .I (g25240));
INVX1 gate11889(.O (g26238), .I (I34180));
INVX1 gate11890(.O (I34183), .I (g25241));
INVX1 gate11891(.O (g26239), .I (I34183));
INVX1 gate11892(.O (I34189), .I (g25242));
INVX1 gate11893(.O (g26245), .I (I34189));
INVX1 gate11894(.O (I34192), .I (g25243));
INVX1 gate11895(.O (g26246), .I (I34192));
INVX1 gate11896(.O (I34195), .I (g25244));
INVX1 gate11897(.O (g26247), .I (I34195));
INVX1 gate11898(.O (I34198), .I (g25245));
INVX1 gate11899(.O (g26248), .I (I34198));
INVX1 gate11900(.O (I34201), .I (g25246));
INVX1 gate11901(.O (g26249), .I (I34201));
INVX1 gate11902(.O (I34204), .I (g25247));
INVX1 gate11903(.O (g26250), .I (I34204));
INVX1 gate11904(.O (I34207), .I (g25969));
INVX1 gate11905(.O (g26251), .I (I34207));
INVX1 gate11906(.O (I34210), .I (g25761));
INVX1 gate11907(.O (g26254), .I (I34210));
INVX1 gate11908(.O (I34220), .I (g25248));
INVX1 gate11909(.O (g26264), .I (I34220));
INVX1 gate11910(.O (g26275), .I (g25315));
INVX1 gate11911(.O (I34230), .I (g25249));
INVX1 gate11912(.O (g26276), .I (I34230));
INVX1 gate11913(.O (I34233), .I (g25250));
INVX1 gate11914(.O (g26277), .I (I34233));
INVX1 gate11915(.O (I34238), .I (g25251));
INVX1 gate11916(.O (g26280), .I (I34238));
INVX1 gate11917(.O (I34241), .I (g25252));
INVX1 gate11918(.O (g26281), .I (I34241));
INVX1 gate11919(.O (I34244), .I (g25253));
INVX1 gate11920(.O (g26282), .I (I34244));
INVX1 gate11921(.O (I34254), .I (g25185));
INVX1 gate11922(.O (g26294), .I (I34254));
INVX1 gate11923(.O (I34266), .I (g25255));
INVX1 gate11924(.O (g26308), .I (I34266));
INVX1 gate11925(.O (g26313), .I (g25324));
INVX1 gate11926(.O (I34274), .I (g25256));
INVX1 gate11927(.O (g26314), .I (I34274));
INVX1 gate11928(.O (I34277), .I (g25257));
INVX1 gate11929(.O (g26315), .I (I34277));
INVX1 gate11930(.O (I34296), .I (g25189));
INVX1 gate11931(.O (g26341), .I (I34296));
INVX1 gate11932(.O (I34306), .I (g25259));
INVX1 gate11933(.O (g26349), .I (I34306));
INVX1 gate11934(.O (I34313), .I (g25265));
INVX1 gate11935(.O (g26354), .I (I34313));
INVX1 gate11936(.O (I34316), .I (g25191));
INVX1 gate11937(.O (g26355), .I (I34316));
INVX1 gate11938(.O (I34321), .I (g25928));
INVX1 gate11939(.O (g26358), .I (I34321));
INVX1 gate11940(.O (I34327), .I (g25260));
INVX1 gate11941(.O (g26364), .I (I34327));
INVX1 gate11942(.O (I34343), .I (g25194));
INVX1 gate11943(.O (g26385), .I (I34343));
INVX1 gate11944(.O (I34353), .I (g25927));
INVX1 gate11945(.O (g26393), .I (I34353));
INVX1 gate11946(.O (I34358), .I (g25262));
INVX1 gate11947(.O (g26398), .I (I34358));
INVX1 gate11948(.O (I34363), .I (g25930));
INVX1 gate11949(.O (g26401), .I (I34363));
INVX1 gate11950(.O (I34369), .I (g25263));
INVX1 gate11951(.O (g26407), .I (I34369));
INVX1 gate11952(.O (I34385), .I (g25197));
INVX1 gate11953(.O (g26428), .I (I34385));
INVX1 gate11954(.O (I34388), .I (g25200));
INVX1 gate11955(.O (g26429), .I (I34388));
INVX1 gate11956(.O (I34392), .I (g25266));
INVX1 gate11957(.O (g26433), .I (I34392));
INVX1 gate11958(.O (I34395), .I (g25929));
INVX1 gate11959(.O (g26434), .I (I34395));
INVX1 gate11960(.O (I34400), .I (g25267));
INVX1 gate11961(.O (g26439), .I (I34400));
INVX1 gate11962(.O (I34405), .I (g25933));
INVX1 gate11963(.O (g26442), .I (I34405));
INVX1 gate11964(.O (I34411), .I (g25268));
INVX1 gate11965(.O (g26448), .I (I34411));
INVX1 gate11966(.O (I34421), .I (g25203));
INVX1 gate11967(.O (g26461), .I (I34421));
INVX1 gate11968(.O (I34425), .I (g25270));
INVX1 gate11969(.O (g26465), .I (I34425));
INVX1 gate11970(.O (I34428), .I (g25931));
INVX1 gate11971(.O (g26466), .I (I34428));
INVX1 gate11972(.O (I34433), .I (g25271));
INVX1 gate11973(.O (g26471), .I (I34433));
INVX1 gate11974(.O (I34438), .I (g25936));
INVX1 gate11975(.O (g26474), .I (I34438));
INVX1 gate11976(.O (I34444), .I (g25272));
INVX1 gate11977(.O (g26480), .I (I34444));
INVX1 gate11978(.O (g26481), .I (g25764));
INVX1 gate11979(.O (I34449), .I (g25205));
INVX1 gate11980(.O (g26485), .I (I34449));
INVX1 gate11981(.O (I34453), .I (g25279));
INVX1 gate11982(.O (g26489), .I (I34453));
INVX1 gate11983(.O (I34456), .I (g25934));
INVX1 gate11984(.O (g26490), .I (I34456));
INVX1 gate11985(.O (I34461), .I (g25280));
INVX1 gate11986(.O (g26495), .I (I34461));
INVX1 gate11987(.O (I34464), .I (g25199));
INVX1 gate11988(.O (g26496), .I (I34464));
INVX1 gate11989(.O (g26497), .I (g25818));
INVX1 gate11990(.O (I34469), .I (g25210));
INVX1 gate11991(.O (g26501), .I (I34469));
INVX1 gate11992(.O (I34473), .I (g25288));
INVX1 gate11993(.O (g26505), .I (I34473));
INVX1 gate11994(.O (I34476), .I (g25201));
INVX1 gate11995(.O (g26506), .I (I34476));
INVX1 gate11996(.O (I34479), .I (g25202));
INVX1 gate11997(.O (g26507), .I (I34479));
INVX1 gate11998(.O (g26508), .I (g25312));
INVX1 gate11999(.O (g26512), .I (g25853));
INVX1 gate12000(.O (g26516), .I (g25320));
INVX1 gate12001(.O (g26520), .I (g25874));
INVX1 gate12002(.O (g26521), .I (g25331));
INVX1 gate12003(.O (g26525), .I (g25340));
INVX1 gate12004(.O (g26533), .I (g25454));
INVX1 gate12005(.O (g26538), .I (g25458));
INVX1 gate12006(.O (g26539), .I (g25463));
INVX1 gate12007(.O (g26540), .I (g25467));
INVX1 gate12008(.O (g26542), .I (g25472));
INVX1 gate12009(.O (g26543), .I (g25476));
INVX1 gate12010(.O (g26544), .I (g25479));
INVX1 gate12011(.O (g26546), .I (g25484));
INVX1 gate12012(.O (I34505), .I (g25450));
INVX1 gate12013(.O (g26548), .I (I34505));
INVX1 gate12014(.O (g26549), .I (g25421));
INVX1 gate12015(.O (g26550), .I (g25493));
INVX1 gate12016(.O (g26551), .I (g25496));
INVX1 gate12017(.O (g26552), .I (g25499));
INVX1 gate12018(.O (g26554), .I (g25502));
INVX1 gate12019(.O (g26555), .I (g25507));
INVX1 gate12020(.O (g26556), .I (g25510));
INVX1 gate12021(.O (g26558), .I (g25515));
INVX1 gate12022(.O (g26561), .I (g25524));
INVX1 gate12023(.O (g26562), .I (g25527));
INVX1 gate12024(.O (g26563), .I (g25530));
INVX1 gate12025(.O (g26564), .I (g25533));
INVX1 gate12026(.O (g26565), .I (g25536));
INVX1 gate12027(.O (g26566), .I (g25540));
INVX1 gate12028(.O (g26567), .I (g25543));
INVX1 gate12029(.O (g26568), .I (g25546));
INVX1 gate12030(.O (g26570), .I (g25549));
INVX1 gate12031(.O (g26571), .I (g25554));
INVX1 gate12032(.O (g26572), .I (g25557));
INVX1 gate12033(.O (g26574), .I (g25562));
INVX1 gate12034(.O (I34535), .I (g25451));
INVX1 gate12035(.O (g26576), .I (I34535));
INVX1 gate12036(.O (g26577), .I (g25436));
INVX1 gate12037(.O (g26578), .I (g25573));
INVX1 gate12038(.O (g26579), .I (g25576));
INVX1 gate12039(.O (g26580), .I (g25579));
INVX1 gate12040(.O (g26581), .I (g25582));
INVX1 gate12041(.O (g26582), .I (g25585));
INVX1 gate12042(.O (g26584), .I (g25590));
INVX1 gate12043(.O (g26585), .I (g25593));
INVX1 gate12044(.O (g26586), .I (g25596));
INVX1 gate12045(.O (g26587), .I (g25599));
INVX1 gate12046(.O (g26588), .I (g25602));
INVX1 gate12047(.O (g26589), .I (g25606));
INVX1 gate12048(.O (g26590), .I (g25609));
INVX1 gate12049(.O (g26591), .I (g25612));
INVX1 gate12050(.O (g26593), .I (g25615));
INVX1 gate12051(.O (g26594), .I (g25620));
INVX1 gate12052(.O (g26595), .I (g25623));
INVX1 gate12053(.O (g26597), .I (g25443));
INVX1 gate12054(.O (g26598), .I (g25634));
INVX1 gate12055(.O (g26599), .I (g25637));
INVX1 gate12056(.O (g26600), .I (g25640));
INVX1 gate12057(.O (g26601), .I (g25643));
INVX1 gate12058(.O (g26602), .I (g25652));
INVX1 gate12059(.O (g26603), .I (g25655));
INVX1 gate12060(.O (g26604), .I (g25658));
INVX1 gate12061(.O (g26605), .I (g25661));
INVX1 gate12062(.O (g26606), .I (g25664));
INVX1 gate12063(.O (g26608), .I (g25669));
INVX1 gate12064(.O (g26609), .I (g25672));
INVX1 gate12065(.O (g26610), .I (g25675));
INVX1 gate12066(.O (g26611), .I (g25678));
INVX1 gate12067(.O (g26612), .I (g25681));
INVX1 gate12068(.O (g26613), .I (g25685));
INVX1 gate12069(.O (g26614), .I (g25688));
INVX1 gate12070(.O (g26615), .I (g25691));
INVX1 gate12071(.O (g26617), .I (g25694));
INVX1 gate12072(.O (I34579), .I (g25452));
INVX1 gate12073(.O (g26618), .I (I34579));
INVX1 gate12074(.O (g26619), .I (g25700));
INVX1 gate12075(.O (g26620), .I (g25703));
INVX1 gate12076(.O (g26621), .I (g25711));
INVX1 gate12077(.O (g26622), .I (g25714));
INVX1 gate12078(.O (g26623), .I (g25717));
INVX1 gate12079(.O (g26624), .I (g25720));
INVX1 gate12080(.O (g26625), .I (g25729));
INVX1 gate12081(.O (g26626), .I (g25732));
INVX1 gate12082(.O (g26627), .I (g25735));
INVX1 gate12083(.O (g26628), .I (g25738));
INVX1 gate12084(.O (g26629), .I (g25741));
INVX1 gate12085(.O (g26631), .I (g25746));
INVX1 gate12086(.O (g26632), .I (g25749));
INVX1 gate12087(.O (g26633), .I (g25752));
INVX1 gate12088(.O (g26634), .I (g25755));
INVX1 gate12089(.O (g26635), .I (g25758));
INVX1 gate12090(.O (g26636), .I (g25767));
INVX1 gate12091(.O (g26637), .I (g25773));
INVX1 gate12092(.O (g26638), .I (g25776));
INVX1 gate12093(.O (g26639), .I (g25784));
INVX1 gate12094(.O (g26640), .I (g25787));
INVX1 gate12095(.O (g26641), .I (g25790));
INVX1 gate12096(.O (g26642), .I (g25793));
INVX1 gate12097(.O (g26643), .I (g25802));
INVX1 gate12098(.O (g26644), .I (g25805));
INVX1 gate12099(.O (g26645), .I (g25808));
INVX1 gate12100(.O (g26646), .I (g25811));
INVX1 gate12101(.O (g26647), .I (g25814));
INVX1 gate12102(.O (g26648), .I (g25821));
INVX1 gate12103(.O (g26649), .I (g25827));
INVX1 gate12104(.O (g26650), .I (g25830));
INVX1 gate12105(.O (g26651), .I (g25838));
INVX1 gate12106(.O (g26652), .I (g25841));
INVX1 gate12107(.O (g26653), .I (g25844));
INVX1 gate12108(.O (g26654), .I (g25847));
INVX1 gate12109(.O (g26656), .I (g25856));
INVX1 gate12110(.O (g26657), .I (g25862));
INVX1 gate12111(.O (g26658), .I (g25865));
INVX1 gate12112(.O (g26662), .I (g25877));
INVX1 gate12113(.O (I34641), .I (g26086));
INVX1 gate12114(.O (g26678), .I (I34641));
INVX1 gate12115(.O (I34644), .I (g26159));
INVX1 gate12116(.O (g26679), .I (I34644));
INVX1 gate12117(.O (I34647), .I (g26164));
INVX1 gate12118(.O (g26680), .I (I34647));
INVX1 gate12119(.O (I34650), .I (g26172));
INVX1 gate12120(.O (g26681), .I (I34650));
INVX1 gate12121(.O (I34653), .I (g26165));
INVX1 gate12122(.O (g26682), .I (I34653));
INVX1 gate12123(.O (I34656), .I (g26173));
INVX1 gate12124(.O (g26683), .I (I34656));
INVX1 gate12125(.O (I34659), .I (g26190));
INVX1 gate12126(.O (g26684), .I (I34659));
INVX1 gate12127(.O (I34662), .I (g26174));
INVX1 gate12128(.O (g26685), .I (I34662));
INVX1 gate12129(.O (I34665), .I (g26191));
INVX1 gate12130(.O (g26686), .I (I34665));
INVX1 gate12131(.O (I34668), .I (g26210));
INVX1 gate12132(.O (g26687), .I (I34668));
INVX1 gate12133(.O (I34671), .I (g26192));
INVX1 gate12134(.O (g26688), .I (I34671));
INVX1 gate12135(.O (I34674), .I (g26211));
INVX1 gate12136(.O (g26689), .I (I34674));
INVX1 gate12137(.O (I34677), .I (g26232));
INVX1 gate12138(.O (g26690), .I (I34677));
INVX1 gate12139(.O (I34680), .I (g26294));
INVX1 gate12140(.O (g26691), .I (I34680));
INVX1 gate12141(.O (I34683), .I (g26364));
INVX1 gate12142(.O (g26692), .I (I34683));
INVX1 gate12143(.O (I34686), .I (g26398));
INVX1 gate12144(.O (g26693), .I (I34686));
INVX1 gate12145(.O (I34689), .I (g26433));
INVX1 gate12146(.O (g26694), .I (I34689));
INVX1 gate12147(.O (I34692), .I (g26102));
INVX1 gate12148(.O (g26695), .I (I34692));
INVX1 gate12149(.O (I34695), .I (g26167));
INVX1 gate12150(.O (g26696), .I (I34695));
INVX1 gate12151(.O (I34698), .I (g26181));
INVX1 gate12152(.O (g26697), .I (I34698));
INVX1 gate12153(.O (I34701), .I (g26193));
INVX1 gate12154(.O (g26698), .I (I34701));
INVX1 gate12155(.O (I34704), .I (g26182));
INVX1 gate12156(.O (g26699), .I (I34704));
INVX1 gate12157(.O (I34707), .I (g26194));
INVX1 gate12158(.O (g26700), .I (I34707));
INVX1 gate12159(.O (I34710), .I (g26214));
INVX1 gate12160(.O (g26701), .I (I34710));
INVX1 gate12161(.O (I34713), .I (g26195));
INVX1 gate12162(.O (g26702), .I (I34713));
INVX1 gate12163(.O (I34716), .I (g26215));
INVX1 gate12164(.O (g26703), .I (I34716));
INVX1 gate12165(.O (I34719), .I (g26238));
INVX1 gate12166(.O (g26704), .I (I34719));
INVX1 gate12167(.O (I34722), .I (g26216));
INVX1 gate12168(.O (g26705), .I (I34722));
INVX1 gate12169(.O (I34725), .I (g26239));
INVX1 gate12170(.O (g26706), .I (I34725));
INVX1 gate12171(.O (I34728), .I (g26264));
INVX1 gate12172(.O (g26707), .I (I34728));
INVX1 gate12173(.O (I34731), .I (g26341));
INVX1 gate12174(.O (g26708), .I (I34731));
INVX1 gate12175(.O (I34734), .I (g26407));
INVX1 gate12176(.O (g26709), .I (I34734));
INVX1 gate12177(.O (I34737), .I (g26439));
INVX1 gate12178(.O (g26710), .I (I34737));
INVX1 gate12179(.O (I34740), .I (g26465));
INVX1 gate12180(.O (g26711), .I (I34740));
INVX1 gate12181(.O (I34743), .I (g26118));
INVX1 gate12182(.O (g26712), .I (I34743));
INVX1 gate12183(.O (I34746), .I (g26187));
INVX1 gate12184(.O (g26713), .I (I34746));
INVX1 gate12185(.O (I34749), .I (g26205));
INVX1 gate12186(.O (g26714), .I (I34749));
INVX1 gate12187(.O (I34752), .I (g26220));
INVX1 gate12188(.O (g26715), .I (I34752));
INVX1 gate12189(.O (I34755), .I (g26206));
INVX1 gate12190(.O (g26716), .I (I34755));
INVX1 gate12191(.O (I34758), .I (g26221));
INVX1 gate12192(.O (g26717), .I (I34758));
INVX1 gate12193(.O (I34761), .I (g26245));
INVX1 gate12194(.O (g26718), .I (I34761));
INVX1 gate12195(.O (I34764), .I (g26222));
INVX1 gate12196(.O (g26719), .I (I34764));
INVX1 gate12197(.O (I34767), .I (g26246));
INVX1 gate12198(.O (g26720), .I (I34767));
INVX1 gate12199(.O (I34770), .I (g26276));
INVX1 gate12200(.O (g26721), .I (I34770));
INVX1 gate12201(.O (I34773), .I (g26247));
INVX1 gate12202(.O (g26722), .I (I34773));
INVX1 gate12203(.O (I34776), .I (g26277));
INVX1 gate12204(.O (g26723), .I (I34776));
INVX1 gate12205(.O (I34779), .I (g26308));
INVX1 gate12206(.O (g26724), .I (I34779));
INVX1 gate12207(.O (I34782), .I (g26385));
INVX1 gate12208(.O (g26725), .I (I34782));
INVX1 gate12209(.O (I34785), .I (g26448));
INVX1 gate12210(.O (g26726), .I (I34785));
INVX1 gate12211(.O (I34788), .I (g26471));
INVX1 gate12212(.O (g26727), .I (I34788));
INVX1 gate12213(.O (I34791), .I (g26489));
INVX1 gate12214(.O (g26728), .I (I34791));
INVX1 gate12215(.O (I34794), .I (g26125));
INVX1 gate12216(.O (g26729), .I (I34794));
INVX1 gate12217(.O (I34797), .I (g26208));
INVX1 gate12218(.O (g26730), .I (I34797));
INVX1 gate12219(.O (I34800), .I (g26229));
INVX1 gate12220(.O (g26731), .I (I34800));
INVX1 gate12221(.O (I34803), .I (g26248));
INVX1 gate12222(.O (g26732), .I (I34803));
INVX1 gate12223(.O (I34806), .I (g26230));
INVX1 gate12224(.O (g26733), .I (I34806));
INVX1 gate12225(.O (I34809), .I (g26249));
INVX1 gate12226(.O (g26734), .I (I34809));
INVX1 gate12227(.O (I34812), .I (g26280));
INVX1 gate12228(.O (g26735), .I (I34812));
INVX1 gate12229(.O (I34815), .I (g26250));
INVX1 gate12230(.O (g26736), .I (I34815));
INVX1 gate12231(.O (I34818), .I (g26281));
INVX1 gate12232(.O (g26737), .I (I34818));
INVX1 gate12233(.O (I34821), .I (g26314));
INVX1 gate12234(.O (g26738), .I (I34821));
INVX1 gate12235(.O (I34824), .I (g26282));
INVX1 gate12236(.O (g26739), .I (I34824));
INVX1 gate12237(.O (I34827), .I (g26315));
INVX1 gate12238(.O (g26740), .I (I34827));
INVX1 gate12239(.O (I34830), .I (g26349));
INVX1 gate12240(.O (g26741), .I (I34830));
INVX1 gate12241(.O (I34833), .I (g26428));
INVX1 gate12242(.O (g26742), .I (I34833));
INVX1 gate12243(.O (I34836), .I (g26480));
INVX1 gate12244(.O (g26743), .I (I34836));
INVX1 gate12245(.O (I34839), .I (g26495));
INVX1 gate12246(.O (g26744), .I (I34839));
INVX1 gate12247(.O (I34842), .I (g26505));
INVX1 gate12248(.O (g26745), .I (I34842));
INVX1 gate12249(.O (I34845), .I (g26496));
INVX1 gate12250(.O (g26746), .I (I34845));
INVX1 gate12251(.O (I34848), .I (g26506));
INVX1 gate12252(.O (g26747), .I (I34848));
INVX1 gate12253(.O (I34851), .I (g26354));
INVX1 gate12254(.O (g26748), .I (I34851));
INVX1 gate12255(.O (I34854), .I (g26507));
INVX1 gate12256(.O (g26749), .I (I34854));
INVX1 gate12257(.O (I34857), .I (g26355));
INVX1 gate12258(.O (g26750), .I (I34857));
INVX1 gate12259(.O (I34860), .I (g26548));
INVX1 gate12260(.O (g26751), .I (I34860));
INVX1 gate12261(.O (I34863), .I (g26576));
INVX1 gate12262(.O (g26752), .I (I34863));
INVX1 gate12263(.O (I34866), .I (g26618));
INVX1 gate12264(.O (g26753), .I (I34866));
INVX1 gate12265(.O (I34872), .I (g26217));
INVX1 gate12266(.O (g26757), .I (I34872));
INVX1 gate12267(.O (I34879), .I (g26240));
INVX1 gate12268(.O (g26762), .I (I34879));
INVX1 gate12269(.O (I34901), .I (g26295));
INVX1 gate12270(.O (g26782), .I (I34901));
INVX1 gate12271(.O (I34909), .I (g26265));
INVX1 gate12272(.O (g26788), .I (I34909));
INVX1 gate12273(.O (I34916), .I (g26240));
INVX1 gate12274(.O (g26793), .I (I34916));
INVX1 gate12275(.O (I34921), .I (g26217));
INVX1 gate12276(.O (g26796), .I (I34921));
INVX1 gate12277(.O (I34946), .I (g26534));
INVX1 gate12278(.O (g26819), .I (I34946));
INVX1 gate12279(.O (I34957), .I (g26541));
INVX1 gate12280(.O (g26828), .I (I34957));
INVX1 gate12281(.O (I34961), .I (g26545));
INVX1 gate12282(.O (g26830), .I (I34961));
INVX1 gate12283(.O (I34964), .I (g26547));
INVX1 gate12284(.O (g26831), .I (I34964));
INVX1 gate12285(.O (I34967), .I (g26553));
INVX1 gate12286(.O (g26832), .I (I34967));
INVX1 gate12287(.O (I34971), .I (g26557));
INVX1 gate12288(.O (g26834), .I (I34971));
INVX1 gate12289(.O (I34974), .I (g26168));
INVX1 gate12290(.O (g26835), .I (I34974));
INVX1 gate12291(.O (I34977), .I (g26559));
INVX1 gate12292(.O (g26836), .I (I34977));
INVX1 gate12293(.O (I34980), .I (g26458));
INVX1 gate12294(.O (g26837), .I (I34980));
INVX1 gate12295(.O (I34983), .I (g26569));
INVX1 gate12296(.O (g26840), .I (I34983));
INVX1 gate12297(.O (I34986), .I (g26160));
INVX1 gate12298(.O (g26841), .I (I34986));
INVX1 gate12299(.O (I34990), .I (g26573));
INVX1 gate12300(.O (g26843), .I (I34990));
INVX1 gate12301(.O (I34993), .I (g26575));
INVX1 gate12302(.O (g26844), .I (I34993));
INVX1 gate12303(.O (I34997), .I (g26482));
INVX1 gate12304(.O (g26846), .I (I34997));
INVX1 gate12305(.O (I35000), .I (g26336));
INVX1 gate12306(.O (g26849), .I (I35000));
INVX1 gate12307(.O (I35003), .I (g26592));
INVX1 gate12308(.O (g26850), .I (I35003));
INVX1 gate12309(.O (I35007), .I (g26596));
INVX1 gate12310(.O (g26852), .I (I35007));
INVX1 gate12311(.O (I35011), .I (g26304));
INVX1 gate12312(.O (g26854), .I (I35011));
INVX1 gate12313(.O (I35014), .I (g26498));
INVX1 gate12314(.O (g26855), .I (I35014));
INVX1 gate12315(.O (I35017), .I (g26616));
INVX1 gate12316(.O (g26858), .I (I35017));
INVX1 gate12317(.O (I35028), .I (g26513));
INVX1 gate12318(.O (g26861), .I (I35028));
INVX1 gate12319(.O (I35031), .I (g26529));
INVX1 gate12320(.O (g26864), .I (I35031));
INVX1 gate12321(.O (I35049), .I (g26530));
INVX1 gate12322(.O (g26868), .I (I35049));
INVX1 gate12323(.O (I35053), .I (g26655));
INVX1 gate12324(.O (g26872), .I (I35053));
INVX1 gate12325(.O (I35064), .I (g26531));
INVX1 gate12326(.O (g26875), .I (I35064));
INVX1 gate12327(.O (I35067), .I (g26659));
INVX1 gate12328(.O (g26876), .I (I35067));
INVX1 gate12329(.O (I35072), .I (g26661));
INVX1 gate12330(.O (g26881), .I (I35072));
INVX1 gate12331(.O (I35076), .I (g26532));
INVX1 gate12332(.O (g26883), .I (I35076));
INVX1 gate12333(.O (I35079), .I (g26664));
INVX1 gate12334(.O (g26884), .I (I35079));
INVX1 gate12335(.O (I35083), .I (g26665));
INVX1 gate12336(.O (g26886), .I (I35083));
INVX1 gate12337(.O (I35087), .I (g26667));
INVX1 gate12338(.O (g26890), .I (I35087));
INVX1 gate12339(.O (I35092), .I (g26669));
INVX1 gate12340(.O (g26895), .I (I35092));
INVX1 gate12341(.O (I35095), .I (g26670));
INVX1 gate12342(.O (g26896), .I (I35095));
INVX1 gate12343(.O (I35099), .I (g26672));
INVX1 gate12344(.O (g26900), .I (I35099));
INVX1 gate12345(.O (I35106), .I (g26675));
INVX1 gate12346(.O (g26909), .I (I35106));
INVX1 gate12347(.O (I35109), .I (g26676));
INVX1 gate12348(.O (g26910), .I (I35109));
INVX1 gate12349(.O (I35116), .I (g26025));
INVX1 gate12350(.O (g26921), .I (I35116));
INVX1 gate12351(.O (g26922), .I (g26283));
INVX1 gate12352(.O (g26935), .I (g26327));
INVX1 gate12353(.O (g26944), .I (g26374));
INVX1 gate12354(.O (g26950), .I (g26417));
INVX1 gate12355(.O (I35136), .I (g26660));
INVX1 gate12356(.O (g26953), .I (I35136));
INVX1 gate12357(.O (g26954), .I (g26549));
INVX1 gate12358(.O (I35141), .I (g26666));
INVX1 gate12359(.O (g26956), .I (I35141));
INVX1 gate12360(.O (g26957), .I (g26577));
INVX1 gate12361(.O (I35146), .I (g26671));
INVX1 gate12362(.O (g26959), .I (I35146));
INVX1 gate12363(.O (g26960), .I (g26597));
INVX1 gate12364(.O (I35153), .I (g26677));
INVX1 gate12365(.O (g26964), .I (I35153));
INVX1 gate12366(.O (I35172), .I (g26272));
INVX1 gate12367(.O (g26983), .I (I35172));
INVX1 gate12368(.O (g26987), .I (g26056));
INVX1 gate12369(.O (g27010), .I (g26063));
INVX1 gate12370(.O (g27036), .I (g26070));
INVX1 gate12371(.O (g27064), .I (g26076));
INVX1 gate12372(.O (I35254), .I (g26048));
INVX1 gate12373(.O (g27075), .I (I35254));
INVX1 gate12374(.O (I35283), .I (g26031));
INVX1 gate12375(.O (g27102), .I (I35283));
INVX1 gate12376(.O (I35297), .I (g26199));
INVX1 gate12377(.O (g27114), .I (I35297));
INVX1 gate12378(.O (I35301), .I (g26037));
INVX1 gate12379(.O (g27116), .I (I35301));
INVX1 gate12380(.O (I35313), .I (g26534));
INVX1 gate12381(.O (g27126), .I (I35313));
INVX1 gate12382(.O (I35319), .I (g26183));
INVX1 gate12383(.O (g27132), .I (I35319));
INVX1 gate12384(.O (g27133), .I (g26105));
INVX1 gate12385(.O (g27134), .I (g26175));
INVX1 gate12386(.O (g27135), .I (g26178));
INVX1 gate12387(.O (g27136), .I (g26196));
INVX1 gate12388(.O (g27137), .I (g26202));
INVX1 gate12389(.O (g27138), .I (g26223));
INVX1 gate12390(.O (g27139), .I (g26226));
INVX1 gate12391(.O (g27140), .I (g26136));
INVX1 gate12392(.O (g27141), .I (g26251));
INVX1 gate12393(.O (g27142), .I (g26254));
INVX1 gate12394(.O (g27143), .I (g26150));
INVX1 gate12395(.O (I35334), .I (g26106));
INVX1 gate12396(.O (g27145), .I (I35334));
INVX1 gate12397(.O (g27146), .I (g26358));
INVX1 gate12398(.O (g27148), .I (g26393));
INVX1 gate12399(.O (I35341), .I (g26120));
INVX1 gate12400(.O (g27150), .I (I35341));
INVX1 gate12401(.O (g27151), .I (g26401));
INVX1 gate12402(.O (g27153), .I (g26429));
INVX1 gate12403(.O (I35347), .I (g26265));
INVX1 gate12404(.O (g27154), .I (I35347));
INVX1 gate12405(.O (g27155), .I (g26434));
INVX1 gate12406(.O (I35351), .I (g26272));
INVX1 gate12407(.O (g27156), .I (I35351));
INVX1 gate12408(.O (I35355), .I (g26130));
INVX1 gate12409(.O (g27158), .I (I35355));
INVX1 gate12410(.O (g27159), .I (g26442));
INVX1 gate12411(.O (I35360), .I (g26295));
INVX1 gate12412(.O (g27161), .I (I35360));
INVX1 gate12413(.O (g27162), .I (g26461));
INVX1 gate12414(.O (I35364), .I (g26304));
INVX1 gate12415(.O (g27163), .I (I35364));
INVX1 gate12416(.O (g27164), .I (g26466));
INVX1 gate12417(.O (I35369), .I (g26144));
INVX1 gate12418(.O (g27166), .I (I35369));
INVX1 gate12419(.O (g27167), .I (g26474));
INVX1 gate12420(.O (I35373), .I (g26189));
INVX1 gate12421(.O (g27168), .I (I35373));
INVX1 gate12422(.O (I35376), .I (g26336));
INVX1 gate12423(.O (g27171), .I (I35376));
INVX1 gate12424(.O (g27172), .I (g26485));
INVX1 gate12425(.O (g27173), .I (g26490));
INVX1 gate12426(.O (I35383), .I (g26160));
INVX1 gate12427(.O (g27176), .I (I35383));
INVX1 gate12428(.O (g27177), .I (g26501));
INVX1 gate12429(.O (I35389), .I (g26168));
INVX1 gate12430(.O (g27180), .I (I35389));
INVX1 gate12431(.O (I35394), .I (g26183));
INVX1 gate12432(.O (g27183), .I (I35394));
INVX1 gate12433(.O (I35399), .I (g26199));
INVX1 gate12434(.O (g27186), .I (I35399));
INVX1 gate12435(.O (I35404), .I (g26864));
INVX1 gate12436(.O (g27189), .I (I35404));
INVX1 gate12437(.O (I35407), .I (g27145));
INVX1 gate12438(.O (g27190), .I (I35407));
INVX1 gate12439(.O (I35410), .I (g26872));
INVX1 gate12440(.O (g27191), .I (I35410));
INVX1 gate12441(.O (I35413), .I (g26876));
INVX1 gate12442(.O (g27192), .I (I35413));
INVX1 gate12443(.O (I35416), .I (g26884));
INVX1 gate12444(.O (g27193), .I (I35416));
INVX1 gate12445(.O (I35419), .I (g26828));
INVX1 gate12446(.O (g27194), .I (I35419));
INVX1 gate12447(.O (I35422), .I (g26830));
INVX1 gate12448(.O (g27195), .I (I35422));
INVX1 gate12449(.O (I35425), .I (g26832));
INVX1 gate12450(.O (g27196), .I (I35425));
INVX1 gate12451(.O (I35428), .I (g26953));
INVX1 gate12452(.O (g27197), .I (I35428));
INVX1 gate12453(.O (I35431), .I (g26868));
INVX1 gate12454(.O (g27198), .I (I35431));
INVX1 gate12455(.O (I35434), .I (g27150));
INVX1 gate12456(.O (g27199), .I (I35434));
INVX1 gate12457(.O (I35437), .I (g27183));
INVX1 gate12458(.O (g27200), .I (I35437));
INVX1 gate12459(.O (I35440), .I (g27186));
INVX1 gate12460(.O (g27201), .I (I35440));
INVX1 gate12461(.O (I35443), .I (g26757));
INVX1 gate12462(.O (g27202), .I (I35443));
INVX1 gate12463(.O (I35446), .I (g26762));
INVX1 gate12464(.O (g27203), .I (I35446));
INVX1 gate12465(.O (I35449), .I (g27154));
INVX1 gate12466(.O (g27204), .I (I35449));
INVX1 gate12467(.O (I35452), .I (g27161));
INVX1 gate12468(.O (g27205), .I (I35452));
INVX1 gate12469(.O (I35455), .I (g26881));
INVX1 gate12470(.O (g27206), .I (I35455));
INVX1 gate12471(.O (I35458), .I (g26886));
INVX1 gate12472(.O (g27207), .I (I35458));
INVX1 gate12473(.O (I35461), .I (g26895));
INVX1 gate12474(.O (g27208), .I (I35461));
INVX1 gate12475(.O (I35464), .I (g26831));
INVX1 gate12476(.O (g27209), .I (I35464));
INVX1 gate12477(.O (I35467), .I (g26834));
INVX1 gate12478(.O (g27210), .I (I35467));
INVX1 gate12479(.O (I35470), .I (g26840));
INVX1 gate12480(.O (g27211), .I (I35470));
INVX1 gate12481(.O (I35473), .I (g27156));
INVX1 gate12482(.O (g27212), .I (I35473));
INVX1 gate12483(.O (I35476), .I (g27163));
INVX1 gate12484(.O (g27213), .I (I35476));
INVX1 gate12485(.O (I35479), .I (g27171));
INVX1 gate12486(.O (g27214), .I (I35479));
INVX1 gate12487(.O (I35482), .I (g27176));
INVX1 gate12488(.O (g27215), .I (I35482));
INVX1 gate12489(.O (I35485), .I (g27180));
INVX1 gate12490(.O (g27216), .I (I35485));
INVX1 gate12491(.O (I35488), .I (g26819));
INVX1 gate12492(.O (g27217), .I (I35488));
INVX1 gate12493(.O (I35491), .I (g26956));
INVX1 gate12494(.O (g27218), .I (I35491));
INVX1 gate12495(.O (I35494), .I (g26875));
INVX1 gate12496(.O (g27219), .I (I35494));
INVX1 gate12497(.O (I35497), .I (g27158));
INVX1 gate12498(.O (g27220), .I (I35497));
INVX1 gate12499(.O (I35500), .I (g26890));
INVX1 gate12500(.O (g27221), .I (I35500));
INVX1 gate12501(.O (I35503), .I (g26896));
INVX1 gate12502(.O (g27222), .I (I35503));
INVX1 gate12503(.O (I35506), .I (g26909));
INVX1 gate12504(.O (g27223), .I (I35506));
INVX1 gate12505(.O (I35509), .I (g26836));
INVX1 gate12506(.O (g27224), .I (I35509));
INVX1 gate12507(.O (I35512), .I (g26843));
INVX1 gate12508(.O (g27225), .I (I35512));
INVX1 gate12509(.O (I35515), .I (g26850));
INVX1 gate12510(.O (g27226), .I (I35515));
INVX1 gate12511(.O (I35518), .I (g26959));
INVX1 gate12512(.O (g27227), .I (I35518));
INVX1 gate12513(.O (I35521), .I (g26883));
INVX1 gate12514(.O (g27228), .I (I35521));
INVX1 gate12515(.O (I35524), .I (g27166));
INVX1 gate12516(.O (g27229), .I (I35524));
INVX1 gate12517(.O (I35527), .I (g26900));
INVX1 gate12518(.O (g27230), .I (I35527));
INVX1 gate12519(.O (I35530), .I (g26910));
INVX1 gate12520(.O (g27231), .I (I35530));
INVX1 gate12521(.O (I35533), .I (g26921));
INVX1 gate12522(.O (g27232), .I (I35533));
INVX1 gate12523(.O (I35536), .I (g26844));
INVX1 gate12524(.O (g27233), .I (I35536));
INVX1 gate12525(.O (I35539), .I (g26852));
INVX1 gate12526(.O (g27234), .I (I35539));
INVX1 gate12527(.O (I35542), .I (g26858));
INVX1 gate12528(.O (g27235), .I (I35542));
INVX1 gate12529(.O (I35545), .I (g26964));
INVX1 gate12530(.O (g27236), .I (I35545));
INVX1 gate12531(.O (I35548), .I (g27116));
INVX1 gate12532(.O (g27237), .I (I35548));
INVX1 gate12533(.O (I35551), .I (g27075));
INVX1 gate12534(.O (g27238), .I (I35551));
INVX1 gate12535(.O (I35554), .I (g27102));
INVX1 gate12536(.O (g27239), .I (I35554));
INVX1 gate12537(.O (g27349), .I (g27126));
INVX1 gate12538(.O (I35667), .I (g27120));
INVX1 gate12539(.O (g27353), .I (I35667));
INVX1 gate12540(.O (I35673), .I (g27123));
INVX1 gate12541(.O (g27357), .I (I35673));
INVX1 gate12542(.O (I35678), .I (g27129));
INVX1 gate12543(.O (g27360), .I (I35678));
INVX1 gate12544(.O (I35681), .I (g26869));
INVX1 gate12545(.O (g27361), .I (I35681));
INVX1 gate12546(.O (I35686), .I (g27131));
INVX1 gate12547(.O (g27366), .I (I35686));
INVX1 gate12548(.O (I35689), .I (g26878));
INVX1 gate12549(.O (g27367), .I (I35689));
INVX1 gate12550(.O (I35695), .I (g26887));
INVX1 gate12551(.O (g27373), .I (I35695));
INVX1 gate12552(.O (I35698), .I (g26897));
INVX1 gate12553(.O (g27376), .I (I35698));
INVX1 gate12554(.O (I35708), .I (g26974));
INVX1 gate12555(.O (g27380), .I (I35708));
INVX1 gate12556(.O (I35711), .I (g26974));
INVX1 gate12557(.O (g27381), .I (I35711));
INVX1 gate12558(.O (g27383), .I (g27133));
INVX1 gate12559(.O (g27384), .I (g27140));
INVX1 gate12560(.O (I35723), .I (g27168));
INVX1 gate12561(.O (g27385), .I (I35723));
INVX1 gate12562(.O (g27386), .I (g27143));
INVX1 gate12563(.O (I35727), .I (g26902));
INVX1 gate12564(.O (g27387), .I (I35727));
INVX1 gate12565(.O (I35731), .I (g26892));
INVX1 gate12566(.O (g27391), .I (I35731));
INVX1 gate12567(.O (I35737), .I (g26915));
INVX1 gate12568(.O (g27397), .I (I35737));
INVX1 gate12569(.O (I35741), .I (g27118));
INVX1 gate12570(.O (g27401), .I (I35741));
INVX1 gate12571(.O (I35744), .I (g26906));
INVX1 gate12572(.O (g27404), .I (I35744));
INVX1 gate12573(.O (I35750), .I (g26928));
INVX1 gate12574(.O (g27410), .I (I35750));
INVX1 gate12575(.O (I35756), .I (g27117));
INVX1 gate12576(.O (g27416), .I (I35756));
INVX1 gate12577(.O (I35759), .I (g27121));
INVX1 gate12578(.O (g27419), .I (I35759));
INVX1 gate12579(.O (I35762), .I (g26918));
INVX1 gate12580(.O (g27422), .I (I35762));
INVX1 gate12581(.O (I35768), .I (g26941));
INVX1 gate12582(.O (g27428), .I (I35768));
INVX1 gate12583(.O (I35772), .I (g26772));
INVX1 gate12584(.O (g27432), .I (I35772));
INVX1 gate12585(.O (I35777), .I (g27119));
INVX1 gate12586(.O (g27437), .I (I35777));
INVX1 gate12587(.O (I35780), .I (g27124));
INVX1 gate12588(.O (g27440), .I (I35780));
INVX1 gate12589(.O (I35783), .I (g26931));
INVX1 gate12590(.O (g27443), .I (I35783));
INVX1 gate12591(.O (g27449), .I (g26837));
INVX1 gate12592(.O (I35791), .I (g26779));
INVX1 gate12593(.O (g27451), .I (I35791));
INVX1 gate12594(.O (I35796), .I (g27122));
INVX1 gate12595(.O (g27456), .I (I35796));
INVX1 gate12596(.O (I35799), .I (g27130));
INVX1 gate12597(.O (g27459), .I (I35799));
INVX1 gate12598(.O (I35803), .I (g26803));
INVX1 gate12599(.O (g27463), .I (I35803));
INVX1 gate12600(.O (g27465), .I (g26846));
INVX1 gate12601(.O (I35809), .I (g26785));
INVX1 gate12602(.O (g27467), .I (I35809));
INVX1 gate12603(.O (I35814), .I (g27125));
INVX1 gate12604(.O (g27472), .I (I35814));
INVX1 gate12605(.O (I35817), .I (g26922));
INVX1 gate12606(.O (g27475), .I (I35817));
INVX1 gate12607(.O (I35821), .I (g26804));
INVX1 gate12608(.O (g27479), .I (I35821));
INVX1 gate12609(.O (I35824), .I (g26805));
INVX1 gate12610(.O (g27480), .I (I35824));
INVX1 gate12611(.O (I35829), .I (g26806));
INVX1 gate12612(.O (g27483), .I (I35829));
INVX1 gate12613(.O (g27484), .I (g26855));
INVX1 gate12614(.O (I35834), .I (g26792));
INVX1 gate12615(.O (g27486), .I (I35834));
INVX1 gate12616(.O (I35837), .I (g26911));
INVX1 gate12617(.O (g27489), .I (I35837));
INVX1 gate12618(.O (I35841), .I (g26807));
INVX1 gate12619(.O (g27493), .I (I35841));
INVX1 gate12620(.O (I35844), .I (g26808));
INVX1 gate12621(.O (g27494), .I (I35844));
INVX1 gate12622(.O (I35849), .I (g26776));
INVX1 gate12623(.O (g27497), .I (I35849));
INVX1 gate12624(.O (I35852), .I (g26935));
INVX1 gate12625(.O (g27498), .I (I35852));
INVX1 gate12626(.O (I35856), .I (g26809));
INVX1 gate12627(.O (g27502), .I (I35856));
INVX1 gate12628(.O (I35859), .I (g26810));
INVX1 gate12629(.O (g27503), .I (I35859));
INVX1 gate12630(.O (I35863), .I (g26811));
INVX1 gate12631(.O (g27505), .I (I35863));
INVX1 gate12632(.O (g27506), .I (g26861));
INVX1 gate12633(.O (I35868), .I (g26812));
INVX1 gate12634(.O (g27508), .I (I35868));
INVX1 gate12635(.O (I35872), .I (g26925));
INVX1 gate12636(.O (g27510), .I (I35872));
INVX1 gate12637(.O (I35876), .I (g26813));
INVX1 gate12638(.O (g27514), .I (I35876));
INVX1 gate12639(.O (I35879), .I (g26814));
INVX1 gate12640(.O (g27515), .I (I35879));
INVX1 gate12641(.O (I35883), .I (g26781));
INVX1 gate12642(.O (g27517), .I (I35883));
INVX1 gate12643(.O (I35886), .I (g26944));
INVX1 gate12644(.O (g27518), .I (I35886));
INVX1 gate12645(.O (I35890), .I (g26815));
INVX1 gate12646(.O (g27522), .I (I35890));
INVX1 gate12647(.O (I35893), .I (g26816));
INVX1 gate12648(.O (g27523), .I (I35893));
INVX1 gate12649(.O (I35897), .I (g26817));
INVX1 gate12650(.O (g27525), .I (I35897));
INVX1 gate12651(.O (I35900), .I (g26786));
INVX1 gate12652(.O (g27526), .I (I35900));
INVX1 gate12653(.O (I35915), .I (g26818));
INVX1 gate12654(.O (g27533), .I (I35915));
INVX1 gate12655(.O (I35919), .I (g26938));
INVX1 gate12656(.O (g27535), .I (I35919));
INVX1 gate12657(.O (I35923), .I (g26820));
INVX1 gate12658(.O (g27539), .I (I35923));
INVX1 gate12659(.O (I35926), .I (g26821));
INVX1 gate12660(.O (g27540), .I (I35926));
INVX1 gate12661(.O (I35930), .I (g26789));
INVX1 gate12662(.O (g27542), .I (I35930));
INVX1 gate12663(.O (I35933), .I (g26950));
INVX1 gate12664(.O (g27543), .I (I35933));
INVX1 gate12665(.O (I35937), .I (g26822));
INVX1 gate12666(.O (g27547), .I (I35937));
INVX1 gate12667(.O (I35940), .I (g26823));
INVX1 gate12668(.O (g27548), .I (I35940));
INVX1 gate12669(.O (I35953), .I (g26824));
INVX1 gate12670(.O (g27553), .I (I35953));
INVX1 gate12671(.O (I35957), .I (g26947));
INVX1 gate12672(.O (g27555), .I (I35957));
INVX1 gate12673(.O (I35961), .I (g26825));
INVX1 gate12674(.O (g27559), .I (I35961));
INVX1 gate12675(.O (I35964), .I (g26826));
INVX1 gate12676(.O (g27560), .I (I35964));
INVX1 gate12677(.O (I35968), .I (g26795));
INVX1 gate12678(.O (g27562), .I (I35968));
INVX1 gate12679(.O (I35983), .I (g26827));
INVX1 gate12680(.O (g27569), .I (I35983));
INVX1 gate12681(.O (I36008), .I (g26798));
INVX1 gate12682(.O (g27586), .I (I36008));
INVX1 gate12683(.O (g27589), .I (g27168));
INVX1 gate12684(.O (g27590), .I (g27144));
INVX1 gate12685(.O (g27595), .I (g27149));
INVX1 gate12686(.O (g27599), .I (g27147));
INVX1 gate12687(.O (g27604), .I (g27157));
INVX1 gate12688(.O (g27608), .I (g27152));
INVX1 gate12689(.O (g27613), .I (g27165));
INVX1 gate12690(.O (g27617), .I (g27160));
INVX1 gate12691(.O (g27622), .I (g27174));
INVX1 gate12692(.O (I36032), .I (g27113));
INVX1 gate12693(.O (g27632), .I (I36032));
INVX1 gate12694(.O (I36042), .I (g26960));
INVX1 gate12695(.O (g27662), .I (I36042));
INVX1 gate12696(.O (I36046), .I (g26957));
INVX1 gate12697(.O (g27667), .I (I36046));
INVX1 gate12698(.O (I36052), .I (g26954));
INVX1 gate12699(.O (g27674), .I (I36052));
INVX1 gate12700(.O (I36060), .I (g27353));
INVX1 gate12701(.O (g27683), .I (I36060));
INVX1 gate12702(.O (I36063), .I (g27463));
INVX1 gate12703(.O (g27684), .I (I36063));
INVX1 gate12704(.O (I36066), .I (g27479));
INVX1 gate12705(.O (g27685), .I (I36066));
INVX1 gate12706(.O (I36069), .I (g27493));
INVX1 gate12707(.O (g27686), .I (I36069));
INVX1 gate12708(.O (I36072), .I (g27480));
INVX1 gate12709(.O (g27687), .I (I36072));
INVX1 gate12710(.O (I36075), .I (g27494));
INVX1 gate12711(.O (g27688), .I (I36075));
INVX1 gate12712(.O (I36078), .I (g27508));
INVX1 gate12713(.O (g27689), .I (I36078));
INVX1 gate12714(.O (I36081), .I (g27497));
INVX1 gate12715(.O (g27690), .I (I36081));
INVX1 gate12716(.O (I36084), .I (g27357));
INVX1 gate12717(.O (g27691), .I (I36084));
INVX1 gate12718(.O (I36087), .I (g27483));
INVX1 gate12719(.O (g27692), .I (I36087));
INVX1 gate12720(.O (I36090), .I (g27502));
INVX1 gate12721(.O (g27693), .I (I36090));
INVX1 gate12722(.O (I36093), .I (g27514));
INVX1 gate12723(.O (g27694), .I (I36093));
INVX1 gate12724(.O (I36096), .I (g27503));
INVX1 gate12725(.O (g27695), .I (I36096));
INVX1 gate12726(.O (I36099), .I (g27515));
INVX1 gate12727(.O (g27696), .I (I36099));
INVX1 gate12728(.O (I36102), .I (g27533));
INVX1 gate12729(.O (g27697), .I (I36102));
INVX1 gate12730(.O (I36105), .I (g27517));
INVX1 gate12731(.O (g27698), .I (I36105));
INVX1 gate12732(.O (I36108), .I (g27360));
INVX1 gate12733(.O (g27699), .I (I36108));
INVX1 gate12734(.O (I36111), .I (g27505));
INVX1 gate12735(.O (g27700), .I (I36111));
INVX1 gate12736(.O (I36114), .I (g27522));
INVX1 gate12737(.O (g27701), .I (I36114));
INVX1 gate12738(.O (I36117), .I (g27539));
INVX1 gate12739(.O (g27702), .I (I36117));
INVX1 gate12740(.O (I36120), .I (g27523));
INVX1 gate12741(.O (g27703), .I (I36120));
INVX1 gate12742(.O (I36123), .I (g27540));
INVX1 gate12743(.O (g27704), .I (I36123));
INVX1 gate12744(.O (I36126), .I (g27553));
INVX1 gate12745(.O (g27705), .I (I36126));
INVX1 gate12746(.O (I36129), .I (g27542));
INVX1 gate12747(.O (g27706), .I (I36129));
INVX1 gate12748(.O (I36132), .I (g27366));
INVX1 gate12749(.O (g27707), .I (I36132));
INVX1 gate12750(.O (I36135), .I (g27525));
INVX1 gate12751(.O (g27708), .I (I36135));
INVX1 gate12752(.O (I36138), .I (g27547));
INVX1 gate12753(.O (g27709), .I (I36138));
INVX1 gate12754(.O (I36141), .I (g27559));
INVX1 gate12755(.O (g27710), .I (I36141));
INVX1 gate12756(.O (I36144), .I (g27548));
INVX1 gate12757(.O (g27711), .I (I36144));
INVX1 gate12758(.O (I36147), .I (g27560));
INVX1 gate12759(.O (g27712), .I (I36147));
INVX1 gate12760(.O (I36150), .I (g27569));
INVX1 gate12761(.O (g27713), .I (I36150));
INVX1 gate12762(.O (I36153), .I (g27562));
INVX1 gate12763(.O (g27714), .I (I36153));
INVX1 gate12764(.O (I36156), .I (g27586));
INVX1 gate12765(.O (g27715), .I (I36156));
INVX1 gate12766(.O (I36159), .I (g27526));
INVX1 gate12767(.O (g27716), .I (I36159));
INVX1 gate12768(.O (I36162), .I (g27385));
INVX1 gate12769(.O (g27717), .I (I36162));
INVX1 gate12770(.O (g27748), .I (g27632));
INVX1 gate12771(.O (I36213), .I (g27571));
INVX1 gate12772(.O (g27776), .I (I36213));
INVX1 gate12773(.O (I36217), .I (g27580));
INVX1 gate12774(.O (g27780), .I (I36217));
INVX1 gate12775(.O (I36221), .I (g27662));
INVX1 gate12776(.O (g27784), .I (I36221));
INVX1 gate12777(.O (I36224), .I (g27589));
INVX1 gate12778(.O (g27785), .I (I36224));
INVX1 gate12779(.O (I36227), .I (g27594));
INVX1 gate12780(.O (g27786), .I (I36227));
INVX1 gate12781(.O (I36230), .I (g27583));
INVX1 gate12782(.O (g27787), .I (I36230));
INVX1 gate12783(.O (I36234), .I (g27667));
INVX1 gate12784(.O (g27791), .I (I36234));
INVX1 gate12785(.O (I36237), .I (g27662));
INVX1 gate12786(.O (g27792), .I (I36237));
INVX1 gate12787(.O (I36240), .I (g27603));
INVX1 gate12788(.O (g27793), .I (I36240));
INVX1 gate12789(.O (I36243), .I (g27587));
INVX1 gate12790(.O (g27794), .I (I36243));
INVX1 gate12791(.O (I36246), .I (g27674));
INVX1 gate12792(.O (g27797), .I (I36246));
INVX1 gate12793(.O (I36250), .I (g27612));
INVX1 gate12794(.O (g27799), .I (I36250));
INVX1 gate12795(.O (I36253), .I (g27674));
INVX1 gate12796(.O (g27800), .I (I36253));
INVX1 gate12797(.O (I36264), .I (g27621));
INVX1 gate12798(.O (g27805), .I (I36264));
INVX1 gate12799(.O (I36267), .I (g27395));
INVX1 gate12800(.O (g27806), .I (I36267));
INVX1 gate12801(.O (I36280), .I (g27390));
INVX1 gate12802(.O (g27817), .I (I36280));
INVX1 gate12803(.O (I36283), .I (g27408));
INVX1 gate12804(.O (g27820), .I (I36283));
INVX1 gate12805(.O (I36296), .I (g27626));
INVX1 gate12806(.O (g27831), .I (I36296));
INVX1 gate12807(.O (I36307), .I (g27400));
INVX1 gate12808(.O (g27839), .I (I36307));
INVX1 gate12809(.O (I36311), .I (g27426));
INVX1 gate12810(.O (g27843), .I (I36311));
INVX1 gate12811(.O (I36321), .I (g27627));
INVX1 gate12812(.O (g27847), .I (I36321));
INVX1 gate12813(.O (I36327), .I (g27413));
INVX1 gate12814(.O (g27858), .I (I36327));
INVX1 gate12815(.O (I36330), .I (g27447));
INVX1 gate12816(.O (g27861), .I (I36330));
INVX1 gate12817(.O (I36337), .I (g27628));
INVX1 gate12818(.O (g27872), .I (I36337));
INVX1 gate12819(.O (I36341), .I (g27431));
INVX1 gate12820(.O (g27879), .I (I36341));
INVX1 gate12821(.O (I36347), .I (g27630));
INVX1 gate12822(.O (g27889), .I (I36347));
INVX1 gate12823(.O (I36354), .I (g27662));
INVX1 gate12824(.O (g27903), .I (I36354));
INVX1 gate12825(.O (I36358), .I (g27672));
INVX1 gate12826(.O (g27905), .I (I36358));
INVX1 gate12827(.O (I36362), .I (g27667));
INVX1 gate12828(.O (g27907), .I (I36362));
INVX1 gate12829(.O (I36367), .I (g27678));
INVX1 gate12830(.O (g27910), .I (I36367));
INVX1 gate12831(.O (I36371), .I (g27674));
INVX1 gate12832(.O (g27912), .I (I36371));
INVX1 gate12833(.O (I36379), .I (g27682));
INVX1 gate12834(.O (g27918), .I (I36379));
INVX1 gate12835(.O (I36382), .I (g27563));
INVX1 gate12836(.O (g27919), .I (I36382));
INVX1 gate12837(.O (I36390), .I (g27243));
INVX1 gate12838(.O (g27927), .I (I36390));
INVX1 gate12839(.O (I36393), .I (g27572));
INVX1 gate12840(.O (g27928), .I (I36393));
INVX1 gate12841(.O (I36397), .I (g27574));
INVX1 gate12842(.O (g27932), .I (I36397));
INVX1 gate12843(.O (I36404), .I (g27450));
INVX1 gate12844(.O (g27939), .I (I36404));
INVX1 gate12845(.O (I36407), .I (g27581));
INVX1 gate12846(.O (g27942), .I (I36407));
INVX1 gate12847(.O (I36411), .I (g27582));
INVX1 gate12848(.O (g27946), .I (I36411));
INVX1 gate12849(.O (I36417), .I (g27462));
INVX1 gate12850(.O (g27952), .I (I36417));
INVX1 gate12851(.O (I36420), .I (g27253));
INVX1 gate12852(.O (g27955), .I (I36420));
INVX1 gate12853(.O (I36423), .I (g27466));
INVX1 gate12854(.O (g27956), .I (I36423));
INVX1 gate12855(.O (I36426), .I (g27584));
INVX1 gate12856(.O (g27959), .I (I36426));
INVX1 gate12857(.O (I36432), .I (g27585));
INVX1 gate12858(.O (g27965), .I (I36432));
INVX1 gate12859(.O (g27969), .I (g27361));
INVX1 gate12860(.O (I36438), .I (g27255));
INVX1 gate12861(.O (g27971), .I (I36438));
INVX1 gate12862(.O (I36441), .I (g27256));
INVX1 gate12863(.O (g27972), .I (I36441));
INVX1 gate12864(.O (I36444), .I (g27482));
INVX1 gate12865(.O (g27973), .I (I36444));
INVX1 gate12866(.O (I36447), .I (g27257));
INVX1 gate12867(.O (g27976), .I (I36447));
INVX1 gate12868(.O (I36450), .I (g27485));
INVX1 gate12869(.O (g27977), .I (I36450));
INVX1 gate12870(.O (I36454), .I (g27588));
INVX1 gate12871(.O (g27981), .I (I36454));
INVX1 gate12872(.O (I36459), .I (g27258));
INVX1 gate12873(.O (g27986), .I (I36459));
INVX1 gate12874(.O (I36462), .I (g27259));
INVX1 gate12875(.O (g27987), .I (I36462));
INVX1 gate12876(.O (I36465), .I (g27260));
INVX1 gate12877(.O (g27988), .I (I36465));
INVX1 gate12878(.O (I36468), .I (g27261));
INVX1 gate12879(.O (g27989), .I (I36468));
INVX1 gate12880(.O (g27990), .I (g27367));
INVX1 gate12881(.O (I36473), .I (g27262));
INVX1 gate12882(.O (g27992), .I (I36473));
INVX1 gate12883(.O (I36476), .I (g27263));
INVX1 gate12884(.O (g27993), .I (I36476));
INVX1 gate12885(.O (I36479), .I (g27504));
INVX1 gate12886(.O (g27994), .I (I36479));
INVX1 gate12887(.O (I36483), .I (g27264));
INVX1 gate12888(.O (g27998), .I (I36483));
INVX1 gate12889(.O (I36486), .I (g27507));
INVX1 gate12890(.O (g27999), .I (I36486));
INVX1 gate12891(.O (I36490), .I (g27265));
INVX1 gate12892(.O (g28003), .I (I36490));
INVX1 gate12893(.O (I36493), .I (g27266));
INVX1 gate12894(.O (g28004), .I (I36493));
INVX1 gate12895(.O (I36496), .I (g27267));
INVX1 gate12896(.O (g28005), .I (I36496));
INVX1 gate12897(.O (I36499), .I (g27268));
INVX1 gate12898(.O (g28006), .I (I36499));
INVX1 gate12899(.O (I36502), .I (g27269));
INVX1 gate12900(.O (g28007), .I (I36502));
INVX1 gate12901(.O (I36507), .I (g27270));
INVX1 gate12902(.O (g28010), .I (I36507));
INVX1 gate12903(.O (I36510), .I (g27271));
INVX1 gate12904(.O (g28011), .I (I36510));
INVX1 gate12905(.O (I36513), .I (g27272));
INVX1 gate12906(.O (g28012), .I (I36513));
INVX1 gate12907(.O (I36516), .I (g27273));
INVX1 gate12908(.O (g28013), .I (I36516));
INVX1 gate12909(.O (g28014), .I (g27373));
INVX1 gate12910(.O (I36521), .I (g27274));
INVX1 gate12911(.O (g28016), .I (I36521));
INVX1 gate12912(.O (I36524), .I (g27275));
INVX1 gate12913(.O (g28017), .I (I36524));
INVX1 gate12914(.O (I36527), .I (g27524));
INVX1 gate12915(.O (g28018), .I (I36527));
INVX1 gate12916(.O (I36530), .I (g27276));
INVX1 gate12917(.O (g28021), .I (I36530));
INVX1 gate12918(.O (I36533), .I (g27277));
INVX1 gate12919(.O (g28022), .I (I36533));
INVX1 gate12920(.O (I36536), .I (g27278));
INVX1 gate12921(.O (g28023), .I (I36536));
INVX1 gate12922(.O (I36539), .I (g27279));
INVX1 gate12923(.O (g28024), .I (I36539));
INVX1 gate12924(.O (I36542), .I (g27280));
INVX1 gate12925(.O (g28025), .I (I36542));
INVX1 gate12926(.O (I36545), .I (g27281));
INVX1 gate12927(.O (g28026), .I (I36545));
INVX1 gate12928(.O (I36551), .I (g27282));
INVX1 gate12929(.O (g28030), .I (I36551));
INVX1 gate12930(.O (I36554), .I (g27283));
INVX1 gate12931(.O (g28031), .I (I36554));
INVX1 gate12932(.O (I36557), .I (g27284));
INVX1 gate12933(.O (g28032), .I (I36557));
INVX1 gate12934(.O (I36560), .I (g27285));
INVX1 gate12935(.O (g28033), .I (I36560));
INVX1 gate12936(.O (I36563), .I (g27286));
INVX1 gate12937(.O (g28034), .I (I36563));
INVX1 gate12938(.O (I36568), .I (g27287));
INVX1 gate12939(.O (g28037), .I (I36568));
INVX1 gate12940(.O (I36571), .I (g27288));
INVX1 gate12941(.O (g28038), .I (I36571));
INVX1 gate12942(.O (I36574), .I (g27289));
INVX1 gate12943(.O (g28039), .I (I36574));
INVX1 gate12944(.O (I36577), .I (g27290));
INVX1 gate12945(.O (g28040), .I (I36577));
INVX1 gate12946(.O (g28041), .I (g27376));
INVX1 gate12947(.O (I36582), .I (g27291));
INVX1 gate12948(.O (g28043), .I (I36582));
INVX1 gate12949(.O (I36585), .I (g27292));
INVX1 gate12950(.O (g28044), .I (I36585));
INVX1 gate12951(.O (I36588), .I (g27293));
INVX1 gate12952(.O (g28045), .I (I36588));
INVX1 gate12953(.O (I36598), .I (g27294));
INVX1 gate12954(.O (g28047), .I (I36598));
INVX1 gate12955(.O (I36601), .I (g27295));
INVX1 gate12956(.O (g28048), .I (I36601));
INVX1 gate12957(.O (I36604), .I (g27296));
INVX1 gate12958(.O (g28049), .I (I36604));
INVX1 gate12959(.O (I36609), .I (g27297));
INVX1 gate12960(.O (g28052), .I (I36609));
INVX1 gate12961(.O (I36612), .I (g27298));
INVX1 gate12962(.O (g28053), .I (I36612));
INVX1 gate12963(.O (I36615), .I (g27299));
INVX1 gate12964(.O (g28054), .I (I36615));
INVX1 gate12965(.O (I36618), .I (g27300));
INVX1 gate12966(.O (g28055), .I (I36618));
INVX1 gate12967(.O (I36621), .I (g27301));
INVX1 gate12968(.O (g28056), .I (I36621));
INVX1 gate12969(.O (I36627), .I (g27302));
INVX1 gate12970(.O (g28060), .I (I36627));
INVX1 gate12971(.O (I36630), .I (g27303));
INVX1 gate12972(.O (g28061), .I (I36630));
INVX1 gate12973(.O (I36633), .I (g27304));
INVX1 gate12974(.O (g28062), .I (I36633));
INVX1 gate12975(.O (I36636), .I (g27305));
INVX1 gate12976(.O (g28063), .I (I36636));
INVX1 gate12977(.O (I36639), .I (g27306));
INVX1 gate12978(.O (g28064), .I (I36639));
INVX1 gate12979(.O (I36644), .I (g27307));
INVX1 gate12980(.O (g28067), .I (I36644));
INVX1 gate12981(.O (I36647), .I (g27308));
INVX1 gate12982(.O (g28068), .I (I36647));
INVX1 gate12983(.O (I36650), .I (g27309));
INVX1 gate12984(.O (g28069), .I (I36650));
INVX1 gate12985(.O (I36653), .I (g27310));
INVX1 gate12986(.O (g28070), .I (I36653));
INVX1 gate12987(.O (I36656), .I (g27311));
INVX1 gate12988(.O (g28071), .I (I36656));
INVX1 gate12989(.O (I36659), .I (g27312));
INVX1 gate12990(.O (g28072), .I (I36659));
INVX1 gate12991(.O (I36663), .I (g27313));
INVX1 gate12992(.O (g28074), .I (I36663));
INVX1 gate12993(.O (I36673), .I (g27314));
INVX1 gate12994(.O (g28076), .I (I36673));
INVX1 gate12995(.O (I36676), .I (g27315));
INVX1 gate12996(.O (g28077), .I (I36676));
INVX1 gate12997(.O (I36679), .I (g27316));
INVX1 gate12998(.O (g28078), .I (I36679));
INVX1 gate12999(.O (I36684), .I (g27317));
INVX1 gate13000(.O (g28081), .I (I36684));
INVX1 gate13001(.O (I36687), .I (g27318));
INVX1 gate13002(.O (g28082), .I (I36687));
INVX1 gate13003(.O (I36690), .I (g27319));
INVX1 gate13004(.O (g28083), .I (I36690));
INVX1 gate13005(.O (I36693), .I (g27320));
INVX1 gate13006(.O (g28084), .I (I36693));
INVX1 gate13007(.O (I36696), .I (g27321));
INVX1 gate13008(.O (g28085), .I (I36696));
INVX1 gate13009(.O (I36702), .I (g27322));
INVX1 gate13010(.O (g28089), .I (I36702));
INVX1 gate13011(.O (I36705), .I (g27323));
INVX1 gate13012(.O (g28090), .I (I36705));
INVX1 gate13013(.O (I36708), .I (g27324));
INVX1 gate13014(.O (g28091), .I (I36708));
INVX1 gate13015(.O (I36711), .I (g27325));
INVX1 gate13016(.O (g28092), .I (I36711));
INVX1 gate13017(.O (I36714), .I (g27326));
INVX1 gate13018(.O (g28093), .I (I36714));
INVX1 gate13019(.O (I36718), .I (g27327));
INVX1 gate13020(.O (g28095), .I (I36718));
INVX1 gate13021(.O (I36721), .I (g27328));
INVX1 gate13022(.O (g28096), .I (I36721));
INVX1 gate13023(.O (I36724), .I (g27329));
INVX1 gate13024(.O (g28097), .I (I36724));
INVX1 gate13025(.O (I36728), .I (g27330));
INVX1 gate13026(.O (g28099), .I (I36728));
INVX1 gate13027(.O (I36738), .I (g27331));
INVX1 gate13028(.O (g28101), .I (I36738));
INVX1 gate13029(.O (I36741), .I (g27332));
INVX1 gate13030(.O (g28102), .I (I36741));
INVX1 gate13031(.O (I36744), .I (g27333));
INVX1 gate13032(.O (g28103), .I (I36744));
INVX1 gate13033(.O (I36749), .I (g27334));
INVX1 gate13034(.O (g28106), .I (I36749));
INVX1 gate13035(.O (I36752), .I (g27335));
INVX1 gate13036(.O (g28107), .I (I36752));
INVX1 gate13037(.O (I36755), .I (g27336));
INVX1 gate13038(.O (g28108), .I (I36755));
INVX1 gate13039(.O (I36758), .I (g27337));
INVX1 gate13040(.O (g28109), .I (I36758));
INVX1 gate13041(.O (I36761), .I (g27338));
INVX1 gate13042(.O (g28110), .I (I36761));
INVX1 gate13043(.O (I36766), .I (g27339));
INVX1 gate13044(.O (g28113), .I (I36766));
INVX1 gate13045(.O (I36769), .I (g27340));
INVX1 gate13046(.O (g28114), .I (I36769));
INVX1 gate13047(.O (I36772), .I (g27341));
INVX1 gate13048(.O (g28115), .I (I36772));
INVX1 gate13049(.O (I36776), .I (g27342));
INVX1 gate13050(.O (g28117), .I (I36776));
INVX1 gate13051(.O (I36786), .I (g27343));
INVX1 gate13052(.O (g28119), .I (I36786));
INVX1 gate13053(.O (I36789), .I (g27344));
INVX1 gate13054(.O (g28120), .I (I36789));
INVX1 gate13055(.O (I36792), .I (g27345));
INVX1 gate13056(.O (g28121), .I (I36792));
INVX1 gate13057(.O (I36797), .I (g27346));
INVX1 gate13058(.O (g28124), .I (I36797));
INVX1 gate13059(.O (I36800), .I (g27347));
INVX1 gate13060(.O (g28125), .I (I36800));
INVX1 gate13061(.O (I36803), .I (g27348));
INVX1 gate13062(.O (g28126), .I (I36803));
INVX1 gate13063(.O (g28128), .I (g27528));
INVX1 gate13064(.O (I36808), .I (g27354));
INVX1 gate13065(.O (g28132), .I (I36808));
INVX1 gate13066(.O (g28133), .I (g27550));
INVX1 gate13067(.O (g28137), .I (g27566));
INVX1 gate13068(.O (g28141), .I (g27576));
INVX1 gate13069(.O (g28149), .I (g27667));
INVX1 gate13070(.O (g28150), .I (g27387));
INVX1 gate13071(.O (g28151), .I (g27381));
INVX1 gate13072(.O (g28152), .I (g27391));
INVX1 gate13073(.O (g28153), .I (g27397));
INVX1 gate13074(.O (g28154), .I (g27401));
INVX1 gate13075(.O (g28155), .I (g27404));
INVX1 gate13076(.O (g28156), .I (g27410));
INVX1 gate13077(.O (g28158), .I (g27416));
INVX1 gate13078(.O (g28159), .I (g27419));
INVX1 gate13079(.O (g28160), .I (g27422));
INVX1 gate13080(.O (g28161), .I (g27428));
INVX1 gate13081(.O (g28162), .I (g27432));
INVX1 gate13082(.O (g28163), .I (g27437));
INVX1 gate13083(.O (g28164), .I (g27440));
INVX1 gate13084(.O (g28165), .I (g27443));
INVX1 gate13085(.O (g28166), .I (g27451));
INVX1 gate13086(.O (g28167), .I (g27456));
INVX1 gate13087(.O (g28168), .I (g27459));
INVX1 gate13088(.O (g28169), .I (g27467));
INVX1 gate13089(.O (g28170), .I (g27472));
INVX1 gate13090(.O (g28172), .I (g27475));
INVX1 gate13091(.O (g28173), .I (g27486));
INVX1 gate13092(.O (g28174), .I (g27489));
INVX1 gate13093(.O (g28175), .I (g27498));
INVX1 gate13094(.O (g28177), .I (g27510));
INVX1 gate13095(.O (g28178), .I (g27518));
INVX1 gate13096(.O (I36848), .I (g27383));
INVX1 gate13097(.O (g28179), .I (I36848));
INVX1 gate13098(.O (g28186), .I (g27535));
INVX1 gate13099(.O (g28187), .I (g27543));
INVX1 gate13100(.O (g28190), .I (g27555));
INVX1 gate13101(.O (I36860), .I (g27386));
INVX1 gate13102(.O (g28194), .I (I36860));
INVX1 gate13103(.O (I36864), .I (g27384));
INVX1 gate13104(.O (g28200), .I (I36864));
INVX1 gate13105(.O (I36867), .I (g27786));
INVX1 gate13106(.O (g28206), .I (I36867));
INVX1 gate13107(.O (I36870), .I (g27955));
INVX1 gate13108(.O (g28207), .I (I36870));
INVX1 gate13109(.O (I36873), .I (g27971));
INVX1 gate13110(.O (g28208), .I (I36873));
INVX1 gate13111(.O (I36876), .I (g27986));
INVX1 gate13112(.O (g28209), .I (I36876));
INVX1 gate13113(.O (I36879), .I (g27972));
INVX1 gate13114(.O (g28210), .I (I36879));
INVX1 gate13115(.O (I36882), .I (g27987));
INVX1 gate13116(.O (g28211), .I (I36882));
INVX1 gate13117(.O (I36885), .I (g28003));
INVX1 gate13118(.O (g28212), .I (I36885));
INVX1 gate13119(.O (I36888), .I (g27988));
INVX1 gate13120(.O (g28213), .I (I36888));
INVX1 gate13121(.O (I36891), .I (g28004));
INVX1 gate13122(.O (g28214), .I (I36891));
INVX1 gate13123(.O (I36894), .I (g28022));
INVX1 gate13124(.O (g28215), .I (I36894));
INVX1 gate13125(.O (I36897), .I (g28005));
INVX1 gate13126(.O (g28216), .I (I36897));
INVX1 gate13127(.O (I36900), .I (g28023));
INVX1 gate13128(.O (g28217), .I (I36900));
INVX1 gate13129(.O (I36903), .I (g28045));
INVX1 gate13130(.O (g28218), .I (I36903));
INVX1 gate13131(.O (I36906), .I (g27989));
INVX1 gate13132(.O (g28219), .I (I36906));
INVX1 gate13133(.O (I36909), .I (g28006));
INVX1 gate13134(.O (g28220), .I (I36909));
INVX1 gate13135(.O (I36912), .I (g28024));
INVX1 gate13136(.O (g28221), .I (I36912));
INVX1 gate13137(.O (I36915), .I (g28007));
INVX1 gate13138(.O (g28222), .I (I36915));
INVX1 gate13139(.O (I36918), .I (g28025));
INVX1 gate13140(.O (g28223), .I (I36918));
INVX1 gate13141(.O (I36921), .I (g28047));
INVX1 gate13142(.O (g28224), .I (I36921));
INVX1 gate13143(.O (I36924), .I (g28026));
INVX1 gate13144(.O (g28225), .I (I36924));
INVX1 gate13145(.O (I36927), .I (g28048));
INVX1 gate13146(.O (g28226), .I (I36927));
INVX1 gate13147(.O (I36930), .I (g28071));
INVX1 gate13148(.O (g28227), .I (I36930));
INVX1 gate13149(.O (I36933), .I (g28049));
INVX1 gate13150(.O (g28228), .I (I36933));
INVX1 gate13151(.O (I36936), .I (g28072));
INVX1 gate13152(.O (g28229), .I (I36936));
INVX1 gate13153(.O (I36939), .I (g28095));
INVX1 gate13154(.O (g28230), .I (I36939));
INVX1 gate13155(.O (I36942), .I (g27905));
INVX1 gate13156(.O (g28231), .I (I36942));
INVX1 gate13157(.O (I36945), .I (g27793));
INVX1 gate13158(.O (g28232), .I (I36945));
INVX1 gate13159(.O (I36948), .I (g27976));
INVX1 gate13160(.O (g28233), .I (I36948));
INVX1 gate13161(.O (I36951), .I (g27992));
INVX1 gate13162(.O (g28234), .I (I36951));
INVX1 gate13163(.O (I36954), .I (g28010));
INVX1 gate13164(.O (g28235), .I (I36954));
INVX1 gate13165(.O (I36957), .I (g27993));
INVX1 gate13166(.O (g28236), .I (I36957));
INVX1 gate13167(.O (I36960), .I (g28011));
INVX1 gate13168(.O (g28237), .I (I36960));
INVX1 gate13169(.O (I36963), .I (g28030));
INVX1 gate13170(.O (g28238), .I (I36963));
INVX1 gate13171(.O (I36966), .I (g28012));
INVX1 gate13172(.O (g28239), .I (I36966));
INVX1 gate13173(.O (I36969), .I (g28031));
INVX1 gate13174(.O (g28240), .I (I36969));
INVX1 gate13175(.O (I36972), .I (g28052));
INVX1 gate13176(.O (g28241), .I (I36972));
INVX1 gate13177(.O (I36975), .I (g28032));
INVX1 gate13178(.O (g28242), .I (I36975));
INVX1 gate13179(.O (I36978), .I (g28053));
INVX1 gate13180(.O (g28243), .I (I36978));
INVX1 gate13181(.O (I36981), .I (g28074));
INVX1 gate13182(.O (g28244), .I (I36981));
INVX1 gate13183(.O (I36984), .I (g28013));
INVX1 gate13184(.O (g28245), .I (I36984));
INVX1 gate13185(.O (I36987), .I (g28033));
INVX1 gate13186(.O (g28246), .I (I36987));
INVX1 gate13187(.O (I36990), .I (g28054));
INVX1 gate13188(.O (g28247), .I (I36990));
INVX1 gate13189(.O (I36993), .I (g28034));
INVX1 gate13190(.O (g28248), .I (I36993));
INVX1 gate13191(.O (I36996), .I (g28055));
INVX1 gate13192(.O (g28249), .I (I36996));
INVX1 gate13193(.O (I36999), .I (g28076));
INVX1 gate13194(.O (g28250), .I (I36999));
INVX1 gate13195(.O (I37002), .I (g28056));
INVX1 gate13196(.O (g28251), .I (I37002));
INVX1 gate13197(.O (I37005), .I (g28077));
INVX1 gate13198(.O (g28252), .I (I37005));
INVX1 gate13199(.O (I37008), .I (g28096));
INVX1 gate13200(.O (g28253), .I (I37008));
INVX1 gate13201(.O (I37011), .I (g28078));
INVX1 gate13202(.O (g28254), .I (I37011));
INVX1 gate13203(.O (I37014), .I (g28097));
INVX1 gate13204(.O (g28255), .I (I37014));
INVX1 gate13205(.O (I37017), .I (g28113));
INVX1 gate13206(.O (g28256), .I (I37017));
INVX1 gate13207(.O (I37020), .I (g27910));
INVX1 gate13208(.O (g28257), .I (I37020));
INVX1 gate13209(.O (I37023), .I (g27799));
INVX1 gate13210(.O (g28258), .I (I37023));
INVX1 gate13211(.O (I37026), .I (g27998));
INVX1 gate13212(.O (g28259), .I (I37026));
INVX1 gate13213(.O (I37029), .I (g28016));
INVX1 gate13214(.O (g28260), .I (I37029));
INVX1 gate13215(.O (I37032), .I (g28037));
INVX1 gate13216(.O (g28261), .I (I37032));
INVX1 gate13217(.O (I37035), .I (g28017));
INVX1 gate13218(.O (g28262), .I (I37035));
INVX1 gate13219(.O (I37038), .I (g28038));
INVX1 gate13220(.O (g28263), .I (I37038));
INVX1 gate13221(.O (I37041), .I (g28060));
INVX1 gate13222(.O (g28264), .I (I37041));
INVX1 gate13223(.O (I37044), .I (g28039));
INVX1 gate13224(.O (g28265), .I (I37044));
INVX1 gate13225(.O (I37047), .I (g28061));
INVX1 gate13226(.O (g28266), .I (I37047));
INVX1 gate13227(.O (I37050), .I (g28081));
INVX1 gate13228(.O (g28267), .I (I37050));
INVX1 gate13229(.O (I37053), .I (g28062));
INVX1 gate13230(.O (g28268), .I (I37053));
INVX1 gate13231(.O (I37056), .I (g28082));
INVX1 gate13232(.O (g28269), .I (I37056));
INVX1 gate13233(.O (I37059), .I (g28099));
INVX1 gate13234(.O (g28270), .I (I37059));
INVX1 gate13235(.O (I37062), .I (g28040));
INVX1 gate13236(.O (g28271), .I (I37062));
INVX1 gate13237(.O (I37065), .I (g28063));
INVX1 gate13238(.O (g28272), .I (I37065));
INVX1 gate13239(.O (I37068), .I (g28083));
INVX1 gate13240(.O (g28273), .I (I37068));
INVX1 gate13241(.O (I37071), .I (g28064));
INVX1 gate13242(.O (g28274), .I (I37071));
INVX1 gate13243(.O (I37074), .I (g28084));
INVX1 gate13244(.O (g28275), .I (I37074));
INVX1 gate13245(.O (I37077), .I (g28101));
INVX1 gate13246(.O (g28276), .I (I37077));
INVX1 gate13247(.O (I37080), .I (g28085));
INVX1 gate13248(.O (g28277), .I (I37080));
INVX1 gate13249(.O (I37083), .I (g28102));
INVX1 gate13250(.O (g28278), .I (I37083));
INVX1 gate13251(.O (I37086), .I (g28114));
INVX1 gate13252(.O (g28279), .I (I37086));
INVX1 gate13253(.O (I37089), .I (g28103));
INVX1 gate13254(.O (g28280), .I (I37089));
INVX1 gate13255(.O (I37092), .I (g28115));
INVX1 gate13256(.O (g28281), .I (I37092));
INVX1 gate13257(.O (I37095), .I (g28124));
INVX1 gate13258(.O (g28282), .I (I37095));
INVX1 gate13259(.O (I37098), .I (g27918));
INVX1 gate13260(.O (g28283), .I (I37098));
INVX1 gate13261(.O (I37101), .I (g27805));
INVX1 gate13262(.O (g28284), .I (I37101));
INVX1 gate13263(.O (I37104), .I (g28021));
INVX1 gate13264(.O (g28285), .I (I37104));
INVX1 gate13265(.O (I37107), .I (g28043));
INVX1 gate13266(.O (g28286), .I (I37107));
INVX1 gate13267(.O (I37110), .I (g28067));
INVX1 gate13268(.O (g28287), .I (I37110));
INVX1 gate13269(.O (I37113), .I (g28044));
INVX1 gate13270(.O (g28288), .I (I37113));
INVX1 gate13271(.O (I37116), .I (g28068));
INVX1 gate13272(.O (g28289), .I (I37116));
INVX1 gate13273(.O (I37119), .I (g28089));
INVX1 gate13274(.O (g28290), .I (I37119));
INVX1 gate13275(.O (I37122), .I (g28069));
INVX1 gate13276(.O (g28291), .I (I37122));
INVX1 gate13277(.O (I37125), .I (g28090));
INVX1 gate13278(.O (g28292), .I (I37125));
INVX1 gate13279(.O (I37128), .I (g28106));
INVX1 gate13280(.O (g28293), .I (I37128));
INVX1 gate13281(.O (I37131), .I (g28091));
INVX1 gate13282(.O (g28294), .I (I37131));
INVX1 gate13283(.O (I37134), .I (g28107));
INVX1 gate13284(.O (g28295), .I (I37134));
INVX1 gate13285(.O (I37137), .I (g28117));
INVX1 gate13286(.O (g28296), .I (I37137));
INVX1 gate13287(.O (I37140), .I (g28070));
INVX1 gate13288(.O (g28297), .I (I37140));
INVX1 gate13289(.O (I37143), .I (g28092));
INVX1 gate13290(.O (g28298), .I (I37143));
INVX1 gate13291(.O (I37146), .I (g28108));
INVX1 gate13292(.O (g28299), .I (I37146));
INVX1 gate13293(.O (I37149), .I (g28093));
INVX1 gate13294(.O (g28300), .I (I37149));
INVX1 gate13295(.O (I37152), .I (g28109));
INVX1 gate13296(.O (g28301), .I (I37152));
INVX1 gate13297(.O (I37155), .I (g28119));
INVX1 gate13298(.O (g28302), .I (I37155));
INVX1 gate13299(.O (I37158), .I (g28110));
INVX1 gate13300(.O (g28303), .I (I37158));
INVX1 gate13301(.O (I37161), .I (g28120));
INVX1 gate13302(.O (g28304), .I (I37161));
INVX1 gate13303(.O (I37164), .I (g28125));
INVX1 gate13304(.O (g28305), .I (I37164));
INVX1 gate13305(.O (I37167), .I (g28121));
INVX1 gate13306(.O (g28306), .I (I37167));
INVX1 gate13307(.O (I37170), .I (g28126));
INVX1 gate13308(.O (g28307), .I (I37170));
INVX1 gate13309(.O (I37173), .I (g28132));
INVX1 gate13310(.O (g28308), .I (I37173));
INVX1 gate13311(.O (I37176), .I (g27927));
INVX1 gate13312(.O (g28309), .I (I37176));
INVX1 gate13313(.O (I37179), .I (g27784));
INVX1 gate13314(.O (g28310), .I (I37179));
INVX1 gate13315(.O (I37182), .I (g27791));
INVX1 gate13316(.O (g28311), .I (I37182));
INVX1 gate13317(.O (I37185), .I (g27797));
INVX1 gate13318(.O (g28312), .I (I37185));
INVX1 gate13319(.O (I37188), .I (g27785));
INVX1 gate13320(.O (g28313), .I (I37188));
INVX1 gate13321(.O (I37191), .I (g27792));
INVX1 gate13322(.O (g28314), .I (I37191));
INVX1 gate13323(.O (I37194), .I (g27800));
INVX1 gate13324(.O (g28315), .I (I37194));
INVX1 gate13325(.O (I37197), .I (g27903));
INVX1 gate13326(.O (g28316), .I (I37197));
INVX1 gate13327(.O (I37200), .I (g27907));
INVX1 gate13328(.O (g28317), .I (I37200));
INVX1 gate13329(.O (I37203), .I (g27912));
INVX1 gate13330(.O (g28318), .I (I37203));
INVX1 gate13331(.O (I37228), .I (g28194));
INVX1 gate13332(.O (g28341), .I (I37228));
INVX1 gate13333(.O (I37232), .I (g28200));
INVX1 gate13334(.O (g28343), .I (I37232));
INVX1 gate13335(.O (I37238), .I (g28179));
INVX1 gate13336(.O (g28347), .I (I37238));
INVX1 gate13337(.O (I37252), .I (g28200));
INVX1 gate13338(.O (g28359), .I (I37252));
INVX1 gate13339(.O (I37260), .I (g28179));
INVX1 gate13340(.O (g28365), .I (I37260));
INVX1 gate13341(.O (I37266), .I (g28200));
INVX1 gate13342(.O (g28369), .I (I37266));
INVX1 gate13343(.O (I37269), .I (g28145));
INVX1 gate13344(.O (g28370), .I (I37269));
INVX1 gate13345(.O (I37273), .I (g28179));
INVX1 gate13346(.O (g28372), .I (I37273));
INVX1 gate13347(.O (I37277), .I (g28146));
INVX1 gate13348(.O (g28374), .I (I37277));
INVX1 gate13349(.O (I37280), .I (g28179));
INVX1 gate13350(.O (g28375), .I (I37280));
INVX1 gate13351(.O (I37284), .I (g28147));
INVX1 gate13352(.O (g28377), .I (I37284));
INVX1 gate13353(.O (I37291), .I (g28148));
INVX1 gate13354(.O (g28382), .I (I37291));
INVX1 gate13355(.O (I37319), .I (g28149));
INVX1 gate13356(.O (g28390), .I (I37319));
INVX1 gate13357(.O (I37330), .I (g28194));
INVX1 gate13358(.O (g28393), .I (I37330));
INVX1 gate13359(.O (I37334), .I (g28194));
INVX1 gate13360(.O (g28395), .I (I37334));
INVX1 gate13361(.O (g28419), .I (g28151));
INVX1 gate13362(.O (I37379), .I (g28199));
INVX1 gate13363(.O (g28432), .I (I37379));
INVX1 gate13364(.O (I37386), .I (g28194));
INVX1 gate13365(.O (g28437), .I (I37386));
INVX1 gate13366(.O (I37394), .I (g27718));
INVX1 gate13367(.O (g28443), .I (I37394));
INVX1 gate13368(.O (I37400), .I (g28200));
INVX1 gate13369(.O (g28447), .I (I37400));
INVX1 gate13370(.O (I37410), .I (g27722));
INVX1 gate13371(.O (g28455), .I (I37410));
INVX1 gate13372(.O (I37415), .I (g28179));
INVX1 gate13373(.O (g28458), .I (I37415));
INVX1 gate13374(.O (I37426), .I (g27724));
INVX1 gate13375(.O (g28467), .I (I37426));
INVX1 gate13376(.O (g28483), .I (g27776));
INVX1 gate13377(.O (g28491), .I (g27780));
INVX1 gate13378(.O (g28496), .I (g27787));
INVX1 gate13379(.O (I37459), .I (g27759));
INVX1 gate13380(.O (g28498), .I (I37459));
INVX1 gate13381(.O (g28500), .I (g27794));
INVX1 gate13382(.O (I37467), .I (g27760));
INVX1 gate13383(.O (g28524), .I (I37467));
INVX1 gate13384(.O (I37471), .I (g27761));
INVX1 gate13385(.O (g28526), .I (I37471));
INVX1 gate13386(.O (I37474), .I (g27762));
INVX1 gate13387(.O (g28527), .I (I37474));
INVX1 gate13388(.O (I37481), .I (g27763));
INVX1 gate13389(.O (g28552), .I (I37481));
INVX1 gate13390(.O (I37484), .I (g27764));
INVX1 gate13391(.O (g28553), .I (I37484));
INVX1 gate13392(.O (g28554), .I (g27806));
INVX1 gate13393(.O (I37488), .I (g27765));
INVX1 gate13394(.O (g28555), .I (I37488));
INVX1 gate13395(.O (I37494), .I (g27766));
INVX1 gate13396(.O (g28579), .I (I37494));
INVX1 gate13397(.O (I37497), .I (g27767));
INVX1 gate13398(.O (g28580), .I (I37497));
INVX1 gate13399(.O (g28581), .I (g27817));
INVX1 gate13400(.O (g28582), .I (g27820));
INVX1 gate13401(.O (I37502), .I (g27768));
INVX1 gate13402(.O (g28583), .I (I37502));
INVX1 gate13403(.O (I37508), .I (g27769));
INVX1 gate13404(.O (g28607), .I (I37508));
INVX1 gate13405(.O (g28608), .I (g27831));
INVX1 gate13406(.O (g28609), .I (g27839));
INVX1 gate13407(.O (g28610), .I (g27843));
INVX1 gate13408(.O (I37514), .I (g27771));
INVX1 gate13409(.O (g28611), .I (I37514));
INVX1 gate13410(.O (g28612), .I (g28046));
INVX1 gate13411(.O (g28616), .I (g27847));
INVX1 gate13412(.O (g28617), .I (g27858));
INVX1 gate13413(.O (g28618), .I (g27861));
INVX1 gate13414(.O (g28619), .I (g28075));
INVX1 gate13415(.O (g28623), .I (g27872));
INVX1 gate13416(.O (g28624), .I (g27879));
INVX1 gate13417(.O (g28625), .I (g28100));
INVX1 gate13418(.O (g28629), .I (g27889));
INVX1 gate13419(.O (g28630), .I (g28118));
INVX1 gate13420(.O (g28638), .I (g28200));
INVX1 gate13421(.O (g28639), .I (g27919));
INVX1 gate13422(.O (g28640), .I (g27928));
INVX1 gate13423(.O (g28641), .I (g27932));
INVX1 gate13424(.O (g28642), .I (g27939));
INVX1 gate13425(.O (g28643), .I (g27942));
INVX1 gate13426(.O (g28644), .I (g27946));
INVX1 gate13427(.O (g28645), .I (g27952));
INVX1 gate13428(.O (g28646), .I (g27956));
INVX1 gate13429(.O (g28647), .I (g27959));
INVX1 gate13430(.O (g28648), .I (g27965));
INVX1 gate13431(.O (g28649), .I (g27973));
INVX1 gate13432(.O (g28650), .I (g27977));
INVX1 gate13433(.O (g28651), .I (g27981));
INVX1 gate13434(.O (g28652), .I (g27994));
INVX1 gate13435(.O (g28653), .I (g27999));
INVX1 gate13436(.O (g28655), .I (g28018));
INVX1 gate13437(.O (I37566), .I (g28370));
INVX1 gate13438(.O (g28673), .I (I37566));
INVX1 gate13439(.O (I37569), .I (g28498));
INVX1 gate13440(.O (g28674), .I (I37569));
INVX1 gate13441(.O (I37572), .I (g28524));
INVX1 gate13442(.O (g28675), .I (I37572));
INVX1 gate13443(.O (I37575), .I (g28527));
INVX1 gate13444(.O (g28676), .I (I37575));
INVX1 gate13445(.O (I37578), .I (g28432));
INVX1 gate13446(.O (g28677), .I (I37578));
INVX1 gate13447(.O (I37581), .I (g28374));
INVX1 gate13448(.O (g28678), .I (I37581));
INVX1 gate13449(.O (I37584), .I (g28526));
INVX1 gate13450(.O (g28679), .I (I37584));
INVX1 gate13451(.O (I37587), .I (g28552));
INVX1 gate13452(.O (g28680), .I (I37587));
INVX1 gate13453(.O (I37590), .I (g28555));
INVX1 gate13454(.O (g28681), .I (I37590));
INVX1 gate13455(.O (I37593), .I (g28443));
INVX1 gate13456(.O (g28682), .I (I37593));
INVX1 gate13457(.O (I37596), .I (g28377));
INVX1 gate13458(.O (g28683), .I (I37596));
INVX1 gate13459(.O (I37599), .I (g28553));
INVX1 gate13460(.O (g28684), .I (I37599));
INVX1 gate13461(.O (I37602), .I (g28579));
INVX1 gate13462(.O (g28685), .I (I37602));
INVX1 gate13463(.O (I37605), .I (g28583));
INVX1 gate13464(.O (g28686), .I (I37605));
INVX1 gate13465(.O (I37608), .I (g28455));
INVX1 gate13466(.O (g28687), .I (I37608));
INVX1 gate13467(.O (I37611), .I (g28382));
INVX1 gate13468(.O (g28688), .I (I37611));
INVX1 gate13469(.O (I37614), .I (g28580));
INVX1 gate13470(.O (g28689), .I (I37614));
INVX1 gate13471(.O (I37617), .I (g28607));
INVX1 gate13472(.O (g28690), .I (I37617));
INVX1 gate13473(.O (I37620), .I (g28611));
INVX1 gate13474(.O (g28691), .I (I37620));
INVX1 gate13475(.O (I37623), .I (g28467));
INVX1 gate13476(.O (g28692), .I (I37623));
INVX1 gate13477(.O (I37626), .I (g28393));
INVX1 gate13478(.O (g28693), .I (I37626));
INVX1 gate13479(.O (I37629), .I (g28369));
INVX1 gate13480(.O (g28694), .I (I37629));
INVX1 gate13481(.O (I37632), .I (g28372));
INVX1 gate13482(.O (g28695), .I (I37632));
INVX1 gate13483(.O (I37635), .I (g28390));
INVX1 gate13484(.O (g28696), .I (I37635));
INVX1 gate13485(.O (I37638), .I (g28395));
INVX1 gate13486(.O (g28697), .I (I37638));
INVX1 gate13487(.O (I37641), .I (g28375));
INVX1 gate13488(.O (g28698), .I (I37641));
INVX1 gate13489(.O (I37644), .I (g28341));
INVX1 gate13490(.O (g28699), .I (I37644));
INVX1 gate13491(.O (I37647), .I (g28343));
INVX1 gate13492(.O (g28700), .I (I37647));
INVX1 gate13493(.O (I37650), .I (g28347));
INVX1 gate13494(.O (g28701), .I (I37650));
INVX1 gate13495(.O (I37653), .I (g28359));
INVX1 gate13496(.O (g28702), .I (I37653));
INVX1 gate13497(.O (I37656), .I (g28365));
INVX1 gate13498(.O (g28703), .I (I37656));
INVX1 gate13499(.O (I37659), .I (g28437));
INVX1 gate13500(.O (g28704), .I (I37659));
INVX1 gate13501(.O (I37662), .I (g28447));
INVX1 gate13502(.O (g28705), .I (I37662));
INVX1 gate13503(.O (I37665), .I (g28458));
INVX1 gate13504(.O (g28706), .I (I37665));
INVX1 gate13505(.O (g28720), .I (g28495));
INVX1 gate13506(.O (g28721), .I (g28490));
INVX1 gate13507(.O (g28723), .I (g28528));
INVX1 gate13508(.O (g28725), .I (g28499));
INVX1 gate13509(.O (g28727), .I (g28489));
INVX1 gate13510(.O (g28730), .I (g28470));
INVX1 gate13511(.O (g28734), .I (g28525));
INVX1 gate13512(.O (g28740), .I (g28488));
INVX1 gate13513(.O (I37702), .I (g28512));
INVX1 gate13514(.O (g28741), .I (I37702));
INVX1 gate13515(.O (I37712), .I (g28512));
INVX1 gate13516(.O (g28751), .I (I37712));
INVX1 gate13517(.O (I37716), .I (g28540));
INVX1 gate13518(.O (g28755), .I (I37716));
INVX1 gate13519(.O (I37725), .I (g28540));
INVX1 gate13520(.O (g28764), .I (I37725));
INVX1 gate13521(.O (I37729), .I (g28567));
INVX1 gate13522(.O (g28768), .I (I37729));
INVX1 gate13523(.O (I37736), .I (g28567));
INVX1 gate13524(.O (g28775), .I (I37736));
INVX1 gate13525(.O (I37740), .I (g28595));
INVX1 gate13526(.O (g28779), .I (I37740));
INVX1 gate13527(.O (I37746), .I (g28595));
INVX1 gate13528(.O (g28785), .I (I37746));
INVX1 gate13529(.O (I37752), .I (g28512));
INVX1 gate13530(.O (g28791), .I (I37752));
INVX1 gate13531(.O (I37757), .I (g28512));
INVX1 gate13532(.O (g28796), .I (I37757));
INVX1 gate13533(.O (I37760), .I (g28540));
INVX1 gate13534(.O (g28799), .I (I37760));
INVX1 gate13535(.O (I37765), .I (g28512));
INVX1 gate13536(.O (g28804), .I (I37765));
INVX1 gate13537(.O (I37768), .I (g28540));
INVX1 gate13538(.O (g28807), .I (I37768));
INVX1 gate13539(.O (I37771), .I (g28567));
INVX1 gate13540(.O (g28810), .I (I37771));
INVX1 gate13541(.O (I37775), .I (g28540));
INVX1 gate13542(.O (g28814), .I (I37775));
INVX1 gate13543(.O (I37778), .I (g28567));
INVX1 gate13544(.O (g28817), .I (I37778));
INVX1 gate13545(.O (I37781), .I (g28595));
INVX1 gate13546(.O (g28820), .I (I37781));
INVX1 gate13547(.O (I37784), .I (g28567));
INVX1 gate13548(.O (g28823), .I (I37784));
INVX1 gate13549(.O (I37787), .I (g28595));
INVX1 gate13550(.O (g28826), .I (I37787));
INVX1 gate13551(.O (I37790), .I (g28595));
INVX1 gate13552(.O (g28829), .I (I37790));
INVX1 gate13553(.O (I37793), .I (g28638));
INVX1 gate13554(.O (g28832), .I (I37793));
INVX1 gate13555(.O (I37796), .I (g28634));
INVX1 gate13556(.O (g28833), .I (I37796));
INVX1 gate13557(.O (I37800), .I (g28635));
INVX1 gate13558(.O (g28835), .I (I37800));
INVX1 gate13559(.O (I37804), .I (g28636));
INVX1 gate13560(.O (g28837), .I (I37804));
INVX1 gate13561(.O (I37808), .I (g28637));
INVX1 gate13562(.O (g28839), .I (I37808));
INVX1 gate13563(.O (g28855), .I (g28409));
INVX1 gate13564(.O (g28859), .I (g28413));
INVX1 gate13565(.O (g28863), .I (g28417));
INVX1 gate13566(.O (g28867), .I (g28418));
INVX1 gate13567(.O (I37842), .I (g28501));
INVX1 gate13568(.O (g28871), .I (I37842));
INVX1 gate13569(.O (I37846), .I (g28501));
INVX1 gate13570(.O (g28877), .I (I37846));
INVX1 gate13571(.O (I37851), .I (g28668));
INVX1 gate13572(.O (g28882), .I (I37851));
INVX1 gate13573(.O (I37854), .I (g28529));
INVX1 gate13574(.O (g28883), .I (I37854));
INVX1 gate13575(.O (I37858), .I (g28501));
INVX1 gate13576(.O (g28889), .I (I37858));
INVX1 gate13577(.O (I37863), .I (g28529));
INVX1 gate13578(.O (g28894), .I (I37863));
INVX1 gate13579(.O (I37868), .I (g28321));
INVX1 gate13580(.O (g28899), .I (I37868));
INVX1 gate13581(.O (I37871), .I (g28556));
INVX1 gate13582(.O (g28900), .I (I37871));
INVX1 gate13583(.O (I37875), .I (g28501));
INVX1 gate13584(.O (g28906), .I (I37875));
INVX1 gate13585(.O (I37880), .I (g28529));
INVX1 gate13586(.O (g28911), .I (I37880));
INVX1 gate13587(.O (I37885), .I (g28556));
INVX1 gate13588(.O (g28916), .I (I37885));
INVX1 gate13589(.O (I37891), .I (g28325));
INVX1 gate13590(.O (g28924), .I (I37891));
INVX1 gate13591(.O (I37894), .I (g28584));
INVX1 gate13592(.O (g28925), .I (I37894));
INVX1 gate13593(.O (I37897), .I (g28501));
INVX1 gate13594(.O (g28928), .I (I37897));
INVX1 gate13595(.O (I37901), .I (g28529));
INVX1 gate13596(.O (g28932), .I (I37901));
INVX1 gate13597(.O (I37906), .I (g28556));
INVX1 gate13598(.O (g28937), .I (I37906));
INVX1 gate13599(.O (I37912), .I (g28584));
INVX1 gate13600(.O (g28945), .I (I37912));
INVX1 gate13601(.O (I37917), .I (g28328));
INVX1 gate13602(.O (g28950), .I (I37917));
INVX1 gate13603(.O (I37920), .I (g28501));
INVX1 gate13604(.O (g28951), .I (I37920));
INVX1 gate13605(.O (I37924), .I (g28529));
INVX1 gate13606(.O (g28955), .I (I37924));
INVX1 gate13607(.O (I37928), .I (g28556));
INVX1 gate13608(.O (g28959), .I (I37928));
INVX1 gate13609(.O (I37934), .I (g28584));
INVX1 gate13610(.O (g28967), .I (I37934));
INVX1 gate13611(.O (I37939), .I (g28501));
INVX1 gate13612(.O (g28972), .I (I37939));
INVX1 gate13613(.O (I37942), .I (g28501));
INVX1 gate13614(.O (g28975), .I (I37942));
INVX1 gate13615(.O (I37946), .I (g28529));
INVX1 gate13616(.O (g28979), .I (I37946));
INVX1 gate13617(.O (I37950), .I (g28556));
INVX1 gate13618(.O (g28983), .I (I37950));
INVX1 gate13619(.O (I37956), .I (g28584));
INVX1 gate13620(.O (g28993), .I (I37956));
INVX1 gate13621(.O (I37961), .I (g28501));
INVX1 gate13622(.O (g28998), .I (I37961));
INVX1 gate13623(.O (I37965), .I (g28529));
INVX1 gate13624(.O (g29002), .I (I37965));
INVX1 gate13625(.O (I37968), .I (g28529));
INVX1 gate13626(.O (g29005), .I (I37968));
INVX1 gate13627(.O (I37973), .I (g28556));
INVX1 gate13628(.O (g29010), .I (I37973));
INVX1 gate13629(.O (I37978), .I (g28584));
INVX1 gate13630(.O (g29019), .I (I37978));
INVX1 gate13631(.O (I37982), .I (g28501));
INVX1 gate13632(.O (g29023), .I (I37982));
INVX1 gate13633(.O (I37986), .I (g28529));
INVX1 gate13634(.O (g29027), .I (I37986));
INVX1 gate13635(.O (I37991), .I (g28556));
INVX1 gate13636(.O (g29032), .I (I37991));
INVX1 gate13637(.O (I37994), .I (g28556));
INVX1 gate13638(.O (g29035), .I (I37994));
INVX1 gate13639(.O (I37999), .I (g28584));
INVX1 gate13640(.O (g29042), .I (I37999));
INVX1 gate13641(.O (I38003), .I (g28529));
INVX1 gate13642(.O (g29046), .I (I38003));
INVX1 gate13643(.O (I38007), .I (g28556));
INVX1 gate13644(.O (g29050), .I (I38007));
INVX1 gate13645(.O (I38011), .I (g28584));
INVX1 gate13646(.O (g29054), .I (I38011));
INVX1 gate13647(.O (I38014), .I (g28584));
INVX1 gate13648(.O (g29057), .I (I38014));
INVX1 gate13649(.O (I38018), .I (g28342));
INVX1 gate13650(.O (g29061), .I (I38018));
INVX1 gate13651(.O (I38024), .I (g28556));
INVX1 gate13652(.O (g29065), .I (I38024));
INVX1 gate13653(.O (I38028), .I (g28584));
INVX1 gate13654(.O (g29069), .I (I38028));
INVX1 gate13655(.O (I38032), .I (g28344));
INVX1 gate13656(.O (g29073), .I (I38032));
INVX1 gate13657(.O (I38035), .I (g28345));
INVX1 gate13658(.O (g29074), .I (I38035));
INVX1 gate13659(.O (I38038), .I (g28346));
INVX1 gate13660(.O (g29075), .I (I38038));
INVX1 gate13661(.O (I38042), .I (g28584));
INVX1 gate13662(.O (g29077), .I (I38042));
INVX1 gate13663(.O (I38046), .I (g28348));
INVX1 gate13664(.O (g29081), .I (I38046));
INVX1 gate13665(.O (I38049), .I (g28349));
INVX1 gate13666(.O (g29082), .I (I38049));
INVX1 gate13667(.O (I38053), .I (g28350));
INVX1 gate13668(.O (g29084), .I (I38053));
INVX1 gate13669(.O (I38056), .I (g28351));
INVX1 gate13670(.O (g29085), .I (I38056));
INVX1 gate13671(.O (I38059), .I (g28352));
INVX1 gate13672(.O (g29086), .I (I38059));
INVX1 gate13673(.O (I38064), .I (g28353));
INVX1 gate13674(.O (g29089), .I (I38064));
INVX1 gate13675(.O (I38068), .I (g28354));
INVX1 gate13676(.O (g29091), .I (I38068));
INVX1 gate13677(.O (I38071), .I (g28355));
INVX1 gate13678(.O (g29092), .I (I38071));
INVX1 gate13679(.O (I38074), .I (g28356));
INVX1 gate13680(.O (g29093), .I (I38074));
INVX1 gate13681(.O (I38077), .I (g28357));
INVX1 gate13682(.O (g29094), .I (I38077));
INVX1 gate13683(.O (I38080), .I (g28358));
INVX1 gate13684(.O (g29095), .I (I38080));
INVX1 gate13685(.O (I38085), .I (g28360));
INVX1 gate13686(.O (g29098), .I (I38085));
INVX1 gate13687(.O (I38088), .I (g28361));
INVX1 gate13688(.O (g29099), .I (I38088));
INVX1 gate13689(.O (I38091), .I (g28362));
INVX1 gate13690(.O (g29100), .I (I38091));
INVX1 gate13691(.O (I38094), .I (g28363));
INVX1 gate13692(.O (g29101), .I (I38094));
INVX1 gate13693(.O (I38097), .I (g28364));
INVX1 gate13694(.O (g29102), .I (I38097));
INVX1 gate13695(.O (I38101), .I (g28366));
INVX1 gate13696(.O (g29104), .I (I38101));
INVX1 gate13697(.O (I38104), .I (g28367));
INVX1 gate13698(.O (g29105), .I (I38104));
INVX1 gate13699(.O (I38107), .I (g28368));
INVX1 gate13700(.O (g29106), .I (I38107));
INVX1 gate13701(.O (I38111), .I (g28371));
INVX1 gate13702(.O (g29108), .I (I38111));
INVX1 gate13703(.O (I38119), .I (g28420));
INVX1 gate13704(.O (g29117), .I (I38119));
INVX1 gate13705(.O (I38122), .I (g28421));
INVX1 gate13706(.O (g29118), .I (I38122));
INVX1 gate13707(.O (I38125), .I (g28425));
INVX1 gate13708(.O (g29119), .I (I38125));
INVX1 gate13709(.O (I38128), .I (g28419));
INVX1 gate13710(.O (g29120), .I (I38128));
INVX1 gate13711(.O (I38136), .I (g28833));
INVX1 gate13712(.O (g29131), .I (I38136));
INVX1 gate13713(.O (I38139), .I (g29061));
INVX1 gate13714(.O (g29132), .I (I38139));
INVX1 gate13715(.O (I38142), .I (g29073));
INVX1 gate13716(.O (g29133), .I (I38142));
INVX1 gate13717(.O (I38145), .I (g29081));
INVX1 gate13718(.O (g29134), .I (I38145));
INVX1 gate13719(.O (I38148), .I (g29074));
INVX1 gate13720(.O (g29135), .I (I38148));
INVX1 gate13721(.O (I38151), .I (g29082));
INVX1 gate13722(.O (g29136), .I (I38151));
INVX1 gate13723(.O (I38154), .I (g29089));
INVX1 gate13724(.O (g29137), .I (I38154));
INVX1 gate13725(.O (I38157), .I (g28882));
INVX1 gate13726(.O (g29138), .I (I38157));
INVX1 gate13727(.O (I38160), .I (g28835));
INVX1 gate13728(.O (g29139), .I (I38160));
INVX1 gate13729(.O (I38163), .I (g29075));
INVX1 gate13730(.O (g29140), .I (I38163));
INVX1 gate13731(.O (I38166), .I (g29084));
INVX1 gate13732(.O (g29141), .I (I38166));
INVX1 gate13733(.O (I38169), .I (g29091));
INVX1 gate13734(.O (g29142), .I (I38169));
INVX1 gate13735(.O (I38172), .I (g29085));
INVX1 gate13736(.O (g29143), .I (I38172));
INVX1 gate13737(.O (I38175), .I (g29092));
INVX1 gate13738(.O (g29144), .I (I38175));
INVX1 gate13739(.O (I38178), .I (g29098));
INVX1 gate13740(.O (g29145), .I (I38178));
INVX1 gate13741(.O (I38181), .I (g28899));
INVX1 gate13742(.O (g29146), .I (I38181));
INVX1 gate13743(.O (I38184), .I (g28837));
INVX1 gate13744(.O (g29147), .I (I38184));
INVX1 gate13745(.O (I38187), .I (g29086));
INVX1 gate13746(.O (g29148), .I (I38187));
INVX1 gate13747(.O (I38190), .I (g29093));
INVX1 gate13748(.O (g29149), .I (I38190));
INVX1 gate13749(.O (I38193), .I (g29099));
INVX1 gate13750(.O (g29150), .I (I38193));
INVX1 gate13751(.O (I38196), .I (g29094));
INVX1 gate13752(.O (g29151), .I (I38196));
INVX1 gate13753(.O (I38199), .I (g29100));
INVX1 gate13754(.O (g29152), .I (I38199));
INVX1 gate13755(.O (I38202), .I (g29104));
INVX1 gate13756(.O (g29153), .I (I38202));
INVX1 gate13757(.O (I38205), .I (g28924));
INVX1 gate13758(.O (g29154), .I (I38205));
INVX1 gate13759(.O (I38208), .I (g28839));
INVX1 gate13760(.O (g29155), .I (I38208));
INVX1 gate13761(.O (I38211), .I (g29095));
INVX1 gate13762(.O (g29156), .I (I38211));
INVX1 gate13763(.O (I38214), .I (g29101));
INVX1 gate13764(.O (g29157), .I (I38214));
INVX1 gate13765(.O (I38217), .I (g29105));
INVX1 gate13766(.O (g29158), .I (I38217));
INVX1 gate13767(.O (I38220), .I (g29102));
INVX1 gate13768(.O (g29159), .I (I38220));
INVX1 gate13769(.O (I38223), .I (g29106));
INVX1 gate13770(.O (g29160), .I (I38223));
INVX1 gate13771(.O (I38226), .I (g29108));
INVX1 gate13772(.O (g29161), .I (I38226));
INVX1 gate13773(.O (I38229), .I (g28950));
INVX1 gate13774(.O (g29162), .I (I38229));
INVX1 gate13775(.O (I38232), .I (g29117));
INVX1 gate13776(.O (g29163), .I (I38232));
INVX1 gate13777(.O (I38235), .I (g29118));
INVX1 gate13778(.O (g29164), .I (I38235));
INVX1 gate13779(.O (I38238), .I (g29119));
INVX1 gate13780(.O (g29165), .I (I38238));
INVX1 gate13781(.O (I38241), .I (g28832));
INVX1 gate13782(.O (g29166), .I (I38241));
INVX1 gate13783(.O (I38245), .I (g28920));
INVX1 gate13784(.O (g29168), .I (I38245));
INVX1 gate13785(.O (I38250), .I (g28941));
INVX1 gate13786(.O (g29171), .I (I38250));
INVX1 gate13787(.O (I38258), .I (g28963));
INVX1 gate13788(.O (g29177), .I (I38258));
INVX1 gate13789(.O (I38272), .I (g29013));
INVX1 gate13790(.O (g29189), .I (I38272));
INVX1 gate13791(.O (I38275), .I (g28987));
INVX1 gate13792(.O (g29190), .I (I38275));
INVX1 gate13793(.O (I38278), .I (g28963));
INVX1 gate13794(.O (g29191), .I (I38278));
INVX1 gate13795(.O (g29192), .I (g28954));
INVX1 gate13796(.O (I38282), .I (g28941));
INVX1 gate13797(.O (g29193), .I (I38282));
INVX1 gate13798(.O (I38321), .I (g29113));
INVX1 gate13799(.O (g29230), .I (I38321));
INVX1 gate13800(.O (I38330), .I (g29120));
INVX1 gate13801(.O (g29237), .I (I38330));
INVX1 gate13802(.O (I38339), .I (g29120));
INVX1 gate13803(.O (g29244), .I (I38339));
INVX1 gate13804(.O (I38342), .I (g28886));
INVX1 gate13805(.O (g29245), .I (I38342));
INVX1 gate13806(.O (I38345), .I (g29109));
INVX1 gate13807(.O (g29246), .I (I38345));
INVX1 gate13808(.O (I38348), .I (g28874));
INVX1 gate13809(.O (g29247), .I (I38348));
INVX1 gate13810(.O (I38352), .I (g29110));
INVX1 gate13811(.O (g29249), .I (I38352));
INVX1 gate13812(.O (I38355), .I (g29039));
INVX1 gate13813(.O (g29250), .I (I38355));
INVX1 gate13814(.O (I38360), .I (g29111));
INVX1 gate13815(.O (g29253), .I (I38360));
INVX1 gate13816(.O (I38363), .I (g29016));
INVX1 gate13817(.O (g29254), .I (I38363));
INVX1 gate13818(.O (I38369), .I (g29112));
INVX1 gate13819(.O (g29258), .I (I38369));
INVX1 gate13820(.O (g29266), .I (g28741));
INVX1 gate13821(.O (I38386), .I (g28734));
INVX1 gate13822(.O (g29267), .I (I38386));
INVX1 gate13823(.O (g29268), .I (g28751));
INVX1 gate13824(.O (g29269), .I (g28755));
INVX1 gate13825(.O (I38391), .I (g28730));
INVX1 gate13826(.O (g29270), .I (I38391));
INVX1 gate13827(.O (g29271), .I (g28764));
INVX1 gate13828(.O (g29272), .I (g28768));
INVX1 gate13829(.O (I38396), .I (g28727));
INVX1 gate13830(.O (g29273), .I (I38396));
INVX1 gate13831(.O (g29274), .I (g28775));
INVX1 gate13832(.O (g29275), .I (g28779));
INVX1 gate13833(.O (I38401), .I (g28725));
INVX1 gate13834(.O (g29276), .I (I38401));
INVX1 gate13835(.O (g29277), .I (g28785));
INVX1 gate13836(.O (I38405), .I (g28723));
INVX1 gate13837(.O (g29278), .I (I38405));
INVX1 gate13838(.O (I38408), .I (g28721));
INVX1 gate13839(.O (g29279), .I (I38408));
INVX1 gate13840(.O (g29280), .I (g28791));
INVX1 gate13841(.O (I38412), .I (g28720));
INVX1 gate13842(.O (g29281), .I (I38412));
INVX1 gate13843(.O (g29282), .I (g28796));
INVX1 gate13844(.O (g29283), .I (g28799));
INVX1 gate13845(.O (g29285), .I (g28804));
INVX1 gate13846(.O (g29286), .I (g28807));
INVX1 gate13847(.O (g29287), .I (g28810));
INVX1 gate13848(.O (I38421), .I (g28740));
INVX1 gate13849(.O (g29288), .I (I38421));
INVX1 gate13850(.O (g29290), .I (g28814));
INVX1 gate13851(.O (g29291), .I (g28817));
INVX1 gate13852(.O (g29292), .I (g28820));
INVX1 gate13853(.O (I38428), .I (g28732));
INVX1 gate13854(.O (g29293), .I (I38428));
INVX1 gate13855(.O (g29295), .I (g28823));
INVX1 gate13856(.O (g29296), .I (g28826));
INVX1 gate13857(.O (I38434), .I (g28735));
INVX1 gate13858(.O (g29297), .I (I38434));
INVX1 gate13859(.O (I38437), .I (g28736));
INVX1 gate13860(.O (g29298), .I (I38437));
INVX1 gate13861(.O (I38440), .I (g28738));
INVX1 gate13862(.O (g29299), .I (I38440));
INVX1 gate13863(.O (g29301), .I (g28829));
INVX1 gate13864(.O (I38447), .I (g28744));
INVX1 gate13865(.O (g29304), .I (I38447));
INVX1 gate13866(.O (I38450), .I (g28745));
INVX1 gate13867(.O (g29305), .I (I38450));
INVX1 gate13868(.O (I38453), .I (g28746));
INVX1 gate13869(.O (g29306), .I (I38453));
INVX1 gate13870(.O (I38456), .I (g28747));
INVX1 gate13871(.O (g29307), .I (I38456));
INVX1 gate13872(.O (I38459), .I (g28749));
INVX1 gate13873(.O (g29308), .I (I38459));
INVX1 gate13874(.O (I38462), .I (g29120));
INVX1 gate13875(.O (g29309), .I (I38462));
INVX1 gate13876(.O (I38466), .I (g28754));
INVX1 gate13877(.O (g29311), .I (I38466));
INVX1 gate13878(.O (I38471), .I (g28758));
INVX1 gate13879(.O (g29314), .I (I38471));
INVX1 gate13880(.O (I38474), .I (g28759));
INVX1 gate13881(.O (g29315), .I (I38474));
INVX1 gate13882(.O (I38477), .I (g28760));
INVX1 gate13883(.O (g29316), .I (I38477));
INVX1 gate13884(.O (I38480), .I (g28761));
INVX1 gate13885(.O (g29317), .I (I38480));
INVX1 gate13886(.O (I38483), .I (g28990));
INVX1 gate13887(.O (g29318), .I (I38483));
INVX1 gate13888(.O (I38486), .I (g28763));
INVX1 gate13889(.O (g29319), .I (I38486));
INVX1 gate13890(.O (I38491), .I (g28767));
INVX1 gate13891(.O (g29322), .I (I38491));
INVX1 gate13892(.O (I38496), .I (g28771));
INVX1 gate13893(.O (g29325), .I (I38496));
INVX1 gate13894(.O (I38499), .I (g28772));
INVX1 gate13895(.O (g29326), .I (I38499));
INVX1 gate13896(.O (I38502), .I (g28773));
INVX1 gate13897(.O (g29327), .I (I38502));
INVX1 gate13898(.O (I38505), .I (g28774));
INVX1 gate13899(.O (g29328), .I (I38505));
INVX1 gate13900(.O (I38510), .I (g28778));
INVX1 gate13901(.O (g29331), .I (I38510));
INVX1 gate13902(.O (I38515), .I (g28782));
INVX1 gate13903(.O (g29334), .I (I38515));
INVX1 gate13904(.O (I38518), .I (g28783));
INVX1 gate13905(.O (g29335), .I (I38518));
INVX1 gate13906(.O (I38524), .I (g28788));
INVX1 gate13907(.O (g29339), .I (I38524));
INVX1 gate13908(.O (I38536), .I (g28920));
INVX1 gate13909(.O (g29349), .I (I38536));
INVX1 gate13910(.O (I38539), .I (g29113));
INVX1 gate13911(.O (g29350), .I (I38539));
INVX1 gate13912(.O (g29356), .I (g29120));
INVX1 gate13913(.O (g29358), .I (g29120));
INVX1 gate13914(.O (I38548), .I (g28903));
INVX1 gate13915(.O (g29359), .I (I38548));
INVX1 gate13916(.O (g29360), .I (g28871));
INVX1 gate13917(.O (g29361), .I (g28877));
INVX1 gate13918(.O (g29362), .I (g28883));
INVX1 gate13919(.O (g29363), .I (g28889));
INVX1 gate13920(.O (g29364), .I (g28894));
INVX1 gate13921(.O (g29365), .I (g28900));
INVX1 gate13922(.O (g29366), .I (g28906));
INVX1 gate13923(.O (g29367), .I (g28911));
INVX1 gate13924(.O (g29368), .I (g28916));
INVX1 gate13925(.O (g29369), .I (g28925));
INVX1 gate13926(.O (g29370), .I (g28928));
INVX1 gate13927(.O (g29371), .I (g28932));
INVX1 gate13928(.O (g29372), .I (g28937));
INVX1 gate13929(.O (g29373), .I (g28945));
INVX1 gate13930(.O (g29374), .I (g28951));
INVX1 gate13931(.O (g29375), .I (g28955));
INVX1 gate13932(.O (g29376), .I (g28959));
INVX1 gate13933(.O (g29377), .I (g28967));
INVX1 gate13934(.O (g29378), .I (g28972));
INVX1 gate13935(.O (g29379), .I (g28975));
INVX1 gate13936(.O (g29380), .I (g28979));
INVX1 gate13937(.O (g29381), .I (g28983));
INVX1 gate13938(.O (g29382), .I (g28993));
INVX1 gate13939(.O (g29383), .I (g28998));
INVX1 gate13940(.O (g29384), .I (g29002));
INVX1 gate13941(.O (g29385), .I (g29005));
INVX1 gate13942(.O (g29386), .I (g29010));
INVX1 gate13943(.O (g29387), .I (g29019));
INVX1 gate13944(.O (g29388), .I (g29023));
INVX1 gate13945(.O (g29389), .I (g29027));
INVX1 gate13946(.O (g29390), .I (g29032));
INVX1 gate13947(.O (g29391), .I (g29035));
INVX1 gate13948(.O (g29392), .I (g29042));
INVX1 gate13949(.O (g29393), .I (g29046));
INVX1 gate13950(.O (g29394), .I (g29050));
INVX1 gate13951(.O (g29395), .I (g29054));
INVX1 gate13952(.O (g29396), .I (g29057));
INVX1 gate13953(.O (g29397), .I (g29065));
INVX1 gate13954(.O (g29398), .I (g29069));
INVX1 gate13955(.O (I38591), .I (g28987));
INVX1 gate13956(.O (g29400), .I (I38591));
INVX1 gate13957(.O (I38594), .I (g28990));
INVX1 gate13958(.O (g29401), .I (I38594));
INVX1 gate13959(.O (g29402), .I (g29077));
INVX1 gate13960(.O (I38599), .I (g29013));
INVX1 gate13961(.O (g29404), .I (I38599));
INVX1 gate13962(.O (I38602), .I (g29016));
INVX1 gate13963(.O (g29405), .I (I38602));
INVX1 gate13964(.O (I38606), .I (g29039));
INVX1 gate13965(.O (g29407), .I (I38606));
INVX1 gate13966(.O (I38609), .I (g28874));
INVX1 gate13967(.O (g29408), .I (I38609));
INVX1 gate13968(.O (I38613), .I (g28886));
INVX1 gate13969(.O (g29410), .I (I38613));
INVX1 gate13970(.O (I38617), .I (g28903));
INVX1 gate13971(.O (g29412), .I (I38617));
INVX1 gate13972(.O (I38620), .I (g29246));
INVX1 gate13973(.O (g29413), .I (I38620));
INVX1 gate13974(.O (I38623), .I (g29293));
INVX1 gate13975(.O (g29414), .I (I38623));
INVX1 gate13976(.O (I38626), .I (g29297));
INVX1 gate13977(.O (g29415), .I (I38626));
INVX1 gate13978(.O (I38629), .I (g29304));
INVX1 gate13979(.O (g29416), .I (I38629));
INVX1 gate13980(.O (I38632), .I (g29298));
INVX1 gate13981(.O (g29417), .I (I38632));
INVX1 gate13982(.O (I38635), .I (g29305));
INVX1 gate13983(.O (g29418), .I (I38635));
INVX1 gate13984(.O (I38638), .I (g29311));
INVX1 gate13985(.O (g29419), .I (I38638));
INVX1 gate13986(.O (I38641), .I (g29249));
INVX1 gate13987(.O (g29420), .I (I38641));
INVX1 gate13988(.O (I38644), .I (g29299));
INVX1 gate13989(.O (g29421), .I (I38644));
INVX1 gate13990(.O (I38647), .I (g29306));
INVX1 gate13991(.O (g29422), .I (I38647));
INVX1 gate13992(.O (I38650), .I (g29314));
INVX1 gate13993(.O (g29423), .I (I38650));
INVX1 gate13994(.O (I38653), .I (g29307));
INVX1 gate13995(.O (g29424), .I (I38653));
INVX1 gate13996(.O (I38656), .I (g29315));
INVX1 gate13997(.O (g29425), .I (I38656));
INVX1 gate13998(.O (I38659), .I (g29322));
INVX1 gate13999(.O (g29426), .I (I38659));
INVX1 gate14000(.O (I38662), .I (g29253));
INVX1 gate14001(.O (g29427), .I (I38662));
INVX1 gate14002(.O (I38665), .I (g29412));
INVX1 gate14003(.O (g29428), .I (I38665));
INVX1 gate14004(.O (I38668), .I (g29168));
INVX1 gate14005(.O (g29429), .I (I38668));
INVX1 gate14006(.O (I38671), .I (g29171));
INVX1 gate14007(.O (g29430), .I (I38671));
INVX1 gate14008(.O (I38674), .I (g29177));
INVX1 gate14009(.O (g29431), .I (I38674));
INVX1 gate14010(.O (I38677), .I (g29400));
INVX1 gate14011(.O (g29432), .I (I38677));
INVX1 gate14012(.O (I38680), .I (g29404));
INVX1 gate14013(.O (g29433), .I (I38680));
INVX1 gate14014(.O (I38683), .I (g29308));
INVX1 gate14015(.O (g29434), .I (I38683));
INVX1 gate14016(.O (I38686), .I (g29316));
INVX1 gate14017(.O (g29435), .I (I38686));
INVX1 gate14018(.O (I38689), .I (g29325));
INVX1 gate14019(.O (g29436), .I (I38689));
INVX1 gate14020(.O (I38692), .I (g29317));
INVX1 gate14021(.O (g29437), .I (I38692));
INVX1 gate14022(.O (I38695), .I (g29326));
INVX1 gate14023(.O (g29438), .I (I38695));
INVX1 gate14024(.O (I38698), .I (g29331));
INVX1 gate14025(.O (g29439), .I (I38698));
INVX1 gate14026(.O (I38701), .I (g29401));
INVX1 gate14027(.O (g29440), .I (I38701));
INVX1 gate14028(.O (I38704), .I (g29405));
INVX1 gate14029(.O (g29441), .I (I38704));
INVX1 gate14030(.O (I38707), .I (g29407));
INVX1 gate14031(.O (g29442), .I (I38707));
INVX1 gate14032(.O (I38710), .I (g29408));
INVX1 gate14033(.O (g29443), .I (I38710));
INVX1 gate14034(.O (I38713), .I (g29410));
INVX1 gate14035(.O (g29444), .I (I38713));
INVX1 gate14036(.O (I38716), .I (g29230));
INVX1 gate14037(.O (g29445), .I (I38716));
INVX1 gate14038(.O (I38719), .I (g29258));
INVX1 gate14039(.O (g29446), .I (I38719));
INVX1 gate14040(.O (I38722), .I (g29319));
INVX1 gate14041(.O (g29447), .I (I38722));
INVX1 gate14042(.O (I38725), .I (g29327));
INVX1 gate14043(.O (g29448), .I (I38725));
INVX1 gate14044(.O (I38728), .I (g29334));
INVX1 gate14045(.O (g29449), .I (I38728));
INVX1 gate14046(.O (I38731), .I (g29328));
INVX1 gate14047(.O (g29450), .I (I38731));
INVX1 gate14048(.O (I38734), .I (g29335));
INVX1 gate14049(.O (g29451), .I (I38734));
INVX1 gate14050(.O (I38737), .I (g29339));
INVX1 gate14051(.O (g29452), .I (I38737));
INVX1 gate14052(.O (I38740), .I (g29288));
INVX1 gate14053(.O (g29453), .I (I38740));
INVX1 gate14054(.O (I38743), .I (g29267));
INVX1 gate14055(.O (g29454), .I (I38743));
INVX1 gate14056(.O (I38746), .I (g29270));
INVX1 gate14057(.O (g29455), .I (I38746));
INVX1 gate14058(.O (I38749), .I (g29273));
INVX1 gate14059(.O (g29456), .I (I38749));
INVX1 gate14060(.O (I38752), .I (g29276));
INVX1 gate14061(.O (g29457), .I (I38752));
INVX1 gate14062(.O (I38755), .I (g29278));
INVX1 gate14063(.O (g29458), .I (I38755));
INVX1 gate14064(.O (I38758), .I (g29279));
INVX1 gate14065(.O (g29459), .I (I38758));
INVX1 gate14066(.O (I38761), .I (g29281));
INVX1 gate14067(.O (g29460), .I (I38761));
INVX1 gate14068(.O (I38764), .I (g29237));
INVX1 gate14069(.O (g29461), .I (I38764));
INVX1 gate14070(.O (I38767), .I (g29244));
INVX1 gate14071(.O (g29462), .I (I38767));
INVX1 gate14072(.O (I38770), .I (g29309));
INVX1 gate14073(.O (g29463), .I (I38770));
INVX1 gate14074(.O (g29491), .I (g29350));
INVX1 gate14075(.O (I38801), .I (g29358));
INVX1 gate14076(.O (g29495), .I (I38801));
INVX1 gate14077(.O (I38804), .I (g29353));
INVX1 gate14078(.O (g29496), .I (I38804));
INVX1 gate14079(.O (I38807), .I (g29356));
INVX1 gate14080(.O (g29497), .I (I38807));
INVX1 gate14081(.O (I38817), .I (g29354));
INVX1 gate14082(.O (g29499), .I (I38817));
INVX1 gate14083(.O (I38827), .I (g29355));
INVX1 gate14084(.O (g29501), .I (I38827));
INVX1 gate14085(.O (I38838), .I (g29357));
INVX1 gate14086(.O (g29504), .I (I38838));
INVX1 gate14087(.O (I38848), .I (g29167));
INVX1 gate14088(.O (g29506), .I (I38848));
INVX1 gate14089(.O (I38851), .I (g29169));
INVX1 gate14090(.O (g29507), .I (I38851));
INVX1 gate14091(.O (I38854), .I (g29170));
INVX1 gate14092(.O (g29508), .I (I38854));
INVX1 gate14093(.O (I38857), .I (g29172));
INVX1 gate14094(.O (g29509), .I (I38857));
INVX1 gate14095(.O (I38860), .I (g29173));
INVX1 gate14096(.O (g29510), .I (I38860));
INVX1 gate14097(.O (I38863), .I (g29178));
INVX1 gate14098(.O (g29511), .I (I38863));
INVX1 gate14099(.O (I38866), .I (g29179));
INVX1 gate14100(.O (g29512), .I (I38866));
INVX1 gate14101(.O (I38869), .I (g29181));
INVX1 gate14102(.O (g29513), .I (I38869));
INVX1 gate14103(.O (I38872), .I (g29182));
INVX1 gate14104(.O (g29514), .I (I38872));
INVX1 gate14105(.O (I38875), .I (g29184));
INVX1 gate14106(.O (g29515), .I (I38875));
INVX1 gate14107(.O (I38878), .I (g29185));
INVX1 gate14108(.O (g29516), .I (I38878));
INVX1 gate14109(.O (I38881), .I (g29187));
INVX1 gate14110(.O (g29517), .I (I38881));
INVX1 gate14111(.O (I38885), .I (g29192));
INVX1 gate14112(.O (g29519), .I (I38885));
INVX1 gate14113(.O (I38898), .I (g29194));
INVX1 gate14114(.O (g29530), .I (I38898));
INVX1 gate14115(.O (I38905), .I (g29197));
INVX1 gate14116(.O (g29535), .I (I38905));
INVX1 gate14117(.O (I38909), .I (g29198));
INVX1 gate14118(.O (g29537), .I (I38909));
INVX1 gate14119(.O (I38916), .I (g29201));
INVX1 gate14120(.O (g29542), .I (I38916));
INVX1 gate14121(.O (I38920), .I (g29204));
INVX1 gate14122(.O (g29544), .I (I38920));
INVX1 gate14123(.O (I38924), .I (g29205));
INVX1 gate14124(.O (g29546), .I (I38924));
INVX1 gate14125(.O (I38931), .I (g29209));
INVX1 gate14126(.O (g29551), .I (I38931));
INVX1 gate14127(.O (I38936), .I (g29212));
INVX1 gate14128(.O (g29554), .I (I38936));
INVX1 gate14129(.O (I38940), .I (g29213));
INVX1 gate14130(.O (g29556), .I (I38940));
INVX1 gate14131(.O (I38947), .I (g29218));
INVX1 gate14132(.O (g29561), .I (I38947));
INVX1 gate14133(.O (I38951), .I (g29221));
INVX1 gate14134(.O (g29563), .I (I38951));
INVX1 gate14135(.O (I38958), .I (g29226));
INVX1 gate14136(.O (g29568), .I (I38958));
INVX1 gate14137(.O (I38975), .I (g29348));
INVX1 gate14138(.O (g29583), .I (I38975));
INVX1 gate14139(.O (I38999), .I (g29496));
INVX1 gate14140(.O (g29627), .I (I38999));
INVX1 gate14141(.O (I39002), .I (g29506));
INVX1 gate14142(.O (g29628), .I (I39002));
INVX1 gate14143(.O (I39005), .I (g29507));
INVX1 gate14144(.O (g29629), .I (I39005));
INVX1 gate14145(.O (I39008), .I (g29509));
INVX1 gate14146(.O (g29630), .I (I39008));
INVX1 gate14147(.O (I39011), .I (g29530));
INVX1 gate14148(.O (g29631), .I (I39011));
INVX1 gate14149(.O (I39014), .I (g29535));
INVX1 gate14150(.O (g29632), .I (I39014));
INVX1 gate14151(.O (I39017), .I (g29542));
INVX1 gate14152(.O (g29633), .I (I39017));
INVX1 gate14153(.O (I39020), .I (g29499));
INVX1 gate14154(.O (g29634), .I (I39020));
INVX1 gate14155(.O (I39023), .I (g29508));
INVX1 gate14156(.O (g29635), .I (I39023));
INVX1 gate14157(.O (I39026), .I (g29510));
INVX1 gate14158(.O (g29636), .I (I39026));
INVX1 gate14159(.O (I39029), .I (g29512));
INVX1 gate14160(.O (g29637), .I (I39029));
INVX1 gate14161(.O (I39032), .I (g29537));
INVX1 gate14162(.O (g29638), .I (I39032));
INVX1 gate14163(.O (I39035), .I (g29544));
INVX1 gate14164(.O (g29639), .I (I39035));
INVX1 gate14165(.O (I39038), .I (g29551));
INVX1 gate14166(.O (g29640), .I (I39038));
INVX1 gate14167(.O (I39041), .I (g29501));
INVX1 gate14168(.O (g29641), .I (I39041));
INVX1 gate14169(.O (I39044), .I (g29511));
INVX1 gate14170(.O (g29642), .I (I39044));
INVX1 gate14171(.O (I39047), .I (g29513));
INVX1 gate14172(.O (g29643), .I (I39047));
INVX1 gate14173(.O (I39050), .I (g29515));
INVX1 gate14174(.O (g29644), .I (I39050));
INVX1 gate14175(.O (I39053), .I (g29546));
INVX1 gate14176(.O (g29645), .I (I39053));
INVX1 gate14177(.O (I39056), .I (g29554));
INVX1 gate14178(.O (g29646), .I (I39056));
INVX1 gate14179(.O (I39059), .I (g29561));
INVX1 gate14180(.O (g29647), .I (I39059));
INVX1 gate14181(.O (I39062), .I (g29504));
INVX1 gate14182(.O (g29648), .I (I39062));
INVX1 gate14183(.O (I39065), .I (g29514));
INVX1 gate14184(.O (g29649), .I (I39065));
INVX1 gate14185(.O (I39068), .I (g29516));
INVX1 gate14186(.O (g29650), .I (I39068));
INVX1 gate14187(.O (I39071), .I (g29517));
INVX1 gate14188(.O (g29651), .I (I39071));
INVX1 gate14189(.O (I39074), .I (g29556));
INVX1 gate14190(.O (g29652), .I (I39074));
INVX1 gate14191(.O (I39077), .I (g29563));
INVX1 gate14192(.O (g29653), .I (I39077));
INVX1 gate14193(.O (I39080), .I (g29568));
INVX1 gate14194(.O (g29654), .I (I39080));
INVX1 gate14195(.O (I39083), .I (g29519));
INVX1 gate14196(.O (g29655), .I (I39083));
INVX1 gate14197(.O (I39086), .I (g29497));
INVX1 gate14198(.O (g29656), .I (I39086));
INVX1 gate14199(.O (I39089), .I (g29495));
INVX1 gate14200(.O (g29657), .I (I39089));
INVX1 gate14201(.O (g29658), .I (g29574));
INVX1 gate14202(.O (g29659), .I (g29571));
INVX1 gate14203(.O (g29660), .I (g29578));
INVX1 gate14204(.O (g29661), .I (g29576));
INVX1 gate14205(.O (g29662), .I (g29570));
INVX1 gate14206(.O (g29664), .I (g29552));
INVX1 gate14207(.O (g29666), .I (g29577));
INVX1 gate14208(.O (g29668), .I (g29569));
INVX1 gate14209(.O (g29673), .I (g29583));
INVX1 gate14210(.O (I39121), .I (g29579));
INVX1 gate14211(.O (g29689), .I (I39121));
INVX1 gate14212(.O (I39124), .I (g29606));
INVX1 gate14213(.O (g29690), .I (I39124));
INVX1 gate14214(.O (I39127), .I (g29608));
INVX1 gate14215(.O (g29691), .I (I39127));
INVX1 gate14216(.O (I39130), .I (g29580));
INVX1 gate14217(.O (g29692), .I (I39130));
INVX1 gate14218(.O (I39133), .I (g29609));
INVX1 gate14219(.O (g29693), .I (I39133));
INVX1 gate14220(.O (I39136), .I (g29611));
INVX1 gate14221(.O (g29694), .I (I39136));
INVX1 gate14222(.O (I39139), .I (g29612));
INVX1 gate14223(.O (g29695), .I (I39139));
INVX1 gate14224(.O (I39142), .I (g29581));
INVX1 gate14225(.O (g29696), .I (I39142));
INVX1 gate14226(.O (I39145), .I (g29613));
INVX1 gate14227(.O (g29697), .I (I39145));
INVX1 gate14228(.O (I39148), .I (g29616));
INVX1 gate14229(.O (g29698), .I (I39148));
INVX1 gate14230(.O (I39151), .I (g29617));
INVX1 gate14231(.O (g29699), .I (I39151));
INVX1 gate14232(.O (I39154), .I (g29582));
INVX1 gate14233(.O (g29700), .I (I39154));
INVX1 gate14234(.O (I39157), .I (g29618));
INVX1 gate14235(.O (g29701), .I (I39157));
INVX1 gate14236(.O (I39160), .I (g29620));
INVX1 gate14237(.O (g29702), .I (I39160));
INVX1 gate14238(.O (I39164), .I (g29621));
INVX1 gate14239(.O (g29704), .I (I39164));
INVX1 gate14240(.O (I39168), .I (g29623));
INVX1 gate14241(.O (g29708), .I (I39168));
INVX1 gate14242(.O (g29716), .I (g29498));
INVX1 gate14243(.O (g29724), .I (g29500));
INVX1 gate14244(.O (g29726), .I (g29503));
INVX1 gate14245(.O (g29739), .I (g29505));
INVX1 gate14246(.O (I39234), .I (g29689));
INVX1 gate14247(.O (g29794), .I (I39234));
INVX1 gate14248(.O (I39237), .I (g29690));
INVX1 gate14249(.O (g29795), .I (I39237));
INVX1 gate14250(.O (I39240), .I (g29691));
INVX1 gate14251(.O (g29796), .I (I39240));
INVX1 gate14252(.O (I39243), .I (g29694));
INVX1 gate14253(.O (g29797), .I (I39243));
INVX1 gate14254(.O (I39246), .I (g29692));
INVX1 gate14255(.O (g29798), .I (I39246));
INVX1 gate14256(.O (I39249), .I (g29693));
INVX1 gate14257(.O (g29799), .I (I39249));
INVX1 gate14258(.O (I39252), .I (g29695));
INVX1 gate14259(.O (g29800), .I (I39252));
INVX1 gate14260(.O (I39255), .I (g29698));
INVX1 gate14261(.O (g29801), .I (I39255));
INVX1 gate14262(.O (I39258), .I (g29696));
INVX1 gate14263(.O (g29802), .I (I39258));
INVX1 gate14264(.O (I39261), .I (g29697));
INVX1 gate14265(.O (g29803), .I (I39261));
INVX1 gate14266(.O (I39264), .I (g29699));
INVX1 gate14267(.O (g29804), .I (I39264));
INVX1 gate14268(.O (I39267), .I (g29702));
INVX1 gate14269(.O (g29805), .I (I39267));
INVX1 gate14270(.O (I39270), .I (g29700));
INVX1 gate14271(.O (g29806), .I (I39270));
INVX1 gate14272(.O (I39273), .I (g29701));
INVX1 gate14273(.O (g29807), .I (I39273));
INVX1 gate14274(.O (I39276), .I (g29704));
INVX1 gate14275(.O (g29808), .I (I39276));
INVX1 gate14276(.O (I39279), .I (g29708));
INVX1 gate14277(.O (g29809), .I (I39279));
INVX1 gate14278(.O (g29823), .I (g29663));
INVX1 gate14279(.O (g29829), .I (g29665));
INVX1 gate14280(.O (g29835), .I (g29667));
INVX1 gate14281(.O (g29840), .I (g29669));
INVX1 gate14282(.O (g29844), .I (g29670));
INVX1 gate14283(.O (g29848), .I (g29761));
INVX1 gate14284(.O (g29849), .I (g29671));
INVX1 gate14285(.O (g29853), .I (g29672));
INVX1 gate14286(.O (g29857), .I (g29676));
INVX1 gate14287(.O (g29861), .I (g29677));
INVX1 gate14288(.O (g29865), .I (g29678));
INVX1 gate14289(.O (g29869), .I (g29679));
INVX1 gate14290(.O (g29873), .I (g29680));
INVX1 gate14291(.O (g29877), .I (g29681));
INVX1 gate14292(.O (g29881), .I (g29682));
INVX1 gate14293(.O (g29885), .I (g29683));
INVX1 gate14294(.O (g29889), .I (g29684));
INVX1 gate14295(.O (g29893), .I (g29685));
INVX1 gate14296(.O (g29897), .I (g29686));
INVX1 gate14297(.O (g29901), .I (g29687));
INVX1 gate14298(.O (g29905), .I (g29688));
INVX1 gate14299(.O (I39398), .I (g29664));
INVX1 gate14300(.O (g29932), .I (I39398));
INVX1 gate14301(.O (I39401), .I (g29662));
INVX1 gate14302(.O (g29933), .I (I39401));
INVX1 gate14303(.O (I39404), .I (g29661));
INVX1 gate14304(.O (g29934), .I (I39404));
INVX1 gate14305(.O (I39407), .I (g29660));
INVX1 gate14306(.O (g29935), .I (I39407));
INVX1 gate14307(.O (I39411), .I (g29659));
INVX1 gate14308(.O (g29937), .I (I39411));
INVX1 gate14309(.O (I39414), .I (g29658));
INVX1 gate14310(.O (g29938), .I (I39414));
INVX1 gate14311(.O (I39418), .I (g29668));
INVX1 gate14312(.O (g29940), .I (I39418));
INVX1 gate14313(.O (I39423), .I (g29666));
INVX1 gate14314(.O (g29943), .I (I39423));
INVX1 gate14315(.O (I39454), .I (g29940));
INVX1 gate14316(.O (g29972), .I (I39454));
INVX1 gate14317(.O (I39457), .I (g29943));
INVX1 gate14318(.O (g29973), .I (I39457));
INVX1 gate14319(.O (I39460), .I (g29932));
INVX1 gate14320(.O (g29974), .I (I39460));
INVX1 gate14321(.O (I39463), .I (g29933));
INVX1 gate14322(.O (g29975), .I (I39463));
INVX1 gate14323(.O (I39466), .I (g29934));
INVX1 gate14324(.O (g29976), .I (I39466));
INVX1 gate14325(.O (I39469), .I (g29935));
INVX1 gate14326(.O (g29977), .I (I39469));
INVX1 gate14327(.O (I39472), .I (g29937));
INVX1 gate14328(.O (g29978), .I (I39472));
INVX1 gate14329(.O (I39475), .I (g29938));
INVX1 gate14330(.O (g29979), .I (I39475));
INVX1 gate14331(.O (g30036), .I (g29912));
INVX1 gate14332(.O (g30040), .I (g29914));
INVX1 gate14333(.O (g30044), .I (g29916));
INVX1 gate14334(.O (g30048), .I (g29920));
INVX1 gate14335(.O (I39550), .I (g29848));
INVX1 gate14336(.O (g30052), .I (I39550));
INVX1 gate14337(.O (I39573), .I (g29936));
INVX1 gate14338(.O (g30076), .I (I39573));
INVX1 gate14339(.O (I39577), .I (g29939));
INVX1 gate14340(.O (g30078), .I (I39577));
INVX1 gate14341(.O (I39585), .I (g29941));
INVX1 gate14342(.O (g30084), .I (I39585));
INVX1 gate14343(.O (I39622), .I (g30052));
INVX1 gate14344(.O (g30119), .I (I39622));
INVX1 gate14345(.O (I39625), .I (g30076));
INVX1 gate14346(.O (g30120), .I (I39625));
INVX1 gate14347(.O (I39628), .I (g30078));
INVX1 gate14348(.O (g30121), .I (I39628));
INVX1 gate14349(.O (I39631), .I (g30084));
INVX1 gate14350(.O (g30122), .I (I39631));
INVX1 gate14351(.O (I39635), .I (g30055));
INVX1 gate14352(.O (g30124), .I (I39635));
INVX1 gate14353(.O (I39638), .I (g30056));
INVX1 gate14354(.O (g30125), .I (I39638));
INVX1 gate14355(.O (I39641), .I (g30057));
INVX1 gate14356(.O (g30126), .I (I39641));
INVX1 gate14357(.O (I39647), .I (g30058));
INVX1 gate14358(.O (g30130), .I (I39647));
INVX1 gate14359(.O (g30134), .I (g30010));
INVX1 gate14360(.O (g30139), .I (g30011));
INVX1 gate14361(.O (g30143), .I (g30012));
INVX1 gate14362(.O (g30147), .I (g30013));
INVX1 gate14363(.O (g30151), .I (g30014));
INVX1 gate14364(.O (g30155), .I (g30015));
INVX1 gate14365(.O (g30159), .I (g30016));
INVX1 gate14366(.O (g30163), .I (g30017));
INVX1 gate14367(.O (g30167), .I (g30018));
INVX1 gate14368(.O (g30171), .I (g30019));
INVX1 gate14369(.O (g30175), .I (g30020));
INVX1 gate14370(.O (g30179), .I (g30021));
INVX1 gate14371(.O (g30183), .I (g30022));
INVX1 gate14372(.O (g30187), .I (g30023));
INVX1 gate14373(.O (g30191), .I (g30024));
INVX1 gate14374(.O (g30195), .I (g30025));
INVX1 gate14375(.O (g30199), .I (g30026));
INVX1 gate14376(.O (g30203), .I (g30027));
INVX1 gate14377(.O (g30207), .I (g30028));
INVX1 gate14378(.O (g30211), .I (g30029));
INVX1 gate14379(.O (I39674), .I (g30072));
INVX1 gate14380(.O (g30215), .I (I39674));
INVX1 gate14381(.O (g30229), .I (g30030));
INVX1 gate14382(.O (g30233), .I (g30031));
INVX1 gate14383(.O (g30237), .I (g30032));
INVX1 gate14384(.O (g30241), .I (g30033));
INVX1 gate14385(.O (I39761), .I (g30072));
INVX1 gate14386(.O (g30306), .I (I39761));
INVX1 gate14387(.O (I39764), .I (g30060));
INVX1 gate14388(.O (g30307), .I (I39764));
INVX1 gate14389(.O (I39767), .I (g30061));
INVX1 gate14390(.O (g30308), .I (I39767));
INVX1 gate14391(.O (I39770), .I (g30063));
INVX1 gate14392(.O (g30309), .I (I39770));
INVX1 gate14393(.O (I39773), .I (g30064));
INVX1 gate14394(.O (g30310), .I (I39773));
INVX1 gate14395(.O (I39776), .I (g30066));
INVX1 gate14396(.O (g30311), .I (I39776));
INVX1 gate14397(.O (I39779), .I (g30053));
INVX1 gate14398(.O (g30312), .I (I39779));
INVX1 gate14399(.O (I39782), .I (g30054));
INVX1 gate14400(.O (g30313), .I (I39782));
INVX1 gate14401(.O (I39785), .I (g30124));
INVX1 gate14402(.O (g30314), .I (I39785));
INVX1 gate14403(.O (I39788), .I (g30125));
INVX1 gate14404(.O (g30315), .I (I39788));
INVX1 gate14405(.O (I39791), .I (g30126));
INVX1 gate14406(.O (g30316), .I (I39791));
INVX1 gate14407(.O (I39794), .I (g30130));
INVX1 gate14408(.O (g30317), .I (I39794));
INVX1 gate14409(.O (I39797), .I (g30307));
INVX1 gate14410(.O (g30318), .I (I39797));
INVX1 gate14411(.O (I39800), .I (g30309));
INVX1 gate14412(.O (g30319), .I (I39800));
INVX1 gate14413(.O (I39803), .I (g30308));
INVX1 gate14414(.O (g30320), .I (I39803));
INVX1 gate14415(.O (I39806), .I (g30310));
INVX1 gate14416(.O (g30321), .I (I39806));
INVX1 gate14417(.O (I39809), .I (g30311));
INVX1 gate14418(.O (g30322), .I (I39809));
INVX1 gate14419(.O (I39812), .I (g30312));
INVX1 gate14420(.O (g30323), .I (I39812));
INVX1 gate14421(.O (I39815), .I (g30313));
INVX1 gate14422(.O (g30324), .I (I39815));
INVX1 gate14423(.O (I39818), .I (g30215));
INVX1 gate14424(.O (g30325), .I (I39818));
INVX1 gate14425(.O (I39821), .I (g30267));
INVX1 gate14426(.O (g30326), .I (I39821));
INVX1 gate14427(.O (I39825), .I (g30268));
INVX1 gate14428(.O (g30328), .I (I39825));
INVX1 gate14429(.O (I39828), .I (g30269));
INVX1 gate14430(.O (g30329), .I (I39828));
INVX1 gate14431(.O (I39832), .I (g30270));
INVX1 gate14432(.O (g30331), .I (I39832));
INVX1 gate14433(.O (I39835), .I (g30271));
INVX1 gate14434(.O (g30332), .I (I39835));
INVX1 gate14435(.O (I39840), .I (g30272));
INVX1 gate14436(.O (g30335), .I (I39840));
INVX1 gate14437(.O (I39843), .I (g30273));
INVX1 gate14438(.O (g30336), .I (I39843));
INVX1 gate14439(.O (I39848), .I (g30274));
INVX1 gate14440(.O (g30339), .I (I39848));
INVX1 gate14441(.O (I39853), .I (g30275));
INVX1 gate14442(.O (g30342), .I (I39853));
INVX1 gate14443(.O (I39856), .I (g30276));
INVX1 gate14444(.O (g30343), .I (I39856));
INVX1 gate14445(.O (I39859), .I (g30277));
INVX1 gate14446(.O (g30344), .I (I39859));
INVX1 gate14447(.O (I39863), .I (g30278));
INVX1 gate14448(.O (g30346), .I (I39863));
INVX1 gate14449(.O (I39866), .I (g30279));
INVX1 gate14450(.O (g30347), .I (I39866));
INVX1 gate14451(.O (I39870), .I (g30280));
INVX1 gate14452(.O (g30349), .I (I39870));
INVX1 gate14453(.O (I39873), .I (g30281));
INVX1 gate14454(.O (g30350), .I (I39873));
INVX1 gate14455(.O (I39878), .I (g30282));
INVX1 gate14456(.O (g30353), .I (I39878));
INVX1 gate14457(.O (I39881), .I (g30283));
INVX1 gate14458(.O (g30354), .I (I39881));
INVX1 gate14459(.O (I39886), .I (g30284));
INVX1 gate14460(.O (g30357), .I (I39886));
INVX1 gate14461(.O (I39889), .I (g30285));
INVX1 gate14462(.O (g30358), .I (I39889));
INVX1 gate14463(.O (I39892), .I (g30286));
INVX1 gate14464(.O (g30359), .I (I39892));
INVX1 gate14465(.O (I39895), .I (g30287));
INVX1 gate14466(.O (g30360), .I (I39895));
INVX1 gate14467(.O (I39899), .I (g30288));
INVX1 gate14468(.O (g30362), .I (I39899));
INVX1 gate14469(.O (I39902), .I (g30289));
INVX1 gate14470(.O (g30363), .I (I39902));
INVX1 gate14471(.O (I39906), .I (g30290));
INVX1 gate14472(.O (g30365), .I (I39906));
INVX1 gate14473(.O (I39909), .I (g30291));
INVX1 gate14474(.O (g30366), .I (I39909));
INVX1 gate14475(.O (I39913), .I (g30292));
INVX1 gate14476(.O (g30368), .I (I39913));
INVX1 gate14477(.O (I39916), .I (g30293));
INVX1 gate14478(.O (g30369), .I (I39916));
INVX1 gate14479(.O (I39919), .I (g30294));
INVX1 gate14480(.O (g30370), .I (I39919));
INVX1 gate14481(.O (I39922), .I (g30295));
INVX1 gate14482(.O (g30371), .I (I39922));
INVX1 gate14483(.O (I39926), .I (g30296));
INVX1 gate14484(.O (g30373), .I (I39926));
INVX1 gate14485(.O (I39930), .I (g30297));
INVX1 gate14486(.O (g30375), .I (I39930));
INVX1 gate14487(.O (I39933), .I (g30298));
INVX1 gate14488(.O (g30376), .I (I39933));
INVX1 gate14489(.O (I39936), .I (g30299));
INVX1 gate14490(.O (g30377), .I (I39936));
INVX1 gate14491(.O (I39939), .I (g30300));
INVX1 gate14492(.O (g30378), .I (I39939));
INVX1 gate14493(.O (I39942), .I (g30301));
INVX1 gate14494(.O (g30379), .I (I39942));
INVX1 gate14495(.O (I39945), .I (g30302));
INVX1 gate14496(.O (g30380), .I (I39945));
INVX1 gate14497(.O (I39948), .I (g30303));
INVX1 gate14498(.O (g30381), .I (I39948));
INVX1 gate14499(.O (I39951), .I (g30304));
INVX1 gate14500(.O (g30382), .I (I39951));
INVX1 gate14501(.O (g30383), .I (g30306));
INVX1 gate14502(.O (I39976), .I (g30245));
INVX1 gate14503(.O (g30408), .I (I39976));
INVX1 gate14504(.O (I39982), .I (g30305));
INVX1 gate14505(.O (g30412), .I (I39982));
INVX1 gate14506(.O (I39985), .I (g30246));
INVX1 gate14507(.O (g30435), .I (I39985));
INVX1 gate14508(.O (I39991), .I (g30247));
INVX1 gate14509(.O (g30439), .I (I39991));
INVX1 gate14510(.O (I39997), .I (g30248));
INVX1 gate14511(.O (g30443), .I (I39997));
INVX1 gate14512(.O (I40002), .I (g30249));
INVX1 gate14513(.O (g30446), .I (I40002));
INVX1 gate14514(.O (I40008), .I (g30250));
INVX1 gate14515(.O (g30450), .I (I40008));
INVX1 gate14516(.O (I40016), .I (g30251));
INVX1 gate14517(.O (g30456), .I (I40016));
INVX1 gate14518(.O (I40021), .I (g30252));
INVX1 gate14519(.O (g30459), .I (I40021));
INVX1 gate14520(.O (I40027), .I (g30253));
INVX1 gate14521(.O (g30463), .I (I40027));
INVX1 gate14522(.O (I40032), .I (g30254));
INVX1 gate14523(.O (g30466), .I (I40032));
INVX1 gate14524(.O (I40039), .I (g30255));
INVX1 gate14525(.O (g30471), .I (I40039));
INVX1 gate14526(.O (I40044), .I (g30256));
INVX1 gate14527(.O (g30474), .I (I40044));
INVX1 gate14528(.O (I40051), .I (g30257));
INVX1 gate14529(.O (g30479), .I (I40051));
INVX1 gate14530(.O (I40054), .I (g30258));
INVX1 gate14531(.O (g30480), .I (I40054));
INVX1 gate14532(.O (I40059), .I (g30259));
INVX1 gate14533(.O (g30483), .I (I40059));
INVX1 gate14534(.O (I40066), .I (g30260));
INVX1 gate14535(.O (g30488), .I (I40066));
INVX1 gate14536(.O (I40071), .I (g30261));
INVX1 gate14537(.O (g30491), .I (I40071));
INVX1 gate14538(.O (I40075), .I (g30262));
INVX1 gate14539(.O (g30493), .I (I40075));
INVX1 gate14540(.O (I40078), .I (g30263));
INVX1 gate14541(.O (g30494), .I (I40078));
INVX1 gate14542(.O (I40083), .I (g30264));
INVX1 gate14543(.O (g30497), .I (I40083));
INVX1 gate14544(.O (I40086), .I (g30265));
INVX1 gate14545(.O (g30498), .I (I40086));
INVX1 gate14546(.O (I40091), .I (g30266));
INVX1 gate14547(.O (g30501), .I (I40091));
INVX1 gate14548(.O (I40098), .I (g30491));
INVX1 gate14549(.O (g30506), .I (I40098));
INVX1 gate14550(.O (I40101), .I (g30326));
INVX1 gate14551(.O (g30507), .I (I40101));
INVX1 gate14552(.O (I40104), .I (g30342));
INVX1 gate14553(.O (g30508), .I (I40104));
INVX1 gate14554(.O (I40107), .I (g30343));
INVX1 gate14555(.O (g30509), .I (I40107));
INVX1 gate14556(.O (I40110), .I (g30357));
INVX1 gate14557(.O (g30510), .I (I40110));
INVX1 gate14558(.O (I40113), .I (g30368));
INVX1 gate14559(.O (g30511), .I (I40113));
INVX1 gate14560(.O (I40116), .I (g30408));
INVX1 gate14561(.O (g30512), .I (I40116));
INVX1 gate14562(.O (I40119), .I (g30435));
INVX1 gate14563(.O (g30513), .I (I40119));
INVX1 gate14564(.O (I40122), .I (g30443));
INVX1 gate14565(.O (g30514), .I (I40122));
INVX1 gate14566(.O (I40125), .I (g30466));
INVX1 gate14567(.O (g30515), .I (I40125));
INVX1 gate14568(.O (I40128), .I (g30479));
INVX1 gate14569(.O (g30516), .I (I40128));
INVX1 gate14570(.O (I40131), .I (g30493));
INVX1 gate14571(.O (g30517), .I (I40131));
INVX1 gate14572(.O (I40134), .I (g30480));
INVX1 gate14573(.O (g30518), .I (I40134));
INVX1 gate14574(.O (I40137), .I (g30494));
INVX1 gate14575(.O (g30519), .I (I40137));
INVX1 gate14576(.O (I40140), .I (g30328));
INVX1 gate14577(.O (g30520), .I (I40140));
INVX1 gate14578(.O (I40143), .I (g30329));
INVX1 gate14579(.O (g30521), .I (I40143));
INVX1 gate14580(.O (I40146), .I (g30344));
INVX1 gate14581(.O (g30522), .I (I40146));
INVX1 gate14582(.O (I40149), .I (g30358));
INVX1 gate14583(.O (g30523), .I (I40149));
INVX1 gate14584(.O (I40152), .I (g30359));
INVX1 gate14585(.O (g30524), .I (I40152));
INVX1 gate14586(.O (I40155), .I (g30369));
INVX1 gate14587(.O (g30525), .I (I40155));
INVX1 gate14588(.O (I40158), .I (g30376));
INVX1 gate14589(.O (g30526), .I (I40158));
INVX1 gate14590(.O (I40161), .I (g30439));
INVX1 gate14591(.O (g30527), .I (I40161));
INVX1 gate14592(.O (I40164), .I (g30446));
INVX1 gate14593(.O (g30528), .I (I40164));
INVX1 gate14594(.O (I40167), .I (g30456));
INVX1 gate14595(.O (g30529), .I (I40167));
INVX1 gate14596(.O (I40170), .I (g30483));
INVX1 gate14597(.O (g30530), .I (I40170));
INVX1 gate14598(.O (I40173), .I (g30497));
INVX1 gate14599(.O (g30531), .I (I40173));
INVX1 gate14600(.O (I40176), .I (g30331));
INVX1 gate14601(.O (g30532), .I (I40176));
INVX1 gate14602(.O (I40179), .I (g30498));
INVX1 gate14603(.O (g30533), .I (I40179));
INVX1 gate14604(.O (I40182), .I (g30332));
INVX1 gate14605(.O (g30534), .I (I40182));
INVX1 gate14606(.O (I40185), .I (g30346));
INVX1 gate14607(.O (g30535), .I (I40185));
INVX1 gate14608(.O (I40188), .I (g30347));
INVX1 gate14609(.O (g30536), .I (I40188));
INVX1 gate14610(.O (I40191), .I (g30360));
INVX1 gate14611(.O (g30537), .I (I40191));
INVX1 gate14612(.O (I40194), .I (g30370));
INVX1 gate14613(.O (g30538), .I (I40194));
INVX1 gate14614(.O (I40197), .I (g30371));
INVX1 gate14615(.O (g30539), .I (I40197));
INVX1 gate14616(.O (I40200), .I (g30377));
INVX1 gate14617(.O (g30540), .I (I40200));
INVX1 gate14618(.O (I40203), .I (g30380));
INVX1 gate14619(.O (g30541), .I (I40203));
INVX1 gate14620(.O (I40206), .I (g30450));
INVX1 gate14621(.O (g30542), .I (I40206));
INVX1 gate14622(.O (I40209), .I (g30459));
INVX1 gate14623(.O (g30543), .I (I40209));
INVX1 gate14624(.O (I40212), .I (g30471));
INVX1 gate14625(.O (g30544), .I (I40212));
INVX1 gate14626(.O (I40215), .I (g30501));
INVX1 gate14627(.O (g30545), .I (I40215));
INVX1 gate14628(.O (I40218), .I (g30335));
INVX1 gate14629(.O (g30546), .I (I40218));
INVX1 gate14630(.O (I40221), .I (g30349));
INVX1 gate14631(.O (g30547), .I (I40221));
INVX1 gate14632(.O (I40224), .I (g30336));
INVX1 gate14633(.O (g30548), .I (I40224));
INVX1 gate14634(.O (I40227), .I (g30350));
INVX1 gate14635(.O (g30549), .I (I40227));
INVX1 gate14636(.O (I40230), .I (g30362));
INVX1 gate14637(.O (g30550), .I (I40230));
INVX1 gate14638(.O (I40233), .I (g30363));
INVX1 gate14639(.O (g30551), .I (I40233));
INVX1 gate14640(.O (I40236), .I (g30373));
INVX1 gate14641(.O (g30552), .I (I40236));
INVX1 gate14642(.O (I40239), .I (g30378));
INVX1 gate14643(.O (g30553), .I (I40239));
INVX1 gate14644(.O (I40242), .I (g30379));
INVX1 gate14645(.O (g30554), .I (I40242));
INVX1 gate14646(.O (I40245), .I (g30381));
INVX1 gate14647(.O (g30555), .I (I40245));
INVX1 gate14648(.O (I40248), .I (g30382));
INVX1 gate14649(.O (g30556), .I (I40248));
INVX1 gate14650(.O (I40251), .I (g30463));
INVX1 gate14651(.O (g30557), .I (I40251));
INVX1 gate14652(.O (I40254), .I (g30474));
INVX1 gate14653(.O (g30558), .I (I40254));
INVX1 gate14654(.O (I40257), .I (g30488));
INVX1 gate14655(.O (g30559), .I (I40257));
INVX1 gate14656(.O (I40260), .I (g30339));
INVX1 gate14657(.O (g30560), .I (I40260));
INVX1 gate14658(.O (I40263), .I (g30353));
INVX1 gate14659(.O (g30561), .I (I40263));
INVX1 gate14660(.O (I40266), .I (g30365));
INVX1 gate14661(.O (g30562), .I (I40266));
INVX1 gate14662(.O (I40269), .I (g30354));
INVX1 gate14663(.O (g30563), .I (I40269));
INVX1 gate14664(.O (I40272), .I (g30366));
INVX1 gate14665(.O (g30564), .I (I40272));
INVX1 gate14666(.O (I40275), .I (g30375));
INVX1 gate14667(.O (g30565), .I (I40275));
INVX1 gate14668(.O (g30567), .I (g30403));
INVX1 gate14669(.O (g30568), .I (g30402));
INVX1 gate14670(.O (g30569), .I (g30406));
INVX1 gate14671(.O (g30570), .I (g30404));
INVX1 gate14672(.O (g30571), .I (g30401));
INVX1 gate14673(.O (g30572), .I (g30399));
INVX1 gate14674(.O (g30573), .I (g30405));
INVX1 gate14675(.O (g30574), .I (g30400));
INVX1 gate14676(.O (g30575), .I (g30412));
INVX1 gate14677(.O (I40288), .I (g30455));
INVX1 gate14678(.O (g30578), .I (I40288));
INVX1 gate14679(.O (I40291), .I (g30468));
INVX1 gate14680(.O (g30579), .I (I40291));
INVX1 gate14681(.O (I40294), .I (g30470));
INVX1 gate14682(.O (g30580), .I (I40294));
INVX1 gate14683(.O (I40297), .I (g30482));
INVX1 gate14684(.O (g30581), .I (I40297));
INVX1 gate14685(.O (I40300), .I (g30485));
INVX1 gate14686(.O (g30582), .I (I40300));
INVX1 gate14687(.O (I40303), .I (g30487));
INVX1 gate14688(.O (g30583), .I (I40303));
INVX1 gate14689(.O (I40307), .I (g30500));
INVX1 gate14690(.O (g30585), .I (I40307));
INVX1 gate14691(.O (I40310), .I (g30503));
INVX1 gate14692(.O (g30586), .I (I40310));
INVX1 gate14693(.O (I40313), .I (g30505));
INVX1 gate14694(.O (g30587), .I (I40313));
INVX1 gate14695(.O (I40317), .I (g30338));
INVX1 gate14696(.O (g30591), .I (I40317));
INVX1 gate14697(.O (I40320), .I (g30341));
INVX1 gate14698(.O (g30592), .I (I40320));
INVX1 gate14699(.O (I40326), .I (g30356));
INVX1 gate14700(.O (g30600), .I (I40326));
INVX1 gate14701(.O (I40420), .I (g30578));
INVX1 gate14702(.O (g30710), .I (I40420));
INVX1 gate14703(.O (I40423), .I (g30579));
INVX1 gate14704(.O (g30711), .I (I40423));
INVX1 gate14705(.O (I40426), .I (g30581));
INVX1 gate14706(.O (g30712), .I (I40426));
INVX1 gate14707(.O (I40429), .I (g30580));
INVX1 gate14708(.O (g30713), .I (I40429));
INVX1 gate14709(.O (I40432), .I (g30582));
INVX1 gate14710(.O (g30714), .I (I40432));
INVX1 gate14711(.O (I40435), .I (g30585));
INVX1 gate14712(.O (g30715), .I (I40435));
INVX1 gate14713(.O (I40438), .I (g30583));
INVX1 gate14714(.O (g30716), .I (I40438));
INVX1 gate14715(.O (I40441), .I (g30586));
INVX1 gate14716(.O (g30717), .I (I40441));
INVX1 gate14717(.O (I40444), .I (g30591));
INVX1 gate14718(.O (g30718), .I (I40444));
INVX1 gate14719(.O (I40447), .I (g30587));
INVX1 gate14720(.O (g30719), .I (I40447));
INVX1 gate14721(.O (I40450), .I (g30592));
INVX1 gate14722(.O (g30720), .I (I40450));
INVX1 gate14723(.O (I40453), .I (g30600));
INVX1 gate14724(.O (g30721), .I (I40453));
INVX1 gate14725(.O (I40456), .I (g30668));
INVX1 gate14726(.O (g30722), .I (I40456));
INVX1 gate14727(.O (I40459), .I (g30669));
INVX1 gate14728(.O (g30723), .I (I40459));
INVX1 gate14729(.O (I40462), .I (g30670));
INVX1 gate14730(.O (g30724), .I (I40462));
INVX1 gate14731(.O (I40465), .I (g30671));
INVX1 gate14732(.O (g30725), .I (I40465));
INVX1 gate14733(.O (I40468), .I (g30672));
INVX1 gate14734(.O (g30726), .I (I40468));
INVX1 gate14735(.O (I40471), .I (g30673));
INVX1 gate14736(.O (g30727), .I (I40471));
INVX1 gate14737(.O (I40475), .I (g30674));
INVX1 gate14738(.O (g30729), .I (I40475));
INVX1 gate14739(.O (I40478), .I (g30675));
INVX1 gate14740(.O (g30730), .I (I40478));
INVX1 gate14741(.O (I40481), .I (g30676));
INVX1 gate14742(.O (g30731), .I (I40481));
INVX1 gate14743(.O (I40484), .I (g30677));
INVX1 gate14744(.O (g30732), .I (I40484));
INVX1 gate14745(.O (I40487), .I (g30678));
INVX1 gate14746(.O (g30733), .I (I40487));
INVX1 gate14747(.O (I40490), .I (g30679));
INVX1 gate14748(.O (g30734), .I (I40490));
INVX1 gate14749(.O (I40495), .I (g30680));
INVX1 gate14750(.O (g30737), .I (I40495));
INVX1 gate14751(.O (I40498), .I (g30681));
INVX1 gate14752(.O (g30738), .I (I40498));
INVX1 gate14753(.O (I40501), .I (g30682));
INVX1 gate14754(.O (g30739), .I (I40501));
INVX1 gate14755(.O (I40504), .I (g30683));
INVX1 gate14756(.O (g30740), .I (I40504));
INVX1 gate14757(.O (I40507), .I (g30684));
INVX1 gate14758(.O (g30741), .I (I40507));
INVX1 gate14759(.O (I40510), .I (g30686));
INVX1 gate14760(.O (g30742), .I (I40510));
INVX1 gate14761(.O (I40515), .I (g30687));
INVX1 gate14762(.O (g30745), .I (I40515));
INVX1 gate14763(.O (I40518), .I (g30688));
INVX1 gate14764(.O (g30746), .I (I40518));
INVX1 gate14765(.O (I40521), .I (g30689));
INVX1 gate14766(.O (g30747), .I (I40521));
INVX1 gate14767(.O (I40524), .I (g30690));
INVX1 gate14768(.O (g30748), .I (I40524));
INVX1 gate14769(.O (I40527), .I (g30691));
INVX1 gate14770(.O (g30749), .I (I40527));
INVX1 gate14771(.O (I40531), .I (g30692));
INVX1 gate14772(.O (g30751), .I (I40531));
INVX1 gate14773(.O (I40534), .I (g30693));
INVX1 gate14774(.O (g30752), .I (I40534));
INVX1 gate14775(.O (I40537), .I (g30694));
INVX1 gate14776(.O (g30753), .I (I40537));
INVX1 gate14777(.O (I40542), .I (g30695));
INVX1 gate14778(.O (g30756), .I (I40542));
INVX1 gate14779(.O (g30765), .I (g30685));
INVX1 gate14780(.O (I40555), .I (g30699));
INVX1 gate14781(.O (g30767), .I (I40555));
INVX1 gate14782(.O (I40565), .I (g30700));
INVX1 gate14783(.O (g30769), .I (I40565));
INVX1 gate14784(.O (I40568), .I (g30701));
INVX1 gate14785(.O (g30770), .I (I40568));
INVX1 gate14786(.O (I40578), .I (g30702));
INVX1 gate14787(.O (g30772), .I (I40578));
INVX1 gate14788(.O (I40581), .I (g30703));
INVX1 gate14789(.O (g30773), .I (I40581));
INVX1 gate14790(.O (I40584), .I (g30704));
INVX1 gate14791(.O (g30774), .I (I40584));
INVX1 gate14792(.O (I40594), .I (g30705));
INVX1 gate14793(.O (g30776), .I (I40594));
INVX1 gate14794(.O (I40597), .I (g30706));
INVX1 gate14795(.O (g30777), .I (I40597));
INVX1 gate14796(.O (I40600), .I (g30707));
INVX1 gate14797(.O (g30778), .I (I40600));
INVX1 gate14798(.O (I40611), .I (g30708));
INVX1 gate14799(.O (g30781), .I (I40611));
INVX1 gate14800(.O (I40614), .I (g30709));
INVX1 gate14801(.O (g30782), .I (I40614));
INVX1 gate14802(.O (I40618), .I (g30566));
INVX1 gate14803(.O (g30784), .I (I40618));
INVX1 gate14804(.O (I40634), .I (g30571));
INVX1 gate14805(.O (g30792), .I (I40634));
INVX1 gate14806(.O (I40637), .I (g30570));
INVX1 gate14807(.O (g30793), .I (I40637));
INVX1 gate14808(.O (I40640), .I (g30569));
INVX1 gate14809(.O (g30794), .I (I40640));
INVX1 gate14810(.O (I40643), .I (g30568));
INVX1 gate14811(.O (g30795), .I (I40643));
INVX1 gate14812(.O (I40647), .I (g30567));
INVX1 gate14813(.O (g30797), .I (I40647));
INVX1 gate14814(.O (I40651), .I (g30574));
INVX1 gate14815(.O (g30799), .I (I40651));
INVX1 gate14816(.O (I40654), .I (g30573));
INVX1 gate14817(.O (g30800), .I (I40654));
INVX1 gate14818(.O (I40658), .I (g30572));
INVX1 gate14819(.O (g30802), .I (I40658));
INVX1 gate14820(.O (I40661), .I (g30635));
INVX1 gate14821(.O (g30803), .I (I40661));
INVX1 gate14822(.O (I40664), .I (g30636));
INVX1 gate14823(.O (g30804), .I (I40664));
INVX1 gate14824(.O (I40667), .I (g30637));
INVX1 gate14825(.O (g30805), .I (I40667));
INVX1 gate14826(.O (I40670), .I (g30638));
INVX1 gate14827(.O (g30806), .I (I40670));
INVX1 gate14828(.O (I40673), .I (g30639));
INVX1 gate14829(.O (g30807), .I (I40673));
INVX1 gate14830(.O (I40676), .I (g30640));
INVX1 gate14831(.O (g30808), .I (I40676));
INVX1 gate14832(.O (I40679), .I (g30641));
INVX1 gate14833(.O (g30809), .I (I40679));
INVX1 gate14834(.O (I40682), .I (g30642));
INVX1 gate14835(.O (g30810), .I (I40682));
INVX1 gate14836(.O (I40685), .I (g30643));
INVX1 gate14837(.O (g30811), .I (I40685));
INVX1 gate14838(.O (I40688), .I (g30644));
INVX1 gate14839(.O (g30812), .I (I40688));
INVX1 gate14840(.O (I40691), .I (g30645));
INVX1 gate14841(.O (g30813), .I (I40691));
INVX1 gate14842(.O (I40694), .I (g30646));
INVX1 gate14843(.O (g30814), .I (I40694));
INVX1 gate14844(.O (I40697), .I (g30647));
INVX1 gate14845(.O (g30815), .I (I40697));
INVX1 gate14846(.O (I40700), .I (g30648));
INVX1 gate14847(.O (g30816), .I (I40700));
INVX1 gate14848(.O (I40703), .I (g30649));
INVX1 gate14849(.O (g30817), .I (I40703));
INVX1 gate14850(.O (I40706), .I (g30650));
INVX1 gate14851(.O (g30818), .I (I40706));
INVX1 gate14852(.O (I40709), .I (g30651));
INVX1 gate14853(.O (g30819), .I (I40709));
INVX1 gate14854(.O (I40712), .I (g30652));
INVX1 gate14855(.O (g30820), .I (I40712));
INVX1 gate14856(.O (I40715), .I (g30653));
INVX1 gate14857(.O (g30821), .I (I40715));
INVX1 gate14858(.O (I40718), .I (g30654));
INVX1 gate14859(.O (g30822), .I (I40718));
INVX1 gate14860(.O (I40721), .I (g30655));
INVX1 gate14861(.O (g30823), .I (I40721));
INVX1 gate14862(.O (I40724), .I (g30656));
INVX1 gate14863(.O (g30824), .I (I40724));
INVX1 gate14864(.O (I40727), .I (g30657));
INVX1 gate14865(.O (g30825), .I (I40727));
INVX1 gate14866(.O (I40730), .I (g30658));
INVX1 gate14867(.O (g30826), .I (I40730));
INVX1 gate14868(.O (I40733), .I (g30659));
INVX1 gate14869(.O (g30827), .I (I40733));
INVX1 gate14870(.O (I40736), .I (g30660));
INVX1 gate14871(.O (g30828), .I (I40736));
INVX1 gate14872(.O (I40739), .I (g30661));
INVX1 gate14873(.O (g30829), .I (I40739));
INVX1 gate14874(.O (I40742), .I (g30662));
INVX1 gate14875(.O (g30830), .I (I40742));
INVX1 gate14876(.O (I40745), .I (g30663));
INVX1 gate14877(.O (g30831), .I (I40745));
INVX1 gate14878(.O (I40748), .I (g30664));
INVX1 gate14879(.O (g30832), .I (I40748));
INVX1 gate14880(.O (I40751), .I (g30665));
INVX1 gate14881(.O (g30833), .I (I40751));
INVX1 gate14882(.O (I40754), .I (g30666));
INVX1 gate14883(.O (g30834), .I (I40754));
INVX1 gate14884(.O (I40757), .I (g30667));
INVX1 gate14885(.O (g30835), .I (I40757));
INVX1 gate14886(.O (I40760), .I (g30722));
INVX1 gate14887(.O (g30836), .I (I40760));
INVX1 gate14888(.O (I40763), .I (g30729));
INVX1 gate14889(.O (g30837), .I (I40763));
INVX1 gate14890(.O (I40766), .I (g30737));
INVX1 gate14891(.O (g30838), .I (I40766));
INVX1 gate14892(.O (I40769), .I (g30803));
INVX1 gate14893(.O (g30839), .I (I40769));
INVX1 gate14894(.O (I40772), .I (g30804));
INVX1 gate14895(.O (g30840), .I (I40772));
INVX1 gate14896(.O (I40775), .I (g30807));
INVX1 gate14897(.O (g30841), .I (I40775));
INVX1 gate14898(.O (I40778), .I (g30805));
INVX1 gate14899(.O (g30842), .I (I40778));
INVX1 gate14900(.O (I40781), .I (g30808));
INVX1 gate14901(.O (g30843), .I (I40781));
INVX1 gate14902(.O (I40784), .I (g30813));
INVX1 gate14903(.O (g30844), .I (I40784));
INVX1 gate14904(.O (I40787), .I (g30809));
INVX1 gate14905(.O (g30845), .I (I40787));
INVX1 gate14906(.O (I40790), .I (g30814));
INVX1 gate14907(.O (g30846), .I (I40790));
INVX1 gate14908(.O (I40793), .I (g30821));
INVX1 gate14909(.O (g30847), .I (I40793));
INVX1 gate14910(.O (I40796), .I (g30829));
INVX1 gate14911(.O (g30848), .I (I40796));
INVX1 gate14912(.O (I40799), .I (g30723));
INVX1 gate14913(.O (g30849), .I (I40799));
INVX1 gate14914(.O (I40802), .I (g30730));
INVX1 gate14915(.O (g30850), .I (I40802));
INVX1 gate14916(.O (I40805), .I (g30767));
INVX1 gate14917(.O (g30851), .I (I40805));
INVX1 gate14918(.O (I40808), .I (g30769));
INVX1 gate14919(.O (g30852), .I (I40808));
INVX1 gate14920(.O (I40811), .I (g30772));
INVX1 gate14921(.O (g30853), .I (I40811));
INVX1 gate14922(.O (I40814), .I (g30731));
INVX1 gate14923(.O (g30854), .I (I40814));
INVX1 gate14924(.O (I40817), .I (g30738));
INVX1 gate14925(.O (g30855), .I (I40817));
INVX1 gate14926(.O (I40820), .I (g30745));
INVX1 gate14927(.O (g30856), .I (I40820));
INVX1 gate14928(.O (I40823), .I (g30806));
INVX1 gate14929(.O (g30857), .I (I40823));
INVX1 gate14930(.O (I40826), .I (g30810));
INVX1 gate14931(.O (g30858), .I (I40826));
INVX1 gate14932(.O (I40829), .I (g30815));
INVX1 gate14933(.O (g30859), .I (I40829));
INVX1 gate14934(.O (I40832), .I (g30811));
INVX1 gate14935(.O (g30860), .I (I40832));
INVX1 gate14936(.O (I40835), .I (g30816));
INVX1 gate14937(.O (g30861), .I (I40835));
INVX1 gate14938(.O (I40838), .I (g30822));
INVX1 gate14939(.O (g30862), .I (I40838));
INVX1 gate14940(.O (I40841), .I (g30817));
INVX1 gate14941(.O (g30863), .I (I40841));
INVX1 gate14942(.O (I40844), .I (g30823));
INVX1 gate14943(.O (g30864), .I (I40844));
INVX1 gate14944(.O (I40847), .I (g30830));
INVX1 gate14945(.O (g30865), .I (I40847));
INVX1 gate14946(.O (I40850), .I (g30724));
INVX1 gate14947(.O (g30866), .I (I40850));
INVX1 gate14948(.O (I40853), .I (g30732));
INVX1 gate14949(.O (g30867), .I (I40853));
INVX1 gate14950(.O (I40856), .I (g30739));
INVX1 gate14951(.O (g30868), .I (I40856));
INVX1 gate14952(.O (I40859), .I (g30770));
INVX1 gate14953(.O (g30869), .I (I40859));
INVX1 gate14954(.O (I40862), .I (g30773));
INVX1 gate14955(.O (g30870), .I (I40862));
INVX1 gate14956(.O (I40865), .I (g30776));
INVX1 gate14957(.O (g30871), .I (I40865));
INVX1 gate14958(.O (I40868), .I (g30740));
INVX1 gate14959(.O (g30872), .I (I40868));
INVX1 gate14960(.O (I40871), .I (g30746));
INVX1 gate14961(.O (g30873), .I (I40871));
INVX1 gate14962(.O (I40874), .I (g30751));
INVX1 gate14963(.O (g30874), .I (I40874));
INVX1 gate14964(.O (I40877), .I (g30812));
INVX1 gate14965(.O (g30875), .I (I40877));
INVX1 gate14966(.O (I40880), .I (g30818));
INVX1 gate14967(.O (g30876), .I (I40880));
INVX1 gate14968(.O (I40883), .I (g30824));
INVX1 gate14969(.O (g30877), .I (I40883));
INVX1 gate14970(.O (I40886), .I (g30819));
INVX1 gate14971(.O (g30878), .I (I40886));
INVX1 gate14972(.O (I40889), .I (g30825));
INVX1 gate14973(.O (g30879), .I (I40889));
INVX1 gate14974(.O (I40892), .I (g30831));
INVX1 gate14975(.O (g30880), .I (I40892));
INVX1 gate14976(.O (I40895), .I (g30826));
INVX1 gate14977(.O (g30881), .I (I40895));
INVX1 gate14978(.O (I40898), .I (g30832));
INVX1 gate14979(.O (g30882), .I (I40898));
INVX1 gate14980(.O (I40901), .I (g30725));
INVX1 gate14981(.O (g30883), .I (I40901));
INVX1 gate14982(.O (I40904), .I (g30733));
INVX1 gate14983(.O (g30884), .I (I40904));
INVX1 gate14984(.O (I40907), .I (g30741));
INVX1 gate14985(.O (g30885), .I (I40907));
INVX1 gate14986(.O (I40910), .I (g30747));
INVX1 gate14987(.O (g30886), .I (I40910));
INVX1 gate14988(.O (I40913), .I (g30774));
INVX1 gate14989(.O (g30887), .I (I40913));
INVX1 gate14990(.O (I40916), .I (g30777));
INVX1 gate14991(.O (g30888), .I (I40916));
INVX1 gate14992(.O (I40919), .I (g30781));
INVX1 gate14993(.O (g30889), .I (I40919));
INVX1 gate14994(.O (I40922), .I (g30748));
INVX1 gate14995(.O (g30890), .I (I40922));
INVX1 gate14996(.O (I40925), .I (g30752));
INVX1 gate14997(.O (g30891), .I (I40925));
INVX1 gate14998(.O (I40928), .I (g30756));
INVX1 gate14999(.O (g30892), .I (I40928));
INVX1 gate15000(.O (I40931), .I (g30820));
INVX1 gate15001(.O (g30893), .I (I40931));
INVX1 gate15002(.O (I40934), .I (g30827));
INVX1 gate15003(.O (g30894), .I (I40934));
INVX1 gate15004(.O (I40937), .I (g30833));
INVX1 gate15005(.O (g30895), .I (I40937));
INVX1 gate15006(.O (I40940), .I (g30828));
INVX1 gate15007(.O (g30896), .I (I40940));
INVX1 gate15008(.O (I40943), .I (g30834));
INVX1 gate15009(.O (g30897), .I (I40943));
INVX1 gate15010(.O (I40946), .I (g30726));
INVX1 gate15011(.O (g30898), .I (I40946));
INVX1 gate15012(.O (I40949), .I (g30835));
INVX1 gate15013(.O (g30899), .I (I40949));
INVX1 gate15014(.O (I40952), .I (g30727));
INVX1 gate15015(.O (g30900), .I (I40952));
INVX1 gate15016(.O (I40955), .I (g30734));
INVX1 gate15017(.O (g30901), .I (I40955));
INVX1 gate15018(.O (I40958), .I (g30742));
INVX1 gate15019(.O (g30902), .I (I40958));
INVX1 gate15020(.O (I40961), .I (g30749));
INVX1 gate15021(.O (g30903), .I (I40961));
INVX1 gate15022(.O (I40964), .I (g30753));
INVX1 gate15023(.O (g30904), .I (I40964));
INVX1 gate15024(.O (I40967), .I (g30778));
INVX1 gate15025(.O (g30905), .I (I40967));
INVX1 gate15026(.O (I40970), .I (g30782));
INVX1 gate15027(.O (g30906), .I (I40970));
INVX1 gate15028(.O (I40973), .I (g30784));
INVX1 gate15029(.O (g30907), .I (I40973));
INVX1 gate15030(.O (I40976), .I (g30799));
INVX1 gate15031(.O (g30908), .I (I40976));
INVX1 gate15032(.O (I40979), .I (g30800));
INVX1 gate15033(.O (g30909), .I (I40979));
INVX1 gate15034(.O (I40982), .I (g30802));
INVX1 gate15035(.O (g30910), .I (I40982));
INVX1 gate15036(.O (I40985), .I (g30792));
INVX1 gate15037(.O (g30911), .I (I40985));
INVX1 gate15038(.O (I40988), .I (g30793));
INVX1 gate15039(.O (g30912), .I (I40988));
INVX1 gate15040(.O (I40991), .I (g30794));
INVX1 gate15041(.O (g30913), .I (I40991));
INVX1 gate15042(.O (I40994), .I (g30795));
INVX1 gate15043(.O (g30914), .I (I40994));
INVX1 gate15044(.O (I40997), .I (g30797));
INVX1 gate15045(.O (g30915), .I (I40997));
INVX1 gate15046(.O (I41024), .I (g30765));
INVX1 gate15047(.O (g30928), .I (I41024));
INVX1 gate15048(.O (I41035), .I (g30796));
INVX1 gate15049(.O (g30937), .I (I41035));
INVX1 gate15050(.O (I41038), .I (g30798));
INVX1 gate15051(.O (g30938), .I (I41038));
INVX1 gate15052(.O (I41041), .I (g30801));
INVX1 gate15053(.O (g30939), .I (I41041));
INVX1 gate15054(.O (I41044), .I (g30928));
INVX1 gate15055(.O (g30940), .I (I41044));
INVX1 gate15056(.O (I41047), .I (g30937));
INVX1 gate15057(.O (g30941), .I (I41047));
INVX1 gate15058(.O (I41050), .I (g30938));
INVX1 gate15059(.O (g30942), .I (I41050));
INVX1 gate15060(.O (I41053), .I (g30939));
INVX1 gate15061(.O (g30943), .I (I41053));
INVX1 gate15062(.O (g30962), .I (g30958));
INVX1 gate15063(.O (g30963), .I (g30957));
INVX1 gate15064(.O (g30964), .I (g30961));
INVX1 gate15065(.O (g30965), .I (g30959));
INVX1 gate15066(.O (g30966), .I (g30956));
INVX1 gate15067(.O (g30967), .I (g30954));
INVX1 gate15068(.O (g30968), .I (g30960));
INVX1 gate15069(.O (g30969), .I (g30955));
INVX1 gate15070(.O (g30971), .I (g30970));
INVX1 gate15071(.O (I41090), .I (g30965));
INVX1 gate15072(.O (g30972), .I (I41090));
INVX1 gate15073(.O (I41093), .I (g30964));
INVX1 gate15074(.O (g30973), .I (I41093));
INVX1 gate15075(.O (I41096), .I (g30963));
INVX1 gate15076(.O (g30974), .I (I41096));
INVX1 gate15077(.O (I41099), .I (g30962));
INVX1 gate15078(.O (g30975), .I (I41099));
INVX1 gate15079(.O (I41102), .I (g30969));
INVX1 gate15080(.O (g30976), .I (I41102));
INVX1 gate15081(.O (I41105), .I (g30968));
INVX1 gate15082(.O (g30977), .I (I41105));
INVX1 gate15083(.O (I41108), .I (g30967));
INVX1 gate15084(.O (g30978), .I (I41108));
INVX1 gate15085(.O (I41111), .I (g30966));
INVX1 gate15086(.O (g30979), .I (I41111));
INVX1 gate15087(.O (I41114), .I (g30976));
INVX1 gate15088(.O (g30980), .I (I41114));
INVX1 gate15089(.O (I41117), .I (g30977));
INVX1 gate15090(.O (g30981), .I (I41117));
INVX1 gate15091(.O (I41120), .I (g30978));
INVX1 gate15092(.O (g30982), .I (I41120));
INVX1 gate15093(.O (I41123), .I (g30979));
INVX1 gate15094(.O (g30983), .I (I41123));
INVX1 gate15095(.O (I41126), .I (g30972));
INVX1 gate15096(.O (g30984), .I (I41126));
INVX1 gate15097(.O (I41129), .I (g30973));
INVX1 gate15098(.O (g30985), .I (I41129));
INVX1 gate15099(.O (I41132), .I (g30974));
INVX1 gate15100(.O (g30986), .I (I41132));
INVX1 gate15101(.O (I41135), .I (g30975));
INVX1 gate15102(.O (g30987), .I (I41135));
INVX1 gate15103(.O (I41138), .I (g30971));
INVX1 gate15104(.O (g30988), .I (I41138));
INVX1 gate15105(.O (I41141), .I (g30988));
INVX1 gate15106(.O (g30989), .I (I41141));
AN2X1 gate15107(.O (g5630), .I1 (g325), .I2 (g349));
AN2X1 gate15108(.O (g5649), .I1 (g331), .I2 (g351));
AN2X1 gate15109(.O (g5650), .I1 (g325), .I2 (g364));
AN2X1 gate15110(.O (g5658), .I1 (g1012), .I2 (g1036));
AN2X1 gate15111(.O (g5676), .I1 (g337), .I2 (g353));
AN2X1 gate15112(.O (g5677), .I1 (g331), .I2 (g366));
AN2X1 gate15113(.O (g5678), .I1 (g325), .I2 (g379));
AN2X1 gate15114(.O (g5687), .I1 (g1018), .I2 (g1038));
AN2X1 gate15115(.O (g5688), .I1 (g1012), .I2 (g1051));
AN2X1 gate15116(.O (g5696), .I1 (g1706), .I2 (g1730));
AN2X1 gate15117(.O (g5709), .I1 (g337), .I2 (g368));
AN2X1 gate15118(.O (g5710), .I1 (g331), .I2 (g381));
AN2X1 gate15119(.O (g5711), .I1 (g325), .I2 (g394));
AN2X1 gate15120(.O (g5728), .I1 (g1024), .I2 (g1040));
AN2X1 gate15121(.O (g5729), .I1 (g1018), .I2 (g1053));
AN2X1 gate15122(.O (g5730), .I1 (g1012), .I2 (g1066));
AN2X1 gate15123(.O (g5739), .I1 (g1712), .I2 (g1732));
AN2X1 gate15124(.O (g5740), .I1 (g1706), .I2 (g1745));
AN2X1 gate15125(.O (g5748), .I1 (g2400), .I2 (g2424));
AN2X1 gate15126(.O (g5757), .I1 (g337), .I2 (g383));
AN2X1 gate15127(.O (g5758), .I1 (g331), .I2 (g396));
AN2X1 gate15128(.O (g5767), .I1 (g1024), .I2 (g1055));
AN2X1 gate15129(.O (g5768), .I1 (g1018), .I2 (g1068));
AN2X1 gate15130(.O (g5769), .I1 (g1012), .I2 (g1081));
AN2X1 gate15131(.O (g5786), .I1 (g1718), .I2 (g1734));
AN2X1 gate15132(.O (g5787), .I1 (g1712), .I2 (g1747));
AN2X1 gate15133(.O (g5788), .I1 (g1706), .I2 (g1760));
AN2X1 gate15134(.O (g5797), .I1 (g2406), .I2 (g2426));
AN2X1 gate15135(.O (g5798), .I1 (g2400), .I2 (g2439));
AN2X1 gate15136(.O (g5807), .I1 (g337), .I2 (g324));
AN2X1 gate15137(.O (g5816), .I1 (g1024), .I2 (g1070));
AN2X1 gate15138(.O (g5817), .I1 (g1018), .I2 (g1083));
AN2X1 gate15139(.O (g5826), .I1 (g1718), .I2 (g1749));
AN2X1 gate15140(.O (g5827), .I1 (g1712), .I2 (g1762));
AN2X1 gate15141(.O (g5828), .I1 (g1706), .I2 (g1775));
AN2X1 gate15142(.O (g5845), .I1 (g2412), .I2 (g2428));
AN2X1 gate15143(.O (g5846), .I1 (g2406), .I2 (g2441));
AN2X1 gate15144(.O (g5847), .I1 (g2400), .I2 (g2454));
AN2X1 gate15145(.O (g5863), .I1 (g1024), .I2 (g1011));
AN2X1 gate15146(.O (g5872), .I1 (g1718), .I2 (g1764));
AN2X1 gate15147(.O (g5873), .I1 (g1712), .I2 (g1777));
AN2X1 gate15148(.O (g5882), .I1 (g2412), .I2 (g2443));
AN2X1 gate15149(.O (g5883), .I1 (g2406), .I2 (g2456));
AN2X1 gate15150(.O (g5884), .I1 (g2400), .I2 (g2469));
AN2X1 gate15151(.O (g5910), .I1 (g1718), .I2 (g1705));
AN2X1 gate15152(.O (g5919), .I1 (g2412), .I2 (g2458));
AN2X1 gate15153(.O (g5920), .I1 (g2406), .I2 (g2471));
AN2X1 gate15154(.O (g5949), .I1 (g2412), .I2 (g2399));
AN2X1 gate15155(.O (g8327), .I1 (g3254), .I2 (g219));
AN2X1 gate15156(.O (g8328), .I1 (g6314), .I2 (g225));
AN2X1 gate15157(.O (g8329), .I1 (g6232), .I2 (g231));
AN2X1 gate15158(.O (g8339), .I1 (g6519), .I2 (g903));
AN2X1 gate15159(.O (g8340), .I1 (g6369), .I2 (g909));
AN2X1 gate15160(.O (g8350), .I1 (g6574), .I2 (g1594));
AN2X1 gate15161(.O (g8385), .I1 (g3254), .I2 (g228));
AN2X1 gate15162(.O (g8386), .I1 (g6314), .I2 (g234));
AN2X1 gate15163(.O (g8387), .I1 (g6232), .I2 (g240));
AN2X1 gate15164(.O (g8394), .I1 (g3410), .I2 (g906));
AN2X1 gate15165(.O (g8395), .I1 (g6519), .I2 (g912));
AN2X1 gate15166(.O (g8396), .I1 (g6369), .I2 (g918));
AN2X1 gate15167(.O (g8406), .I1 (g6783), .I2 (g1597));
AN2X1 gate15168(.O (g8407), .I1 (g6574), .I2 (g1603));
AN2X1 gate15169(.O (g8417), .I1 (g6838), .I2 (g2288));
AN2X1 gate15170(.O (g8431), .I1 (g3254), .I2 (g237));
AN2X1 gate15171(.O (g8432), .I1 (g6314), .I2 (g243));
AN2X1 gate15172(.O (g8433), .I1 (g6232), .I2 (g249));
AN2X1 gate15173(.O (g8437), .I1 (g3410), .I2 (g915));
AN2X1 gate15174(.O (g8438), .I1 (g6519), .I2 (g921));
AN2X1 gate15175(.O (g8439), .I1 (g6369), .I2 (g927));
AN2X1 gate15176(.O (g8446), .I1 (g3566), .I2 (g1600));
AN2X1 gate15177(.O (g8447), .I1 (g6783), .I2 (g1606));
AN2X1 gate15178(.O (g8448), .I1 (g6574), .I2 (g1612));
AN2X1 gate15179(.O (g8458), .I1 (g7085), .I2 (g2291));
AN2X1 gate15180(.O (g8459), .I1 (g6838), .I2 (g2297));
AN2X1 gate15181(.O (g8463), .I1 (g3254), .I2 (g246));
AN2X1 gate15182(.O (g8464), .I1 (g6314), .I2 (g252));
AN2X1 gate15183(.O (g8465), .I1 (g6232), .I2 (g258));
AN2X1 gate15184(.O (g8466), .I1 (g3410), .I2 (g924));
AN2X1 gate15185(.O (g8467), .I1 (g6519), .I2 (g930));
AN2X1 gate15186(.O (g8468), .I1 (g6369), .I2 (g936));
AN2X1 gate15187(.O (g8472), .I1 (g3566), .I2 (g1609));
AN2X1 gate15188(.O (g8473), .I1 (g6783), .I2 (g1615));
AN2X1 gate15189(.O (g8474), .I1 (g6574), .I2 (g1621));
AN2X1 gate15190(.O (g8481), .I1 (g3722), .I2 (g2294));
AN2X1 gate15191(.O (g8482), .I1 (g7085), .I2 (g2300));
AN2X1 gate15192(.O (g8483), .I1 (g6838), .I2 (g2306));
AN2X1 gate15193(.O (g8484), .I1 (g6232), .I2 (g186));
AN2X1 gate15194(.O (g8485), .I1 (g3254), .I2 (g255));
AN2X1 gate15195(.O (g8486), .I1 (g6314), .I2 (g261));
AN2X1 gate15196(.O (g8487), .I1 (g6232), .I2 (g267));
AN2X1 gate15197(.O (g8488), .I1 (g3410), .I2 (g933));
AN2X1 gate15198(.O (g8489), .I1 (g6519), .I2 (g939));
AN2X1 gate15199(.O (g8490), .I1 (g6369), .I2 (g945));
AN2X1 gate15200(.O (g8491), .I1 (g3566), .I2 (g1618));
AN2X1 gate15201(.O (g8492), .I1 (g6783), .I2 (g1624));
AN2X1 gate15202(.O (g8493), .I1 (g6574), .I2 (g1630));
AN2X1 gate15203(.O (g8497), .I1 (g3722), .I2 (g2303));
AN2X1 gate15204(.O (g8498), .I1 (g7085), .I2 (g2309));
AN2X1 gate15205(.O (g8499), .I1 (g6838), .I2 (g2315));
AN2X1 gate15206(.O (g8500), .I1 (g6314), .I2 (g189));
AN2X1 gate15207(.O (g8501), .I1 (g6232), .I2 (g195));
AN2X1 gate15208(.O (g8502), .I1 (g3254), .I2 (g264));
AN2X1 gate15209(.O (g8503), .I1 (g6314), .I2 (g270));
AN2X1 gate15210(.O (g8504), .I1 (g6369), .I2 (g873));
AN2X1 gate15211(.O (g8505), .I1 (g3410), .I2 (g942));
AN2X1 gate15212(.O (g8506), .I1 (g6519), .I2 (g948));
AN2X1 gate15213(.O (g8507), .I1 (g6369), .I2 (g954));
AN2X1 gate15214(.O (g8508), .I1 (g3566), .I2 (g1627));
AN2X1 gate15215(.O (g8509), .I1 (g6783), .I2 (g1633));
AN2X1 gate15216(.O (g8510), .I1 (g6574), .I2 (g1639));
AN2X1 gate15217(.O (g8511), .I1 (g3722), .I2 (g2312));
AN2X1 gate15218(.O (g8512), .I1 (g7085), .I2 (g2318));
AN2X1 gate15219(.O (g8513), .I1 (g6838), .I2 (g2324));
AN2X1 gate15220(.O (g8515), .I1 (g3254), .I2 (g192));
AN2X1 gate15221(.O (g8516), .I1 (g6314), .I2 (g198));
AN2X1 gate15222(.O (g8517), .I1 (g6232), .I2 (g204));
AN2X1 gate15223(.O (g8518), .I1 (g3254), .I2 (g273));
AN2X1 gate15224(.O (g8519), .I1 (g6519), .I2 (g876));
AN2X1 gate15225(.O (g8520), .I1 (g6369), .I2 (g882));
AN2X1 gate15226(.O (g8521), .I1 (g3410), .I2 (g951));
AN2X1 gate15227(.O (g8522), .I1 (g6519), .I2 (g957));
AN2X1 gate15228(.O (g8523), .I1 (g6574), .I2 (g1567));
AN2X1 gate15229(.O (g8524), .I1 (g3566), .I2 (g1636));
AN2X1 gate15230(.O (g8525), .I1 (g6783), .I2 (g1642));
AN2X1 gate15231(.O (g8526), .I1 (g6574), .I2 (g1648));
AN2X1 gate15232(.O (g8527), .I1 (g3722), .I2 (g2321));
AN2X1 gate15233(.O (g8528), .I1 (g7085), .I2 (g2327));
AN2X1 gate15234(.O (g8529), .I1 (g6838), .I2 (g2333));
AN2X1 gate15235(.O (g8531), .I1 (g3254), .I2 (g201));
AN2X1 gate15236(.O (g8532), .I1 (g6314), .I2 (g207));
AN2X1 gate15237(.O (g8534), .I1 (g3410), .I2 (g879));
AN2X1 gate15238(.O (g8535), .I1 (g6519), .I2 (g885));
AN2X1 gate15239(.O (g8536), .I1 (g6369), .I2 (g891));
AN2X1 gate15240(.O (g8537), .I1 (g3410), .I2 (g960));
AN2X1 gate15241(.O (g8538), .I1 (g6783), .I2 (g1570));
AN2X1 gate15242(.O (g8539), .I1 (g6574), .I2 (g1576));
AN2X1 gate15243(.O (g8540), .I1 (g3566), .I2 (g1645));
AN2X1 gate15244(.O (g8541), .I1 (g6783), .I2 (g1651));
AN2X1 gate15245(.O (g8542), .I1 (g6838), .I2 (g2261));
AN2X1 gate15246(.O (g8543), .I1 (g3722), .I2 (g2330));
AN2X1 gate15247(.O (g8544), .I1 (g7085), .I2 (g2336));
AN2X1 gate15248(.O (g8545), .I1 (g6838), .I2 (g2342));
AN2X1 gate15249(.O (g8546), .I1 (g3254), .I2 (g210));
AN2X1 gate15250(.O (g8548), .I1 (g3410), .I2 (g888));
AN2X1 gate15251(.O (g8549), .I1 (g6519), .I2 (g894));
AN2X1 gate15252(.O (g8551), .I1 (g3566), .I2 (g1573));
AN2X1 gate15253(.O (g8552), .I1 (g6783), .I2 (g1579));
AN2X1 gate15254(.O (g8553), .I1 (g6574), .I2 (g1585));
AN2X1 gate15255(.O (g8554), .I1 (g3566), .I2 (g1654));
AN2X1 gate15256(.O (g8555), .I1 (g7085), .I2 (g2264));
AN2X1 gate15257(.O (g8556), .I1 (g6838), .I2 (g2270));
AN2X1 gate15258(.O (g8557), .I1 (g3722), .I2 (g2339));
AN2X1 gate15259(.O (g8558), .I1 (g7085), .I2 (g2345));
AN2X1 gate15260(.O (g8559), .I1 (g3410), .I2 (g897));
AN2X1 gate15261(.O (g8561), .I1 (g3566), .I2 (g1582));
AN2X1 gate15262(.O (g8562), .I1 (g6783), .I2 (g1588));
AN2X1 gate15263(.O (g8564), .I1 (g3722), .I2 (g2267));
AN2X1 gate15264(.O (g8565), .I1 (g7085), .I2 (g2273));
AN2X1 gate15265(.O (g8566), .I1 (g6838), .I2 (g2279));
AN2X1 gate15266(.O (g8567), .I1 (g3722), .I2 (g2348));
AN2X1 gate15267(.O (g8570), .I1 (g3566), .I2 (g1591));
AN2X1 gate15268(.O (g8572), .I1 (g3722), .I2 (g2276));
AN2X1 gate15269(.O (g8573), .I1 (g7085), .I2 (g2282));
AN2X1 gate15270(.O (g8576), .I1 (g3722), .I2 (g2285));
AN2X1 gate15271(.O (g8601), .I1 (g6643), .I2 (g7153));
AN2X1 gate15272(.O (g8612), .I1 (g3338), .I2 (g6908));
AN2X1 gate15273(.O (g8613), .I1 (g6945), .I2 (g7349));
AN2X1 gate15274(.O (g8621), .I1 (g6486), .I2 (g6672));
AN2X1 gate15275(.O (g8625), .I1 (g3494), .I2 (g7158));
AN2X1 gate15276(.O (g8626), .I1 (g7195), .I2 (g7479));
AN2X1 gate15277(.O (g8631), .I1 (g6751), .I2 (g6974));
AN2X1 gate15278(.O (g8635), .I1 (g3650), .I2 (g7354));
AN2X1 gate15279(.O (g8636), .I1 (g7391), .I2 (g7535));
AN2X1 gate15280(.O (g8650), .I1 (g7053), .I2 (g7224));
AN2X1 gate15281(.O (g8654), .I1 (g3806), .I2 (g7484));
AN2X1 gate15282(.O (g8666), .I1 (g7303), .I2 (g7420));
AN2X1 gate15283(.O (g8676), .I1 (g6643), .I2 (g7838));
AN2X1 gate15284(.O (g8687), .I1 (g3338), .I2 (g7827));
AN2X1 gate15285(.O (g8688), .I1 (g6945), .I2 (g7858));
AN2X1 gate15286(.O (g8703), .I1 (g6486), .I2 (g7819));
AN2X1 gate15287(.O (g8704), .I1 (g6643), .I2 (g7996));
AN2X1 gate15288(.O (g8705), .I1 (g3494), .I2 (g7842));
AN2X1 gate15289(.O (g8706), .I1 (g7195), .I2 (g7888));
AN2X1 gate15290(.O (g8717), .I1 (g3338), .I2 (g7953));
AN2X1 gate15291(.O (g8722), .I1 (g6751), .I2 (g7830));
AN2X1 gate15292(.O (g8723), .I1 (g6945), .I2 (g8071));
AN2X1 gate15293(.O (g8724), .I1 (g3650), .I2 (g7862));
AN2X1 gate15294(.O (g8725), .I1 (g7391), .I2 (g7912));
AN2X1 gate15295(.O (g8751), .I1 (g6486), .I2 (g7906));
AN2X1 gate15296(.O (g8755), .I1 (g3494), .I2 (g8004));
AN2X1 gate15297(.O (g8760), .I1 (g7053), .I2 (g7845));
AN2X1 gate15298(.O (g8761), .I1 (g7195), .I2 (g8156));
AN2X1 gate15299(.O (g8762), .I1 (g3806), .I2 (g7892));
AN2X1 gate15300(.O (g8774), .I1 (g6751), .I2 (g7958));
AN2X1 gate15301(.O (g8778), .I1 (g3650), .I2 (g8079));
AN2X1 gate15302(.O (g8783), .I1 (g7303), .I2 (g7865));
AN2X1 gate15303(.O (g8784), .I1 (g7391), .I2 (g8242));
AN2X1 gate15304(.O (g8797), .I1 (g7053), .I2 (g8009));
AN2X1 gate15305(.O (g8801), .I1 (g3806), .I2 (g8164));
AN2X1 gate15306(.O (g8816), .I1 (g7303), .I2 (g8084));
AN2X1 gate15307(.O (g8841), .I1 (g6486), .I2 (g490));
AN2X1 gate15308(.O (g8842), .I1 (g6512), .I2 (g5508));
AN2X1 gate15309(.O (g8861), .I1 (g6643), .I2 (g493));
AN2X1 gate15310(.O (g8868), .I1 (g6751), .I2 (g1177));
AN2X1 gate15311(.O (g8869), .I1 (g6776), .I2 (g5552));
AN2X1 gate15312(.O (g8892), .I1 (g3338), .I2 (g496));
AN2X1 gate15313(.O (g8899), .I1 (g6945), .I2 (g1180));
AN2X1 gate15314(.O (g8906), .I1 (g7053), .I2 (g1871));
AN2X1 gate15315(.O (g8907), .I1 (g7078), .I2 (g5598));
AN2X1 gate15316(.O (g8932), .I1 (g3494), .I2 (g1183));
AN2X1 gate15317(.O (g8939), .I1 (g7195), .I2 (g1874));
AN2X1 gate15318(.O (g8946), .I1 (g7303), .I2 (g2565));
AN2X1 gate15319(.O (g8947), .I1 (g7328), .I2 (g5615));
AN2X1 gate15320(.O (g8972), .I1 (g3650), .I2 (g1877));
AN2X1 gate15321(.O (g8979), .I1 (g7391), .I2 (g2568));
AN2X1 gate15322(.O (g9004), .I1 (g3806), .I2 (g2571));
AN2X1 gate15323(.O (g9009), .I1 (g6486), .I2 (g565));
AN2X1 gate15324(.O (g9026), .I1 (g5438), .I2 (g7610));
AN2X1 gate15325(.O (g9033), .I1 (g6643), .I2 (g567));
AN2X1 gate15326(.O (g9034), .I1 (g6751), .I2 (g1251));
AN2X1 gate15327(.O (g9047), .I1 (g6448), .I2 (g7616));
AN2X1 gate15328(.O (g9048), .I1 (g3338), .I2 (g489));
AN2X1 gate15329(.O (g9049), .I1 (g5473), .I2 (g7619));
AN2X1 gate15330(.O (g9056), .I1 (g6945), .I2 (g1253));
AN2X1 gate15331(.O (g9057), .I1 (g7053), .I2 (g1945));
AN2X1 gate15332(.O (g9061), .I1 (g3306), .I2 (g7623));
AN2X1 gate15333(.O (g9062), .I1 (g5438), .I2 (g7626));
AN2X1 gate15334(.O (g9063), .I1 (g5438), .I2 (g7629));
AN2X1 gate15335(.O (g9064), .I1 (g6713), .I2 (g7632));
AN2X1 gate15336(.O (g9065), .I1 (g3494), .I2 (g1176));
AN2X1 gate15337(.O (g9066), .I1 (g5512), .I2 (g7635));
AN2X1 gate15338(.O (g9073), .I1 (g7195), .I2 (g1947));
AN2X1 gate15339(.O (g9074), .I1 (g7303), .I2 (g2639));
AN2X1 gate15340(.O (g9075), .I1 (g6448), .I2 (g7643));
AN2X1 gate15341(.O (g9076), .I1 (g5438), .I2 (g7646));
AN2X1 gate15342(.O (g9077), .I1 (g6448), .I2 (g7649));
AN2X1 gate15343(.O (g9078), .I1 (g3462), .I2 (g7652));
AN2X1 gate15344(.O (g9079), .I1 (g5473), .I2 (g7655));
AN2X1 gate15345(.O (g9080), .I1 (g5473), .I2 (g7658));
AN2X1 gate15346(.O (g9081), .I1 (g7015), .I2 (g7661));
AN2X1 gate15347(.O (g9082), .I1 (g3650), .I2 (g1870));
AN2X1 gate15348(.O (g9083), .I1 (g5556), .I2 (g7664));
AN2X1 gate15349(.O (g9090), .I1 (g7391), .I2 (g2641));
AN2X1 gate15350(.O (g9091), .I1 (g3306), .I2 (g7670));
AN2X1 gate15351(.O (g9092), .I1 (g6448), .I2 (g7673));
AN2X1 gate15352(.O (g9093), .I1 (g3306), .I2 (g7676));
AN2X1 gate15353(.O (g9094), .I1 (g6713), .I2 (g7679));
AN2X1 gate15354(.O (g9095), .I1 (g5473), .I2 (g7682));
AN2X1 gate15355(.O (g9096), .I1 (g6713), .I2 (g7685));
AN2X1 gate15356(.O (g9097), .I1 (g3618), .I2 (g7688));
AN2X1 gate15357(.O (g9098), .I1 (g5512), .I2 (g7691));
AN2X1 gate15358(.O (g9099), .I1 (g5512), .I2 (g7694));
AN2X1 gate15359(.O (g9100), .I1 (g7265), .I2 (g7697));
AN2X1 gate15360(.O (g9101), .I1 (g3806), .I2 (g2564));
AN2X1 gate15361(.O (g9102), .I1 (g3306), .I2 (g7703));
AN2X1 gate15362(.O (g9103), .I1 (g3462), .I2 (g7706));
AN2X1 gate15363(.O (g9104), .I1 (g6713), .I2 (g7709));
AN2X1 gate15364(.O (g9105), .I1 (g3462), .I2 (g7712));
AN2X1 gate15365(.O (g9106), .I1 (g7015), .I2 (g7715));
AN2X1 gate15366(.O (g9107), .I1 (g5512), .I2 (g7718));
AN2X1 gate15367(.O (g9108), .I1 (g7015), .I2 (g7721));
AN2X1 gate15368(.O (g9109), .I1 (g3774), .I2 (g7724));
AN2X1 gate15369(.O (g9110), .I1 (g5556), .I2 (g7727));
AN2X1 gate15370(.O (g9111), .I1 (g5556), .I2 (g7730));
AN2X1 gate15371(.O (g9112), .I1 (g3462), .I2 (g7733));
AN2X1 gate15372(.O (g9113), .I1 (g3618), .I2 (g7736));
AN2X1 gate15373(.O (g9114), .I1 (g7015), .I2 (g7739));
AN2X1 gate15374(.O (g9115), .I1 (g3618), .I2 (g7742));
AN2X1 gate15375(.O (g9116), .I1 (g7265), .I2 (g7745));
AN2X1 gate15376(.O (g9117), .I1 (g5556), .I2 (g7748));
AN2X1 gate15377(.O (g9118), .I1 (g7265), .I2 (g7751));
AN2X1 gate15378(.O (g9119), .I1 (g5438), .I2 (g7754));
AN2X1 gate15379(.O (g9120), .I1 (g3618), .I2 (g7757));
AN2X1 gate15380(.O (g9121), .I1 (g3774), .I2 (g7760));
AN2X1 gate15381(.O (g9122), .I1 (g7265), .I2 (g7763));
AN2X1 gate15382(.O (g9123), .I1 (g3774), .I2 (g7766));
AN2X1 gate15383(.O (g9124), .I1 (g6448), .I2 (g7769));
AN2X1 gate15384(.O (g9125), .I1 (g5473), .I2 (g7776));
AN2X1 gate15385(.O (g9126), .I1 (g3774), .I2 (g7779));
AN2X1 gate15386(.O (g9127), .I1 (g3306), .I2 (g7782));
AN2X1 gate15387(.O (g9131), .I1 (g6713), .I2 (g7785));
AN2X1 gate15388(.O (g9132), .I1 (g5512), .I2 (g7792));
AN2X1 gate15389(.O (g9133), .I1 (g3462), .I2 (g7796));
AN2X1 gate15390(.O (g9137), .I1 (g7015), .I2 (g7799));
AN2X1 gate15391(.O (g9138), .I1 (g5556), .I2 (g7806));
AN2X1 gate15392(.O (g9139), .I1 (g3618), .I2 (g7809));
AN2X1 gate15393(.O (g9143), .I1 (g7265), .I2 (g7812));
AN2X1 gate15394(.O (g9145), .I1 (g3774), .I2 (g7823));
AN2X1 gate15395(.O (g9241), .I1 (g6232), .I2 (g7950));
AN2X1 gate15396(.O (g9301), .I1 (g6314), .I2 (g7990));
AN2X1 gate15397(.O (g9302), .I1 (g6232), .I2 (g7993));
AN2X1 gate15398(.O (g9319), .I1 (g6369), .I2 (g8001));
AN2X1 gate15399(.O (g9364), .I1 (g3254), .I2 (g8053));
AN2X1 gate15400(.O (g9365), .I1 (g6314), .I2 (g8056));
AN2X1 gate15401(.O (g9366), .I1 (g6232), .I2 (g8059));
AN2X1 gate15402(.O (g9367), .I1 (g6232), .I2 (g8062));
AN2X1 gate15403(.O (g9382), .I1 (g6519), .I2 (g8065));
AN2X1 gate15404(.O (g9383), .I1 (g6369), .I2 (g8068));
AN2X1 gate15405(.O (g9400), .I1 (g6574), .I2 (g8076));
AN2X1 gate15406(.O (g9438), .I1 (g3254), .I2 (g8123));
AN2X1 gate15407(.O (g9439), .I1 (g6314), .I2 (g8126));
AN2X1 gate15408(.O (g9440), .I1 (g6232), .I2 (g8129));
AN2X1 gate15409(.O (g9441), .I1 (g6314), .I2 (g8132));
AN2X1 gate15410(.O (g9442), .I1 (g6232), .I2 (g8135));
AN2X1 gate15411(.O (g9461), .I1 (g3410), .I2 (g8138));
AN2X1 gate15412(.O (g9462), .I1 (g6519), .I2 (g8141));
AN2X1 gate15413(.O (g9463), .I1 (g6369), .I2 (g8144));
AN2X1 gate15414(.O (g9464), .I1 (g6369), .I2 (g8147));
AN2X1 gate15415(.O (g9479), .I1 (g6783), .I2 (g8150));
AN2X1 gate15416(.O (g9480), .I1 (g6574), .I2 (g8153));
AN2X1 gate15417(.O (g9497), .I1 (g6838), .I2 (g8161));
AN2X1 gate15418(.O (g9518), .I1 (g3254), .I2 (g8191));
AN2X1 gate15419(.O (g9519), .I1 (g6314), .I2 (g8194));
AN2X1 gate15420(.O (g9520), .I1 (g6232), .I2 (g8197));
AN2X1 gate15421(.O (g9521), .I1 (g3254), .I2 (g8200));
AN2X1 gate15422(.O (g9522), .I1 (g6314), .I2 (g8203));
AN2X1 gate15423(.O (g9523), .I1 (g6232), .I2 (g8206));
AN3X1 gate15424(.O (g9534), .I1 (g7772), .I2 (g6135), .I3 (g538));
AN2X1 gate15425(.O (g9580), .I1 (g3410), .I2 (g8209));
AN2X1 gate15426(.O (g9581), .I1 (g6519), .I2 (g8212));
AN2X1 gate15427(.O (g9582), .I1 (g6369), .I2 (g8215));
AN2X1 gate15428(.O (g9583), .I1 (g6519), .I2 (g8218));
AN2X1 gate15429(.O (g9584), .I1 (g6369), .I2 (g8221));
AN2X1 gate15430(.O (g9603), .I1 (g3566), .I2 (g8224));
AN2X1 gate15431(.O (g9604), .I1 (g6783), .I2 (g8227));
AN2X1 gate15432(.O (g9605), .I1 (g6574), .I2 (g8230));
AN2X1 gate15433(.O (g9606), .I1 (g6574), .I2 (g8233));
AN2X1 gate15434(.O (g9621), .I1 (g7085), .I2 (g8236));
AN2X1 gate15435(.O (g9622), .I1 (g6838), .I2 (g8239));
AN2X1 gate15436(.O (g9630), .I1 (g3254), .I2 (g3922));
AN2X1 gate15437(.O (g9631), .I1 (g6314), .I2 (g3925));
AN2X1 gate15438(.O (g9632), .I1 (g6232), .I2 (g3928));
AN2X1 gate15439(.O (g9633), .I1 (g3254), .I2 (g3931));
AN2X1 gate15440(.O (g9634), .I1 (g6314), .I2 (g3934));
AN2X1 gate15441(.O (g9635), .I1 (g6232), .I2 (g3937));
AN4X1 gate15442(.O (I16735), .I1 (g5856), .I2 (g4338), .I3 (g4339), .I4 (g5141));
AN4X1 gate15443(.O (I16736), .I1 (g5713), .I2 (g5958), .I3 (g4735), .I4 (g4736));
AN2X1 gate15444(.O (g9636), .I1 (I16735), .I2 (I16736));
AN2X1 gate15445(.O (g9639), .I1 (g5438), .I2 (g408));
AN2X1 gate15446(.O (g9647), .I1 (g6678), .I2 (g3942));
AN2X1 gate15447(.O (g9648), .I1 (g6678), .I2 (g3945));
AN2X1 gate15448(.O (g9660), .I1 (g3410), .I2 (g3948));
AN2X1 gate15449(.O (g9661), .I1 (g6519), .I2 (g3951));
AN2X1 gate15450(.O (g9662), .I1 (g6369), .I2 (g3954));
AN2X1 gate15451(.O (g9663), .I1 (g3410), .I2 (g3957));
AN2X1 gate15452(.O (g9664), .I1 (g6519), .I2 (g3960));
AN2X1 gate15453(.O (g9665), .I1 (g6369), .I2 (g3963));
AN3X1 gate15454(.O (g9676), .I1 (g7788), .I2 (g6145), .I3 (g1224));
AN2X1 gate15455(.O (g9722), .I1 (g3566), .I2 (g3966));
AN2X1 gate15456(.O (g9723), .I1 (g6783), .I2 (g3969));
AN2X1 gate15457(.O (g9724), .I1 (g6574), .I2 (g3972));
AN2X1 gate15458(.O (g9725), .I1 (g6783), .I2 (g3975));
AN2X1 gate15459(.O (g9726), .I1 (g6574), .I2 (g3978));
AN2X1 gate15460(.O (g9745), .I1 (g3722), .I2 (g3981));
AN2X1 gate15461(.O (g9746), .I1 (g7085), .I2 (g3984));
AN2X1 gate15462(.O (g9747), .I1 (g6838), .I2 (g3987));
AN2X1 gate15463(.O (g9748), .I1 (g6838), .I2 (g3990));
AN2X1 gate15464(.O (g9759), .I1 (g3254), .I2 (g4000));
AN2X1 gate15465(.O (g9760), .I1 (g6314), .I2 (g4003));
AN2X1 gate15466(.O (g9761), .I1 (g6232), .I2 (g4006));
AN2X1 gate15467(.O (g9762), .I1 (g3254), .I2 (g4009));
AN2X1 gate15468(.O (g9763), .I1 (g6314), .I2 (g4012));
AN2X1 gate15469(.O (g9764), .I1 (g6448), .I2 (g411));
AN2X1 gate15470(.O (g9765), .I1 (g5438), .I2 (g417));
AN2X1 gate15471(.O (g9766), .I1 (g5438), .I2 (g4017));
AN2X1 gate15472(.O (g9773), .I1 (g6912), .I2 (g4020));
AN2X1 gate15473(.O (g9774), .I1 (g6678), .I2 (g4023));
AN2X1 gate15474(.O (g9775), .I1 (g6912), .I2 (g4026));
AN2X1 gate15475(.O (g9776), .I1 (g3410), .I2 (g4029));
AN2X1 gate15476(.O (g9777), .I1 (g6519), .I2 (g4032));
AN2X1 gate15477(.O (g9778), .I1 (g6369), .I2 (g4035));
AN2X1 gate15478(.O (g9779), .I1 (g3410), .I2 (g4038));
AN2X1 gate15479(.O (g9780), .I1 (g6519), .I2 (g4041));
AN2X1 gate15480(.O (g9781), .I1 (g6369), .I2 (g4044));
AN4X1 gate15481(.O (I16826), .I1 (g5903), .I2 (g4507), .I3 (g4508), .I4 (g5234));
AN4X1 gate15482(.O (I16827), .I1 (g5771), .I2 (g5987), .I3 (g4911), .I4 (g4912));
AN2X1 gate15483(.O (g9782), .I1 (I16826), .I2 (I16827));
AN2X1 gate15484(.O (g9785), .I1 (g5473), .I2 (g1095));
AN2X1 gate15485(.O (g9793), .I1 (g6980), .I2 (g4049));
AN2X1 gate15486(.O (g9794), .I1 (g6980), .I2 (g4052));
AN2X1 gate15487(.O (g9806), .I1 (g3566), .I2 (g4055));
AN2X1 gate15488(.O (g9807), .I1 (g6783), .I2 (g4058));
AN2X1 gate15489(.O (g9808), .I1 (g6574), .I2 (g4061));
AN2X1 gate15490(.O (g9809), .I1 (g3566), .I2 (g4064));
AN2X1 gate15491(.O (g9810), .I1 (g6783), .I2 (g4067));
AN2X1 gate15492(.O (g9811), .I1 (g6574), .I2 (g4070));
AN3X1 gate15493(.O (g9822), .I1 (g7802), .I2 (g6166), .I3 (g1918));
AN2X1 gate15494(.O (g9868), .I1 (g3722), .I2 (g4073));
AN2X1 gate15495(.O (g9869), .I1 (g7085), .I2 (g4076));
AN2X1 gate15496(.O (g9870), .I1 (g6838), .I2 (g4079));
AN2X1 gate15497(.O (g9871), .I1 (g7085), .I2 (g4082));
AN2X1 gate15498(.O (g9872), .I1 (g6838), .I2 (g4085));
AN2X1 gate15499(.O (g9887), .I1 (g6232), .I2 (g4095));
AN2X1 gate15500(.O (g9888), .I1 (g3254), .I2 (g4098));
AN2X1 gate15501(.O (g9889), .I1 (g6314), .I2 (g4101));
AN2X1 gate15502(.O (g9890), .I1 (g6232), .I2 (g4104));
AN2X1 gate15503(.O (g9891), .I1 (g3254), .I2 (g4107));
AN2X1 gate15504(.O (g9892), .I1 (g3306), .I2 (g414));
AN2X1 gate15505(.O (g9893), .I1 (g6448), .I2 (g420));
AN2X1 gate15506(.O (g9894), .I1 (g6448), .I2 (g4112));
AN2X1 gate15507(.O (g9901), .I1 (g3366), .I2 (g4115));
AN2X1 gate15508(.O (g9902), .I1 (g6912), .I2 (g4118));
AN2X1 gate15509(.O (g9903), .I1 (g6678), .I2 (g4121));
AN2X1 gate15510(.O (g9904), .I1 (g3366), .I2 (g4124));
AN2X1 gate15511(.O (g9905), .I1 (g3410), .I2 (g4127));
AN2X1 gate15512(.O (g9906), .I1 (g6519), .I2 (g4130));
AN2X1 gate15513(.O (g9907), .I1 (g6369), .I2 (g4133));
AN2X1 gate15514(.O (g9908), .I1 (g3410), .I2 (g4136));
AN2X1 gate15515(.O (g9909), .I1 (g6519), .I2 (g4139));
AN2X1 gate15516(.O (g9910), .I1 (g6713), .I2 (g1098));
AN2X1 gate15517(.O (g9911), .I1 (g5473), .I2 (g1104));
AN2X1 gate15518(.O (g9912), .I1 (g5473), .I2 (g4144));
AN2X1 gate15519(.O (g9919), .I1 (g7162), .I2 (g4147));
AN2X1 gate15520(.O (g9920), .I1 (g6980), .I2 (g4150));
AN2X1 gate15521(.O (g9921), .I1 (g7162), .I2 (g4153));
AN2X1 gate15522(.O (g9922), .I1 (g3566), .I2 (g4156));
AN2X1 gate15523(.O (g9923), .I1 (g6783), .I2 (g4159));
AN2X1 gate15524(.O (g9924), .I1 (g6574), .I2 (g4162));
AN2X1 gate15525(.O (g9925), .I1 (g3566), .I2 (g4165));
AN2X1 gate15526(.O (g9926), .I1 (g6783), .I2 (g4168));
AN2X1 gate15527(.O (g9927), .I1 (g6574), .I2 (g4171));
AN4X1 gate15528(.O (I16930), .I1 (g5942), .I2 (g4683), .I3 (g4684), .I4 (g5297));
AN4X1 gate15529(.O (I16931), .I1 (g5830), .I2 (g6024), .I3 (g5070), .I4 (g5071));
AN2X1 gate15530(.O (g9928), .I1 (I16930), .I2 (I16931));
AN2X1 gate15531(.O (g9931), .I1 (g5512), .I2 (g1789));
AN2X1 gate15532(.O (g9939), .I1 (g7230), .I2 (g4176));
AN2X1 gate15533(.O (g9940), .I1 (g7230), .I2 (g4179));
AN2X1 gate15534(.O (g9952), .I1 (g3722), .I2 (g4182));
AN2X1 gate15535(.O (g9953), .I1 (g7085), .I2 (g4185));
AN2X1 gate15536(.O (g9954), .I1 (g6838), .I2 (g4188));
AN2X1 gate15537(.O (g9955), .I1 (g3722), .I2 (g4191));
AN2X1 gate15538(.O (g9956), .I1 (g7085), .I2 (g4194));
AN2X1 gate15539(.O (g9957), .I1 (g6838), .I2 (g4197));
AN3X1 gate15540(.O (g9968), .I1 (g7815), .I2 (g6193), .I3 (g2612));
AN2X1 gate15541(.O (g10007), .I1 (g6314), .I2 (g4205));
AN2X1 gate15542(.O (g10008), .I1 (g6232), .I2 (g4208));
AN2X1 gate15543(.O (g10009), .I1 (g3254), .I2 (g4211));
AN2X1 gate15544(.O (g10010), .I1 (g6314), .I2 (g4214));
AN2X1 gate15545(.O (g10011), .I1 (g5438), .I2 (g4217));
AN2X1 gate15546(.O (g10012), .I1 (g3306), .I2 (g423));
AN2X1 gate15547(.O (g10013), .I1 (g3306), .I2 (g4221));
AN2X1 gate15548(.O (g10014), .I1 (g5438), .I2 (g429));
AN2X1 gate15549(.O (g10024), .I1 (g3398), .I2 (g6912));
AN2X1 gate15550(.O (g10035), .I1 (g3366), .I2 (g4225));
AN2X1 gate15551(.O (g10036), .I1 (g6912), .I2 (g4228));
AN2X1 gate15552(.O (g10037), .I1 (g6678), .I2 (g4231));
AN2X1 gate15553(.O (g10041), .I1 (g6369), .I2 (g4234));
AN2X1 gate15554(.O (g10042), .I1 (g3410), .I2 (g4237));
AN2X1 gate15555(.O (g10043), .I1 (g6519), .I2 (g4240));
AN2X1 gate15556(.O (g10044), .I1 (g6369), .I2 (g4243));
AN2X1 gate15557(.O (g10045), .I1 (g3410), .I2 (g4246));
AN2X1 gate15558(.O (g10046), .I1 (g3462), .I2 (g1101));
AN2X1 gate15559(.O (g10047), .I1 (g6713), .I2 (g1107));
AN2X1 gate15560(.O (g10048), .I1 (g6713), .I2 (g4251));
AN2X1 gate15561(.O (g10055), .I1 (g3522), .I2 (g4254));
AN2X1 gate15562(.O (g10056), .I1 (g7162), .I2 (g4257));
AN2X1 gate15563(.O (g10057), .I1 (g6980), .I2 (g4260));
AN2X1 gate15564(.O (g10058), .I1 (g3522), .I2 (g4263));
AN2X1 gate15565(.O (g10059), .I1 (g3566), .I2 (g4266));
AN2X1 gate15566(.O (g10060), .I1 (g6783), .I2 (g4269));
AN2X1 gate15567(.O (g10061), .I1 (g6574), .I2 (g4272));
AN2X1 gate15568(.O (g10062), .I1 (g3566), .I2 (g4275));
AN2X1 gate15569(.O (g10063), .I1 (g6783), .I2 (g4278));
AN2X1 gate15570(.O (g10064), .I1 (g7015), .I2 (g1792));
AN2X1 gate15571(.O (g10065), .I1 (g5512), .I2 (g1798));
AN2X1 gate15572(.O (g10066), .I1 (g5512), .I2 (g4283));
AN2X1 gate15573(.O (g10073), .I1 (g7358), .I2 (g4286));
AN2X1 gate15574(.O (g10074), .I1 (g7230), .I2 (g4289));
AN2X1 gate15575(.O (g10075), .I1 (g7358), .I2 (g4292));
AN2X1 gate15576(.O (g10076), .I1 (g3722), .I2 (g4295));
AN2X1 gate15577(.O (g10077), .I1 (g7085), .I2 (g4298));
AN2X1 gate15578(.O (g10078), .I1 (g6838), .I2 (g4301));
AN2X1 gate15579(.O (g10079), .I1 (g3722), .I2 (g4304));
AN2X1 gate15580(.O (g10080), .I1 (g7085), .I2 (g4307));
AN2X1 gate15581(.O (g10081), .I1 (g6838), .I2 (g4310));
AN4X1 gate15582(.O (I17042), .I1 (g5976), .I2 (g4860), .I3 (g4861), .I4 (g5334));
AN4X1 gate15583(.O (I17043), .I1 (g5886), .I2 (g6040), .I3 (g5199), .I4 (g5200));
AN2X1 gate15584(.O (g10082), .I1 (I17042), .I2 (I17043));
AN2X1 gate15585(.O (g10085), .I1 (g5556), .I2 (g2483));
AN2X1 gate15586(.O (g10093), .I1 (g7426), .I2 (g4315));
AN2X1 gate15587(.O (g10094), .I1 (g7426), .I2 (g4318));
AN2X1 gate15588(.O (g10101), .I1 (g3254), .I2 (g4329));
AN2X1 gate15589(.O (g10102), .I1 (g6314), .I2 (g4332));
AN2X1 gate15590(.O (g10103), .I1 (g3254), .I2 (g4335));
AN2X1 gate15591(.O (g10104), .I1 (g6448), .I2 (g4340));
AN2X1 gate15592(.O (g10105), .I1 (g5438), .I2 (g4343));
AN2X1 gate15593(.O (g10106), .I1 (g6448), .I2 (g432));
AN2X1 gate15594(.O (g10107), .I1 (g5438), .I2 (g438));
AN2X1 gate15595(.O (g10108), .I1 (g6486), .I2 (g569));
AN2X1 gate15596(.O (g10112), .I1 (g3366), .I2 (g4348));
AN2X1 gate15597(.O (g10113), .I1 (g6912), .I2 (g4351));
AN2X1 gate15598(.O (g10114), .I1 (g6678), .I2 (g4354));
AN2X1 gate15599(.O (g10115), .I1 (g6678), .I2 (g4357));
AN2X1 gate15600(.O (g10116), .I1 (g6519), .I2 (g4360));
AN2X1 gate15601(.O (g10117), .I1 (g6369), .I2 (g4363));
AN2X1 gate15602(.O (g10118), .I1 (g3410), .I2 (g4366));
AN2X1 gate15603(.O (g10119), .I1 (g6519), .I2 (g4369));
AN2X1 gate15604(.O (g10120), .I1 (g5473), .I2 (g4372));
AN2X1 gate15605(.O (g10121), .I1 (g3462), .I2 (g1110));
AN2X1 gate15606(.O (g10122), .I1 (g3462), .I2 (g4376));
AN2X1 gate15607(.O (g10123), .I1 (g5473), .I2 (g1116));
AN2X1 gate15608(.O (g10133), .I1 (g3554), .I2 (g7162));
AN2X1 gate15609(.O (g10144), .I1 (g3522), .I2 (g4380));
AN2X1 gate15610(.O (g10145), .I1 (g7162), .I2 (g4383));
AN2X1 gate15611(.O (g10146), .I1 (g6980), .I2 (g4386));
AN2X1 gate15612(.O (g10150), .I1 (g6574), .I2 (g4389));
AN2X1 gate15613(.O (g10151), .I1 (g3566), .I2 (g4392));
AN2X1 gate15614(.O (g10152), .I1 (g6783), .I2 (g4395));
AN2X1 gate15615(.O (g10153), .I1 (g6574), .I2 (g4398));
AN2X1 gate15616(.O (g10154), .I1 (g3566), .I2 (g4401));
AN2X1 gate15617(.O (g10155), .I1 (g3618), .I2 (g1795));
AN2X1 gate15618(.O (g10156), .I1 (g7015), .I2 (g1801));
AN2X1 gate15619(.O (g10157), .I1 (g7015), .I2 (g4406));
AN2X1 gate15620(.O (g10164), .I1 (g3678), .I2 (g4409));
AN2X1 gate15621(.O (g10165), .I1 (g7358), .I2 (g4412));
AN2X1 gate15622(.O (g10166), .I1 (g7230), .I2 (g4415));
AN2X1 gate15623(.O (g10167), .I1 (g3678), .I2 (g4418));
AN2X1 gate15624(.O (g10168), .I1 (g3722), .I2 (g4421));
AN2X1 gate15625(.O (g10169), .I1 (g7085), .I2 (g4424));
AN2X1 gate15626(.O (g10170), .I1 (g6838), .I2 (g4427));
AN2X1 gate15627(.O (g10171), .I1 (g3722), .I2 (g4430));
AN2X1 gate15628(.O (g10172), .I1 (g7085), .I2 (g4433));
AN2X1 gate15629(.O (g10173), .I1 (g7265), .I2 (g2486));
AN2X1 gate15630(.O (g10174), .I1 (g5556), .I2 (g2492));
AN2X1 gate15631(.O (g10175), .I1 (g5556), .I2 (g4438));
AN2X1 gate15632(.O (g10182), .I1 (g7488), .I2 (g4441));
AN2X1 gate15633(.O (g10183), .I1 (g7426), .I2 (g4444));
AN2X1 gate15634(.O (g10184), .I1 (g7488), .I2 (g4447));
AN4X1 gate15635(.O (I17156), .I1 (g6898), .I2 (g2998), .I3 (g6901), .I4 (g3002));
AN4X1 gate15636(.O (g10186), .I1 (g3013), .I2 (g7466), .I3 (g3024), .I4 (I17156));
AN2X1 gate15637(.O (g10192), .I1 (g3254), .I2 (g4453));
AN2X1 gate15638(.O (g10193), .I1 (g3306), .I2 (g4465));
AN2X1 gate15639(.O (g10194), .I1 (g6448), .I2 (g4468));
AN2X1 gate15640(.O (g10195), .I1 (g5438), .I2 (g4471));
AN2X1 gate15641(.O (g10196), .I1 (g3306), .I2 (g435));
AN2X1 gate15642(.O (g10197), .I1 (g6448), .I2 (g441));
AN2X1 gate15643(.O (g10198), .I1 (g6643), .I2 (g571));
AN2X1 gate15644(.O (g10199), .I1 (g6486), .I2 (g4476));
AN2X1 gate15645(.O (g10200), .I1 (g6486), .I2 (g587));
AN2X1 gate15646(.O (g10201), .I1 (g3366), .I2 (g4480));
AN2X1 gate15647(.O (g10202), .I1 (g6912), .I2 (g4483));
AN2X1 gate15648(.O (g10203), .I1 (g6678), .I2 (g4486));
AN2X1 gate15649(.O (g10204), .I1 (g6912), .I2 (g4489));
AN2X1 gate15650(.O (g10205), .I1 (g6678), .I2 (g4492));
AN2X1 gate15651(.O (g10206), .I1 (g3410), .I2 (g4498));
AN2X1 gate15652(.O (g10207), .I1 (g6519), .I2 (g4501));
AN2X1 gate15653(.O (g10208), .I1 (g3410), .I2 (g4504));
AN2X1 gate15654(.O (g10209), .I1 (g6713), .I2 (g4509));
AN2X1 gate15655(.O (g10210), .I1 (g5473), .I2 (g4512));
AN2X1 gate15656(.O (g10211), .I1 (g6713), .I2 (g1119));
AN2X1 gate15657(.O (g10212), .I1 (g5473), .I2 (g1125));
AN2X1 gate15658(.O (g10213), .I1 (g6751), .I2 (g1255));
AN2X1 gate15659(.O (g10217), .I1 (g3522), .I2 (g4517));
AN2X1 gate15660(.O (g10218), .I1 (g7162), .I2 (g4520));
AN2X1 gate15661(.O (g10219), .I1 (g6980), .I2 (g4523));
AN2X1 gate15662(.O (g10220), .I1 (g6980), .I2 (g4526));
AN2X1 gate15663(.O (g10221), .I1 (g6783), .I2 (g4529));
AN2X1 gate15664(.O (g10222), .I1 (g6574), .I2 (g4532));
AN2X1 gate15665(.O (g10223), .I1 (g3566), .I2 (g4535));
AN2X1 gate15666(.O (g10224), .I1 (g6783), .I2 (g4538));
AN2X1 gate15667(.O (g10225), .I1 (g5512), .I2 (g4541));
AN2X1 gate15668(.O (g10226), .I1 (g3618), .I2 (g1804));
AN2X1 gate15669(.O (g10227), .I1 (g3618), .I2 (g4545));
AN2X1 gate15670(.O (g10228), .I1 (g5512), .I2 (g1810));
AN2X1 gate15671(.O (g10238), .I1 (g3710), .I2 (g7358));
AN2X1 gate15672(.O (g10249), .I1 (g3678), .I2 (g4549));
AN2X1 gate15673(.O (g10250), .I1 (g7358), .I2 (g4552));
AN2X1 gate15674(.O (g10251), .I1 (g7230), .I2 (g4555));
AN2X1 gate15675(.O (g10255), .I1 (g6838), .I2 (g4558));
AN2X1 gate15676(.O (g10256), .I1 (g3722), .I2 (g4561));
AN2X1 gate15677(.O (g10257), .I1 (g7085), .I2 (g4564));
AN2X1 gate15678(.O (g10258), .I1 (g6838), .I2 (g4567));
AN2X1 gate15679(.O (g10259), .I1 (g3722), .I2 (g4570));
AN2X1 gate15680(.O (g10260), .I1 (g3774), .I2 (g2489));
AN2X1 gate15681(.O (g10261), .I1 (g7265), .I2 (g2495));
AN2X1 gate15682(.O (g10262), .I1 (g7265), .I2 (g4575));
AN2X1 gate15683(.O (g10269), .I1 (g3834), .I2 (g4578));
AN2X1 gate15684(.O (g10270), .I1 (g7488), .I2 (g4581));
AN2X1 gate15685(.O (g10271), .I1 (g7426), .I2 (g4584));
AN2X1 gate15686(.O (g10272), .I1 (g3834), .I2 (g4587));
AN2X1 gate15687(.O (g10279), .I1 (g3306), .I2 (g4592));
AN2X1 gate15688(.O (g10280), .I1 (g6448), .I2 (g4595));
AN2X1 gate15689(.O (g10281), .I1 (g5438), .I2 (g4598));
AN2X1 gate15690(.O (g10282), .I1 (g3306), .I2 (g444));
AN2X1 gate15691(.O (g10283), .I1 (g3338), .I2 (g573));
AN2X1 gate15692(.O (g10284), .I1 (g6643), .I2 (g4603));
AN2X1 gate15693(.O (g10285), .I1 (g6486), .I2 (g4606));
AN2X1 gate15694(.O (g10286), .I1 (g6643), .I2 (g590));
AN2X1 gate15695(.O (g10287), .I1 (g6486), .I2 (g596));
AN2X1 gate15696(.O (g10288), .I1 (g3366), .I2 (g4611));
AN2X1 gate15697(.O (g10289), .I1 (g6912), .I2 (g4614));
AN2X1 gate15698(.O (g10290), .I1 (g6678), .I2 (g4617));
AN2X1 gate15699(.O (g10291), .I1 (g3366), .I2 (g4620));
AN2X1 gate15700(.O (g10292), .I1 (g6912), .I2 (g4623));
AN2X1 gate15701(.O (g10293), .I1 (g6678), .I2 (g4626));
AN2X1 gate15702(.O (g10294), .I1 (g3410), .I2 (g4629));
AN2X1 gate15703(.O (g10295), .I1 (g3462), .I2 (g4641));
AN2X1 gate15704(.O (g10296), .I1 (g6713), .I2 (g4644));
AN2X1 gate15705(.O (g10297), .I1 (g5473), .I2 (g4647));
AN2X1 gate15706(.O (g10298), .I1 (g3462), .I2 (g1122));
AN2X1 gate15707(.O (g10299), .I1 (g6713), .I2 (g1128));
AN2X1 gate15708(.O (g10300), .I1 (g6945), .I2 (g1257));
AN2X1 gate15709(.O (g10301), .I1 (g6751), .I2 (g4652));
AN2X1 gate15710(.O (g10302), .I1 (g6751), .I2 (g1273));
AN2X1 gate15711(.O (g10303), .I1 (g3522), .I2 (g4656));
AN2X1 gate15712(.O (g10304), .I1 (g7162), .I2 (g4659));
AN2X1 gate15713(.O (g10305), .I1 (g6980), .I2 (g4662));
AN2X1 gate15714(.O (g10306), .I1 (g7162), .I2 (g4665));
AN2X1 gate15715(.O (g10307), .I1 (g6980), .I2 (g4668));
AN2X1 gate15716(.O (g10308), .I1 (g3566), .I2 (g4674));
AN2X1 gate15717(.O (g10309), .I1 (g6783), .I2 (g4677));
AN2X1 gate15718(.O (g10310), .I1 (g3566), .I2 (g4680));
AN2X1 gate15719(.O (g10311), .I1 (g7015), .I2 (g4685));
AN2X1 gate15720(.O (g10312), .I1 (g5512), .I2 (g4688));
AN2X1 gate15721(.O (g10313), .I1 (g7015), .I2 (g1813));
AN2X1 gate15722(.O (g10314), .I1 (g5512), .I2 (g1819));
AN2X1 gate15723(.O (g10315), .I1 (g7053), .I2 (g1949));
AN2X1 gate15724(.O (g10319), .I1 (g3678), .I2 (g4693));
AN2X1 gate15725(.O (g10320), .I1 (g7358), .I2 (g4696));
AN2X1 gate15726(.O (g10321), .I1 (g7230), .I2 (g4699));
AN2X1 gate15727(.O (g10322), .I1 (g7230), .I2 (g4702));
AN2X1 gate15728(.O (g10323), .I1 (g7085), .I2 (g4705));
AN2X1 gate15729(.O (g10324), .I1 (g6838), .I2 (g4708));
AN2X1 gate15730(.O (g10325), .I1 (g3722), .I2 (g4711));
AN2X1 gate15731(.O (g10326), .I1 (g7085), .I2 (g4714));
AN2X1 gate15732(.O (g10327), .I1 (g5556), .I2 (g4717));
AN2X1 gate15733(.O (g10328), .I1 (g3774), .I2 (g2498));
AN2X1 gate15734(.O (g10329), .I1 (g3774), .I2 (g4721));
AN2X1 gate15735(.O (g10330), .I1 (g5556), .I2 (g2504));
AN2X1 gate15736(.O (g10340), .I1 (g3866), .I2 (g7488));
AN2X1 gate15737(.O (g10351), .I1 (g3834), .I2 (g4725));
AN2X1 gate15738(.O (g10352), .I1 (g7488), .I2 (g4728));
AN2X1 gate15739(.O (g10353), .I1 (g7426), .I2 (g4731));
AN2X1 gate15740(.O (g10360), .I1 (g3306), .I2 (g4737));
AN2X1 gate15741(.O (g10361), .I1 (g6448), .I2 (g4740));
AN2X1 gate15742(.O (g10362), .I1 (g3338), .I2 (g4743));
AN2X1 gate15743(.O (g10363), .I1 (g6643), .I2 (g4746));
AN2X1 gate15744(.O (g10364), .I1 (g6486), .I2 (g4749));
AN2X1 gate15745(.O (g10365), .I1 (g3338), .I2 (g593));
AN2X1 gate15746(.O (g10366), .I1 (g6643), .I2 (g599));
AN2X1 gate15747(.O (g10367), .I1 (g3366), .I2 (g4754));
AN2X1 gate15748(.O (g10368), .I1 (g6912), .I2 (g4757));
AN2X1 gate15749(.O (g10369), .I1 (g6678), .I2 (g4760));
AN2X1 gate15750(.O (g10370), .I1 (g3366), .I2 (g4763));
AN2X1 gate15751(.O (g10371), .I1 (g6912), .I2 (g4766));
AN2X1 gate15752(.O (g10372), .I1 (g3462), .I2 (g4769));
AN2X1 gate15753(.O (g10373), .I1 (g6713), .I2 (g4772));
AN2X1 gate15754(.O (g10374), .I1 (g5473), .I2 (g4775));
AN2X1 gate15755(.O (g10375), .I1 (g3462), .I2 (g1131));
AN2X1 gate15756(.O (g10376), .I1 (g3494), .I2 (g1259));
AN2X1 gate15757(.O (g10377), .I1 (g6945), .I2 (g4780));
AN2X1 gate15758(.O (g10378), .I1 (g6751), .I2 (g4783));
AN2X1 gate15759(.O (g10379), .I1 (g6945), .I2 (g1276));
AN2X1 gate15760(.O (g10380), .I1 (g6751), .I2 (g1282));
AN2X1 gate15761(.O (g10381), .I1 (g3522), .I2 (g4788));
AN2X1 gate15762(.O (g10382), .I1 (g7162), .I2 (g4791));
AN2X1 gate15763(.O (g10383), .I1 (g6980), .I2 (g4794));
AN2X1 gate15764(.O (g10384), .I1 (g3522), .I2 (g4797));
AN2X1 gate15765(.O (g10385), .I1 (g7162), .I2 (g4800));
AN2X1 gate15766(.O (g10386), .I1 (g6980), .I2 (g4803));
AN2X1 gate15767(.O (g10387), .I1 (g3566), .I2 (g4806));
AN2X1 gate15768(.O (g10388), .I1 (g3618), .I2 (g4818));
AN2X1 gate15769(.O (g10389), .I1 (g7015), .I2 (g4821));
AN2X1 gate15770(.O (g10390), .I1 (g5512), .I2 (g4824));
AN2X1 gate15771(.O (g10391), .I1 (g3618), .I2 (g1816));
AN2X1 gate15772(.O (g10392), .I1 (g7015), .I2 (g1822));
AN2X1 gate15773(.O (g10393), .I1 (g7195), .I2 (g1951));
AN2X1 gate15774(.O (g10394), .I1 (g7053), .I2 (g4829));
AN2X1 gate15775(.O (g10395), .I1 (g7053), .I2 (g1967));
AN2X1 gate15776(.O (g10396), .I1 (g3678), .I2 (g4833));
AN2X1 gate15777(.O (g10397), .I1 (g7358), .I2 (g4836));
AN2X1 gate15778(.O (g10398), .I1 (g7230), .I2 (g4839));
AN2X1 gate15779(.O (g10399), .I1 (g7358), .I2 (g4842));
AN2X1 gate15780(.O (g10400), .I1 (g7230), .I2 (g4845));
AN2X1 gate15781(.O (g10401), .I1 (g3722), .I2 (g4851));
AN2X1 gate15782(.O (g10402), .I1 (g7085), .I2 (g4854));
AN2X1 gate15783(.O (g10403), .I1 (g3722), .I2 (g4857));
AN2X1 gate15784(.O (g10404), .I1 (g7265), .I2 (g4862));
AN2X1 gate15785(.O (g10405), .I1 (g5556), .I2 (g4865));
AN2X1 gate15786(.O (g10406), .I1 (g7265), .I2 (g2507));
AN2X1 gate15787(.O (g10407), .I1 (g5556), .I2 (g2513));
AN2X1 gate15788(.O (g10408), .I1 (g7303), .I2 (g2643));
AN2X1 gate15789(.O (g10412), .I1 (g3834), .I2 (g4870));
AN2X1 gate15790(.O (g10413), .I1 (g7488), .I2 (g4873));
AN2X1 gate15791(.O (g10414), .I1 (g7426), .I2 (g4876));
AN2X1 gate15792(.O (g10415), .I1 (g7426), .I2 (g4879));
AN2X1 gate15793(.O (g10422), .I1 (g3306), .I2 (g4882));
AN2X1 gate15794(.O (g10423), .I1 (g5438), .I2 (g4885));
AN2X1 gate15795(.O (g10430), .I1 (g3338), .I2 (g4888));
AN2X1 gate15796(.O (g10431), .I1 (g6643), .I2 (g4891));
AN2X1 gate15797(.O (g10432), .I1 (g6486), .I2 (g4894));
AN2X1 gate15798(.O (g10433), .I1 (g3338), .I2 (g602));
AN2X1 gate15799(.O (g10434), .I1 (g6486), .I2 (g605));
AN2X1 gate15800(.O (g10435), .I1 (g3366), .I2 (g4899));
AN2X1 gate15801(.O (g10436), .I1 (g6912), .I2 (g4902));
AN2X1 gate15802(.O (g10437), .I1 (g6678), .I2 (g4905));
AN2X1 gate15803(.O (g10438), .I1 (g3366), .I2 (g4908));
AN2X1 gate15804(.O (g10439), .I1 (g3462), .I2 (g4913));
AN2X1 gate15805(.O (g10440), .I1 (g6713), .I2 (g4916));
AN2X1 gate15806(.O (g10441), .I1 (g3494), .I2 (g4919));
AN2X1 gate15807(.O (g10442), .I1 (g6945), .I2 (g4922));
AN2X1 gate15808(.O (g10443), .I1 (g6751), .I2 (g4925));
AN2X1 gate15809(.O (g10444), .I1 (g3494), .I2 (g1279));
AN2X1 gate15810(.O (g10445), .I1 (g6945), .I2 (g1285));
AN2X1 gate15811(.O (g10446), .I1 (g3522), .I2 (g4930));
AN2X1 gate15812(.O (g10447), .I1 (g7162), .I2 (g4933));
AN2X1 gate15813(.O (g10448), .I1 (g6980), .I2 (g4936));
AN2X1 gate15814(.O (g10449), .I1 (g3522), .I2 (g4939));
AN2X1 gate15815(.O (g10450), .I1 (g7162), .I2 (g4942));
AN2X1 gate15816(.O (g10451), .I1 (g3618), .I2 (g4945));
AN2X1 gate15817(.O (g10452), .I1 (g7015), .I2 (g4948));
AN2X1 gate15818(.O (g10453), .I1 (g5512), .I2 (g4951));
AN2X1 gate15819(.O (g10454), .I1 (g3618), .I2 (g1825));
AN2X1 gate15820(.O (g10455), .I1 (g3650), .I2 (g1953));
AN2X1 gate15821(.O (g10456), .I1 (g7195), .I2 (g4956));
AN2X1 gate15822(.O (g10457), .I1 (g7053), .I2 (g4959));
AN2X1 gate15823(.O (g10458), .I1 (g7195), .I2 (g1970));
AN2X1 gate15824(.O (g10459), .I1 (g7053), .I2 (g1976));
AN2X1 gate15825(.O (g10460), .I1 (g3678), .I2 (g4964));
AN2X1 gate15826(.O (g10461), .I1 (g7358), .I2 (g4967));
AN2X1 gate15827(.O (g10462), .I1 (g7230), .I2 (g4970));
AN2X1 gate15828(.O (g10463), .I1 (g3678), .I2 (g4973));
AN2X1 gate15829(.O (g10464), .I1 (g7358), .I2 (g4976));
AN2X1 gate15830(.O (g10465), .I1 (g7230), .I2 (g4979));
AN2X1 gate15831(.O (g10466), .I1 (g3722), .I2 (g4982));
AN2X1 gate15832(.O (g10467), .I1 (g3774), .I2 (g4994));
AN2X1 gate15833(.O (g10468), .I1 (g7265), .I2 (g4997));
AN2X1 gate15834(.O (g10469), .I1 (g5556), .I2 (g5000));
AN2X1 gate15835(.O (g10470), .I1 (g3774), .I2 (g2510));
AN2X1 gate15836(.O (g10471), .I1 (g7265), .I2 (g2516));
AN2X1 gate15837(.O (g10472), .I1 (g7391), .I2 (g2645));
AN2X1 gate15838(.O (g10473), .I1 (g7303), .I2 (g5005));
AN2X1 gate15839(.O (g10474), .I1 (g7303), .I2 (g2661));
AN2X1 gate15840(.O (g10475), .I1 (g3834), .I2 (g5009));
AN2X1 gate15841(.O (g10476), .I1 (g7488), .I2 (g5012));
AN2X1 gate15842(.O (g10477), .I1 (g7426), .I2 (g5015));
AN2X1 gate15843(.O (g10478), .I1 (g7488), .I2 (g5018));
AN2X1 gate15844(.O (g10479), .I1 (g7426), .I2 (g5021));
AN3X1 gate15845(.O (I17429), .I1 (g6901), .I2 (g7338), .I3 (g7146));
AN3X1 gate15846(.O (g10480), .I1 (g7466), .I2 (g7342), .I3 (I17429));
AN2X1 gate15847(.O (g10485), .I1 (g6448), .I2 (g5024));
AN2X1 gate15848(.O (g10492), .I1 (g3338), .I2 (g5027));
AN2X1 gate15849(.O (g10493), .I1 (g6643), .I2 (g5030));
AN2X1 gate15850(.O (g10494), .I1 (g6643), .I2 (g608));
AN2X1 gate15851(.O (g10495), .I1 (g6486), .I2 (g614));
AN2X1 gate15852(.O (g10496), .I1 (g3366), .I2 (g5035));
AN2X1 gate15853(.O (g10497), .I1 (g6912), .I2 (g5038));
AN2X1 gate15854(.O (g10498), .I1 (g3462), .I2 (g5041));
AN2X1 gate15855(.O (g10499), .I1 (g5473), .I2 (g5044));
AN2X1 gate15856(.O (g10506), .I1 (g3494), .I2 (g5047));
AN2X1 gate15857(.O (g10507), .I1 (g6945), .I2 (g5050));
AN2X1 gate15858(.O (g10508), .I1 (g6751), .I2 (g5053));
AN2X1 gate15859(.O (g10509), .I1 (g3494), .I2 (g1288));
AN2X1 gate15860(.O (g10510), .I1 (g6751), .I2 (g1291));
AN2X1 gate15861(.O (g10511), .I1 (g3522), .I2 (g5058));
AN2X1 gate15862(.O (g10512), .I1 (g7162), .I2 (g5061));
AN2X1 gate15863(.O (g10513), .I1 (g6980), .I2 (g5064));
AN2X1 gate15864(.O (g10514), .I1 (g3522), .I2 (g5067));
AN2X1 gate15865(.O (g10515), .I1 (g3618), .I2 (g5072));
AN2X1 gate15866(.O (g10516), .I1 (g7015), .I2 (g5075));
AN2X1 gate15867(.O (g10517), .I1 (g3650), .I2 (g5078));
AN2X1 gate15868(.O (g10518), .I1 (g7195), .I2 (g5081));
AN2X1 gate15869(.O (g10519), .I1 (g7053), .I2 (g5084));
AN2X1 gate15870(.O (g10520), .I1 (g3650), .I2 (g1973));
AN2X1 gate15871(.O (g10521), .I1 (g7195), .I2 (g1979));
AN2X1 gate15872(.O (g10522), .I1 (g3678), .I2 (g5089));
AN2X1 gate15873(.O (g10523), .I1 (g7358), .I2 (g5092));
AN2X1 gate15874(.O (g10524), .I1 (g7230), .I2 (g5095));
AN2X1 gate15875(.O (g10525), .I1 (g3678), .I2 (g5098));
AN2X1 gate15876(.O (g10526), .I1 (g7358), .I2 (g5101));
AN2X1 gate15877(.O (g10527), .I1 (g3774), .I2 (g5104));
AN2X1 gate15878(.O (g10528), .I1 (g7265), .I2 (g5107));
AN2X1 gate15879(.O (g10529), .I1 (g5556), .I2 (g5110));
AN2X1 gate15880(.O (g10530), .I1 (g3774), .I2 (g2519));
AN2X1 gate15881(.O (g10531), .I1 (g3806), .I2 (g2647));
AN2X1 gate15882(.O (g10532), .I1 (g7391), .I2 (g5115));
AN2X1 gate15883(.O (g10533), .I1 (g7303), .I2 (g5118));
AN2X1 gate15884(.O (g10534), .I1 (g7391), .I2 (g2664));
AN2X1 gate15885(.O (g10535), .I1 (g7303), .I2 (g2670));
AN2X1 gate15886(.O (g10536), .I1 (g3834), .I2 (g5123));
AN2X1 gate15887(.O (g10537), .I1 (g7488), .I2 (g5126));
AN2X1 gate15888(.O (g10538), .I1 (g7426), .I2 (g5129));
AN2X1 gate15889(.O (g10539), .I1 (g3834), .I2 (g5132));
AN2X1 gate15890(.O (g10540), .I1 (g7488), .I2 (g5135));
AN2X1 gate15891(.O (g10541), .I1 (g7426), .I2 (g5138));
AN2X1 gate15892(.O (g10548), .I1 (g3306), .I2 (g5142));
AN2X1 gate15893(.O (g10555), .I1 (g3338), .I2 (g5145));
AN2X1 gate15894(.O (g10556), .I1 (g3338), .I2 (g611));
AN2X1 gate15895(.O (g10557), .I1 (g6643), .I2 (g617));
AN2X1 gate15896(.O (g10558), .I1 (g3366), .I2 (g5150));
AN2X1 gate15897(.O (g10559), .I1 (g6713), .I2 (g5153));
AN2X1 gate15898(.O (g10566), .I1 (g3494), .I2 (g5156));
AN2X1 gate15899(.O (g10567), .I1 (g6945), .I2 (g5159));
AN2X1 gate15900(.O (g10568), .I1 (g6945), .I2 (g1294));
AN2X1 gate15901(.O (g10569), .I1 (g6751), .I2 (g1300));
AN2X1 gate15902(.O (g10570), .I1 (g3522), .I2 (g5164));
AN2X1 gate15903(.O (g10571), .I1 (g7162), .I2 (g5167));
AN2X1 gate15904(.O (g10572), .I1 (g3618), .I2 (g5170));
AN2X1 gate15905(.O (g10573), .I1 (g5512), .I2 (g5173));
AN2X1 gate15906(.O (g10580), .I1 (g3650), .I2 (g5176));
AN2X1 gate15907(.O (g10581), .I1 (g7195), .I2 (g5179));
AN2X1 gate15908(.O (g10582), .I1 (g7053), .I2 (g5182));
AN2X1 gate15909(.O (g10583), .I1 (g3650), .I2 (g1982));
AN2X1 gate15910(.O (g10584), .I1 (g7053), .I2 (g1985));
AN2X1 gate15911(.O (g10585), .I1 (g3678), .I2 (g5187));
AN2X1 gate15912(.O (g10586), .I1 (g7358), .I2 (g5190));
AN2X1 gate15913(.O (g10587), .I1 (g7230), .I2 (g5193));
AN2X1 gate15914(.O (g10588), .I1 (g3678), .I2 (g5196));
AN2X1 gate15915(.O (g10589), .I1 (g3774), .I2 (g5201));
AN2X1 gate15916(.O (g10590), .I1 (g7265), .I2 (g5204));
AN2X1 gate15917(.O (g10591), .I1 (g3806), .I2 (g5207));
AN2X1 gate15918(.O (g10592), .I1 (g7391), .I2 (g5210));
AN2X1 gate15919(.O (g10593), .I1 (g7303), .I2 (g5213));
AN2X1 gate15920(.O (g10594), .I1 (g3806), .I2 (g2667));
AN2X1 gate15921(.O (g10595), .I1 (g7391), .I2 (g2673));
AN2X1 gate15922(.O (g10596), .I1 (g3834), .I2 (g5218));
AN2X1 gate15923(.O (g10597), .I1 (g7488), .I2 (g5221));
AN2X1 gate15924(.O (g10598), .I1 (g7426), .I2 (g5224));
AN2X1 gate15925(.O (g10599), .I1 (g3834), .I2 (g5227));
AN2X1 gate15926(.O (g10600), .I1 (g7488), .I2 (g5230));
AN2X1 gate15927(.O (g10604), .I1 (g3338), .I2 (g620));
AN2X1 gate15928(.O (g10605), .I1 (g3462), .I2 (g5235));
AN2X1 gate15929(.O (g10612), .I1 (g3494), .I2 (g5238));
AN2X1 gate15930(.O (g10613), .I1 (g3494), .I2 (g1297));
AN2X1 gate15931(.O (g10614), .I1 (g6945), .I2 (g1303));
AN2X1 gate15932(.O (g10615), .I1 (g3522), .I2 (g5243));
AN2X1 gate15933(.O (g10616), .I1 (g7015), .I2 (g5246));
AN2X1 gate15934(.O (g10623), .I1 (g3650), .I2 (g5249));
AN2X1 gate15935(.O (g10624), .I1 (g7195), .I2 (g5252));
AN2X1 gate15936(.O (g10625), .I1 (g7195), .I2 (g1988));
AN2X1 gate15937(.O (g10626), .I1 (g7053), .I2 (g1994));
AN2X1 gate15938(.O (g10627), .I1 (g3678), .I2 (g5257));
AN2X1 gate15939(.O (g10628), .I1 (g7358), .I2 (g5260));
AN2X1 gate15940(.O (g10629), .I1 (g3774), .I2 (g5263));
AN2X1 gate15941(.O (g10630), .I1 (g5556), .I2 (g5266));
AN2X1 gate15942(.O (g10637), .I1 (g3806), .I2 (g5269));
AN2X1 gate15943(.O (g10638), .I1 (g7391), .I2 (g5272));
AN2X1 gate15944(.O (g10639), .I1 (g7303), .I2 (g5275));
AN2X1 gate15945(.O (g10640), .I1 (g3806), .I2 (g2676));
AN2X1 gate15946(.O (g10641), .I1 (g7303), .I2 (g2679));
AN2X1 gate15947(.O (g10642), .I1 (g3834), .I2 (g5280));
AN2X1 gate15948(.O (g10643), .I1 (g7488), .I2 (g5283));
AN2X1 gate15949(.O (g10644), .I1 (g7426), .I2 (g5286));
AN2X1 gate15950(.O (g10645), .I1 (g3834), .I2 (g5289));
AN2X1 gate15951(.O (g10650), .I1 (g6678), .I2 (g5293));
AN2X1 gate15952(.O (g10651), .I1 (g3494), .I2 (g1306));
AN2X1 gate15953(.O (g10652), .I1 (g3618), .I2 (g5298));
AN2X1 gate15954(.O (g10659), .I1 (g3650), .I2 (g5301));
AN2X1 gate15955(.O (g10660), .I1 (g3650), .I2 (g1991));
AN2X1 gate15956(.O (g10661), .I1 (g7195), .I2 (g1997));
AN2X1 gate15957(.O (g10662), .I1 (g3678), .I2 (g5306));
AN2X1 gate15958(.O (g10663), .I1 (g7265), .I2 (g5309));
AN2X1 gate15959(.O (g10670), .I1 (g3806), .I2 (g5312));
AN2X1 gate15960(.O (g10671), .I1 (g7391), .I2 (g5315));
AN2X1 gate15961(.O (g10672), .I1 (g7391), .I2 (g2682));
AN2X1 gate15962(.O (g10673), .I1 (g7303), .I2 (g2688));
AN2X1 gate15963(.O (g10674), .I1 (g3834), .I2 (g5320));
AN2X1 gate15964(.O (g10675), .I1 (g7488), .I2 (g5323));
AN2X1 gate15965(.O (g10678), .I1 (g6912), .I2 (g5327));
AN2X1 gate15966(.O (g10680), .I1 (g6980), .I2 (g5330));
AN2X1 gate15967(.O (g10681), .I1 (g3650), .I2 (g2000));
AN2X1 gate15968(.O (g10682), .I1 (g3774), .I2 (g5335));
AN2X1 gate15969(.O (g10689), .I1 (g3806), .I2 (g5338));
AN2X1 gate15970(.O (g10690), .I1 (g3806), .I2 (g2685));
AN2X1 gate15971(.O (g10691), .I1 (g7391), .I2 (g2691));
AN2X1 gate15972(.O (g10692), .I1 (g3834), .I2 (g5343));
AN4X1 gate15973(.O (g10693), .I1 (g7462), .I2 (g7522), .I3 (g2924), .I4 (g7545));
AN2X1 gate15974(.O (g10704), .I1 (g3366), .I2 (g5352));
AN2X1 gate15975(.O (g10707), .I1 (g7162), .I2 (g5355));
AN2X1 gate15976(.O (g10709), .I1 (g7230), .I2 (g5358));
AN2X1 gate15977(.O (g10710), .I1 (g3806), .I2 (g2694));
AN3X1 gate15978(.O (I17599), .I1 (g7566), .I2 (g7583), .I3 (g7587));
AN3X1 gate15979(.O (g10711), .I1 (g7595), .I2 (g7600), .I3 (I17599));
AN2X1 gate15980(.O (g10724), .I1 (g3522), .I2 (g5369));
AN2X1 gate15981(.O (g10727), .I1 (g7358), .I2 (g5372));
AN2X1 gate15982(.O (g10729), .I1 (g7426), .I2 (g5375));
AN2X1 gate15983(.O (g10745), .I1 (g3678), .I2 (g5382));
AN2X1 gate15984(.O (g10748), .I1 (g7488), .I2 (g5385));
AN2X1 gate15985(.O (g10764), .I1 (g3834), .I2 (g5391));
AN2X1 gate15986(.O (g11347), .I1 (g6232), .I2 (g213));
AN2X1 gate15987(.O (g11420), .I1 (g6314), .I2 (g216));
AN2X1 gate15988(.O (g11421), .I1 (g6232), .I2 (g222));
AN2X1 gate15989(.O (g11431), .I1 (g6369), .I2 (g900));
AN2X1 gate15990(.O (g11607), .I1 (g5871), .I2 (g8360));
AN2X1 gate15991(.O (g11612), .I1 (g5881), .I2 (g8378));
AN2X1 gate15992(.O (g11637), .I1 (g5918), .I2 (g8427));
AN2X1 gate15993(.O (g11771), .I1 (g554), .I2 (g8622));
AN2X1 gate15994(.O (g11788), .I1 (g1240), .I2 (g8632));
AN2X1 gate15995(.O (g11805), .I1 (g6173), .I2 (g8643));
AN2X1 gate15996(.O (g11814), .I1 (g1934), .I2 (g8651));
AN2X1 gate15997(.O (g11816), .I1 (g7869), .I2 (g8655));
AN2X1 gate15998(.O (g11838), .I1 (g6205), .I2 (g8659));
AN2X1 gate15999(.O (g11847), .I1 (g2628), .I2 (g8667));
AN2X1 gate16000(.O (g11851), .I1 (g7849), .I2 (g8670));
AN2X1 gate16001(.O (g11880), .I1 (g6294), .I2 (g8678));
AN2X1 gate16002(.O (g11885), .I1 (g7834), .I2 (g8684));
AN2X1 gate16003(.O (g11922), .I1 (g6431), .I2 (g8690));
AN2X1 gate16004(.O (g11926), .I1 (g8169), .I2 (g8696));
AN2X1 gate16005(.O (g11966), .I1 (g8090), .I2 (g8708));
AN2X1 gate16006(.O (g11967), .I1 (g7967), .I2 (g8711));
AN2X1 gate16007(.O (g12012), .I1 (g8015), .I2 (g8745));
AN2X1 gate16008(.O (g12069), .I1 (g7964), .I2 (g8763));
AN2X1 gate16009(.O (g12070), .I1 (g8018), .I2 (g8766));
AN2X1 gate16010(.O (g12128), .I1 (g7916), .I2 (g8785));
AN2X1 gate16011(.O (g12129), .I1 (g7872), .I2 (g8788));
AN2X1 gate16012(.O (g12186), .I1 (g8093), .I2 (g8805));
AN2X1 gate16013(.O (g12273), .I1 (g8172), .I2 (g8829));
AN2X1 gate16014(.O (g12274), .I1 (g7900), .I2 (g8832));
AN2X1 gate16015(.O (g12307), .I1 (g7919), .I2 (g8853));
AN2X1 gate16016(.O (g12330), .I1 (g8246), .I2 (g8879));
AN2X1 gate16017(.O (g12331), .I1 (g7927), .I2 (g8882));
AN2X1 gate16018(.O (g12353), .I1 (g7852), .I2 (g8915));
AN2X1 gate16019(.O (g12376), .I1 (g7974), .I2 (g8949));
AN2X1 gate16020(.O (g12419), .I1 (g8028), .I2 (g9006));
AN2X1 gate16021(.O (g12429), .I1 (g8101), .I2 (g9044));
AN2X1 gate16022(.O (g12477), .I1 (g7822), .I2 (g9128));
AN2X1 gate16023(.O (g12494), .I1 (g7833), .I2 (g9134));
AN2X1 gate16024(.O (g12514), .I1 (g7848), .I2 (g9140));
AN2X1 gate16025(.O (g12531), .I1 (g7868), .I2 (g9146));
AN2X1 gate16026(.O (g12650), .I1 (g6149), .I2 (g9290));
AN4X1 gate16027(.O (I19937), .I1 (g9507), .I2 (g9427), .I3 (g9356), .I4 (g9293));
AN4X1 gate16028(.O (I19938), .I1 (g9232), .I2 (g9187), .I3 (g9161), .I4 (g9150));
AN2X1 gate16029(.O (g12876), .I1 (I19937), .I2 (I19938));
AN2X1 gate16030(.O (g12908), .I1 (g7899), .I2 (g10004));
AN4X1 gate16031(.O (I19971), .I1 (g9649), .I2 (g9569), .I3 (g9453), .I4 (g9374));
AN4X1 gate16032(.O (I19972), .I1 (g9310), .I2 (g9248), .I3 (g9203), .I4 (g9174));
AN2X1 gate16033(.O (g12916), .I1 (I19971), .I2 (I19972));
AN2X1 gate16034(.O (g12938), .I1 (g8179), .I2 (g10096));
AN4X1 gate16035(.O (I19996), .I1 (g9795), .I2 (g9711), .I3 (g9595), .I4 (g9471));
AN4X1 gate16036(.O (I19997), .I1 (g9391), .I2 (g9326), .I3 (g9264), .I4 (g9216));
AN2X1 gate16037(.O (g12945), .I1 (I19996), .I2 (I19997));
AN2X1 gate16038(.O (g12966), .I1 (g7926), .I2 (g10189));
AN4X1 gate16039(.O (I20021), .I1 (g9941), .I2 (g9857), .I3 (g9737), .I4 (g9613));
AN4X1 gate16040(.O (I20022), .I1 (g9488), .I2 (g9407), .I3 (g9342), .I4 (g9277));
AN2X1 gate16041(.O (g12974), .I1 (I20021), .I2 (I20022));
AN2X1 gate16042(.O (g12989), .I1 (g8254), .I2 (g10273));
AN2X1 gate16043(.O (g12990), .I1 (g8180), .I2 (g10276));
AN2X1 gate16044(.O (g13000), .I1 (g7973), .I2 (g10357));
AN2X1 gate16045(.O (g13004), .I1 (g10186), .I2 (g8317));
AN2X1 gate16046(.O (g13009), .I1 (g3995), .I2 (g10416));
AN2X1 gate16047(.O (g13010), .I1 (g8255), .I2 (g10419));
AN2X1 gate16048(.O (g13023), .I1 (g8027), .I2 (g10482));
AN2X1 gate16049(.O (g13031), .I1 (g7879), .I2 (g10542));
AN2X1 gate16050(.O (g13032), .I1 (g3996), .I2 (g10545));
AN2X1 gate16051(.O (g13042), .I1 (g8100), .I2 (g10601));
AN3X1 gate16052(.O (I20100), .I1 (g10186), .I2 (g3018), .I3 (g3028));
AN3X1 gate16053(.O (g13055), .I1 (g7471), .I2 (g7570), .I3 (I20100));
AN2X1 gate16054(.O (g13056), .I1 (g4092), .I2 (g10646));
AN4X1 gate16055(.O (I20131), .I1 (g8313), .I2 (g7542), .I3 (g2888), .I4 (g7566));
AN4X1 gate16056(.O (I20132), .I1 (g2892), .I2 (g2903), .I3 (g7595), .I4 (g2908));
AN2X1 gate16057(.O (g13082), .I1 (I20131), .I2 (I20132));
AN4X1 gate16058(.O (g13110), .I1 (g10693), .I2 (g2883), .I3 (g7562), .I4 (g10711));
AN2X1 gate16059(.O (g13247), .I1 (g298), .I2 (g11032));
AN2X1 gate16060(.O (g13266), .I1 (g5628), .I2 (g11088));
AN2X1 gate16061(.O (g13270), .I1 (g985), .I2 (g11102));
AN2X1 gate16062(.O (g13289), .I1 (g5647), .I2 (g11141));
AN2X1 gate16063(.O (g13291), .I1 (g5656), .I2 (g11154));
AN2X1 gate16064(.O (g13295), .I1 (g1679), .I2 (g11170));
AN2X1 gate16065(.O (g13316), .I1 (g5675), .I2 (g11210));
AN2X1 gate16066(.O (g13320), .I1 (g5685), .I2 (g11225));
AN2X1 gate16067(.O (g13322), .I1 (g5694), .I2 (g11240));
AN2X1 gate16068(.O (g13326), .I1 (g2373), .I2 (g11256));
AN2X1 gate16069(.O (g13335), .I1 (g5708), .I2 (g11278));
AN2X1 gate16070(.O (g13340), .I1 (g5727), .I2 (g11294));
AN2X1 gate16071(.O (g13343), .I1 (g5737), .I2 (g11309));
AN2X1 gate16072(.O (g13345), .I1 (g5746), .I2 (g11324));
AN2X1 gate16073(.O (g13355), .I1 (g5756), .I2 (g11355));
AN2X1 gate16074(.O (g13360), .I1 (g5766), .I2 (g11373));
AN2X1 gate16075(.O (g13365), .I1 (g5785), .I2 (g11389));
AN2X1 gate16076(.O (g13368), .I1 (g5795), .I2 (g11404));
AN2X1 gate16077(.O (g13385), .I1 (g5815), .I2 (g11441));
AN2X1 gate16078(.O (g13390), .I1 (g5825), .I2 (g11459));
AN2X1 gate16079(.O (g13395), .I1 (g5844), .I2 (g11475));
AN2X1 gate16080(.O (g13477), .I1 (g6016), .I2 (g12191));
AN2X1 gate16081(.O (g13479), .I1 (g6017), .I2 (g12196));
AN2X1 gate16082(.O (g13480), .I1 (g6018), .I2 (g12197));
AN2X1 gate16083(.O (g13481), .I1 (g5864), .I2 (g11603));
AN2X1 gate16084(.O (g13483), .I1 (g6020), .I2 (g12209));
AN2X1 gate16085(.O (g13484), .I1 (g6021), .I2 (g12210));
AN2X1 gate16086(.O (g13485), .I1 (g6022), .I2 (g12211));
AN2X1 gate16087(.O (g13486), .I1 (g6023), .I2 (g12212));
AN2X1 gate16088(.O (g13487), .I1 (g5874), .I2 (g11608));
AN2X1 gate16089(.O (g13488), .I1 (g6025), .I2 (g12218));
AN2X1 gate16090(.O (g13489), .I1 (g6026), .I2 (g12219));
AN2X1 gate16091(.O (g13490), .I1 (g6027), .I2 (g12220));
AN2X1 gate16092(.O (g13491), .I1 (g6028), .I2 (g12221));
AN2X1 gate16093(.O (g13492), .I1 (g2371), .I2 (g12222));
AN2X1 gate16094(.O (g13493), .I1 (g5887), .I2 (g11613));
AN2X1 gate16095(.O (g13496), .I1 (g6032), .I2 (g12246));
AN2X1 gate16096(.O (g13498), .I1 (g6033), .I2 (g12251));
AN2X1 gate16097(.O (g13499), .I1 (g6034), .I2 (g12252));
AN2X1 gate16098(.O (g13500), .I1 (g5911), .I2 (g11633));
AN2X1 gate16099(.O (g13502), .I1 (g6036), .I2 (g12264));
AN2X1 gate16100(.O (g13503), .I1 (g6037), .I2 (g12265));
AN2X1 gate16101(.O (g13504), .I1 (g6038), .I2 (g12266));
AN2X1 gate16102(.O (g13505), .I1 (g6039), .I2 (g12267));
AN2X1 gate16103(.O (g13506), .I1 (g5921), .I2 (g11638));
AN2X1 gate16104(.O (g13513), .I1 (g6043), .I2 (g12289));
AN2X1 gate16105(.O (g13515), .I1 (g6044), .I2 (g12294));
AN2X1 gate16106(.O (g13516), .I1 (g6045), .I2 (g12295));
AN2X1 gate16107(.O (g13517), .I1 (g5950), .I2 (g11656));
AN2X1 gate16108(.O (g13527), .I1 (g6047), .I2 (g12325));
AN2X1 gate16109(.O (g13609), .I1 (g6141), .I2 (g12456));
AN2X1 gate16110(.O (g13619), .I1 (g6162), .I2 (g12466));
AN2X1 gate16111(.O (g13623), .I1 (g5428), .I2 (g12472));
AN2X1 gate16112(.O (g13625), .I1 (g6173), .I2 (g12476));
AN2X1 gate16113(.O (g13631), .I1 (g6189), .I2 (g12481));
AN2X1 gate16114(.O (g13634), .I1 (g12776), .I2 (g8617));
AN2X1 gate16115(.O (g13636), .I1 (g6205), .I2 (g12493));
AN2X1 gate16116(.O (g13642), .I1 (g6221), .I2 (g12498));
AN2X1 gate16117(.O (g13643), .I1 (g5431), .I2 (g12502));
AN2X1 gate16118(.O (g13645), .I1 (g6281), .I2 (g12504));
AN2X1 gate16119(.O (g13646), .I1 (g7772), .I2 (g12505));
AN2X1 gate16120(.O (g13648), .I1 (g6294), .I2 (g12513));
AN2X1 gate16121(.O (g13654), .I1 (g8093), .I2 (g11791));
AN2X1 gate16122(.O (g13655), .I1 (g7540), .I2 (g12518));
AN2X1 gate16123(.O (g13656), .I1 (g12776), .I2 (g8640));
AN2X1 gate16124(.O (g13671), .I1 (g6418), .I2 (g12521));
AN2X1 gate16125(.O (g13672), .I1 (g7788), .I2 (g12522));
AN2X1 gate16126(.O (g13674), .I1 (g6431), .I2 (g12530));
AN2X1 gate16127(.O (g13675), .I1 (g7561), .I2 (g12532));
AN2X1 gate16128(.O (g13676), .I1 (g5434), .I2 (g12533));
AN2X1 gate16129(.O (g13701), .I1 (g6623), .I2 (g12536));
AN2X1 gate16130(.O (g13702), .I1 (g7802), .I2 (g12537));
AN2X1 gate16131(.O (g13703), .I1 (g8018), .I2 (g11848));
AN2X1 gate16132(.O (g13704), .I1 (g7581), .I2 (g12542));
AN2X1 gate16133(.O (g13705), .I1 (g12776), .I2 (g8673));
AN2X1 gate16134(.O (g13738), .I1 (g6887), .I2 (g12545));
AN2X1 gate16135(.O (g13739), .I1 (g7815), .I2 (g12546));
AN2X1 gate16136(.O (g13740), .I1 (g6636), .I2 (g12547));
AN2X1 gate16137(.O (g13755), .I1 (g7347), .I2 (g12551));
AN2X1 gate16138(.O (g13787), .I1 (g7967), .I2 (g11923));
AN2X1 gate16139(.O (g13788), .I1 (g6897), .I2 (g12553));
AN2X1 gate16140(.O (g13789), .I1 (g7140), .I2 (g12554));
AN2X1 gate16141(.O (g13790), .I1 (g7475), .I2 (g12558));
AN2X1 gate16142(.O (g13796), .I1 (g7477), .I2 (g12559));
AN2X1 gate16143(.O (g13815), .I1 (g7139), .I2 (g12560));
AN2X1 gate16144(.O (g13816), .I1 (g7530), .I2 (g12596));
AN2X1 gate16145(.O (g13818), .I1 (g7531), .I2 (g12597));
AN2X1 gate16146(.O (g13824), .I1 (g7533), .I2 (g12598));
AN2X1 gate16147(.O (g13833), .I1 (g7919), .I2 (g12009));
AN2X1 gate16148(.O (g13834), .I1 (g7336), .I2 (g12599));
AN2X1 gate16149(.O (g13835), .I1 (g7461), .I2 (g12600));
AN2X1 gate16150(.O (g13837), .I1 (g7556), .I2 (g12642));
AN2X1 gate16151(.O (g13839), .I1 (g7557), .I2 (g12643));
AN2X1 gate16152(.O (g13845), .I1 (g7559), .I2 (g12644));
AN2X1 gate16153(.O (g13846), .I1 (g7460), .I2 (g12645));
AN2X1 gate16154(.O (g13847), .I1 (g7521), .I2 (g12646));
AN2X1 gate16155(.O (g13851), .I1 (g7579), .I2 (g12688));
AN2X1 gate16156(.O (g13853), .I1 (g7580), .I2 (g12689));
AN2X1 gate16157(.O (g13854), .I1 (g5349), .I2 (g12690));
AN2X1 gate16158(.O (g13855), .I1 (g7541), .I2 (g12691));
AN2X1 gate16159(.O (g13860), .I1 (g7593), .I2 (g12742));
AN2X1 gate16160(.O (g13862), .I1 (g5366), .I2 (g12743));
AN2X1 gate16161(.O (g13865), .I1 (g548), .I2 (g12748));
AN2X1 gate16162(.O (g13870), .I1 (g7582), .I2 (g12768));
AN2X1 gate16163(.O (g13871), .I1 (g7898), .I2 (g12775));
AN2X1 gate16164(.O (g13878), .I1 (g7610), .I2 (g12782));
AN2X1 gate16165(.O (g13880), .I1 (g1234), .I2 (g12790));
AN2X1 gate16166(.O (g13884), .I1 (g7594), .I2 (g12807));
AN2X1 gate16167(.O (g13892), .I1 (g7616), .I2 (g12815));
AN2X1 gate16168(.O (g13900), .I1 (g7619), .I2 (g12821));
AN2X1 gate16169(.O (g13902), .I1 (g1928), .I2 (g12829));
AN2X1 gate16170(.O (g13904), .I1 (g7337), .I2 (g12843));
AN2X1 gate16171(.O (g13905), .I1 (g7925), .I2 (g12847));
AN2X1 gate16172(.O (g13913), .I1 (g7623), .I2 (g12850));
AN2X1 gate16173(.O (g13914), .I1 (g7626), .I2 (g12851));
AN2X1 gate16174(.O (g13933), .I1 (g7632), .I2 (g12853));
AN2X1 gate16175(.O (g13941), .I1 (g7635), .I2 (g12859));
AN2X1 gate16176(.O (g13943), .I1 (g2622), .I2 (g12867));
AN2X1 gate16177(.O (g13944), .I1 (g7141), .I2 (g12874));
AN2X1 gate16178(.O (g13952), .I1 (g7643), .I2 (g12881));
AN2X1 gate16179(.O (g13953), .I1 (g7646), .I2 (g12882));
AN2X1 gate16180(.O (g13969), .I1 (g7652), .I2 (g12891));
AN2X1 gate16181(.O (g13970), .I1 (g7655), .I2 (g12892));
AN2X1 gate16182(.O (g13989), .I1 (g7661), .I2 (g12894));
AN2X1 gate16183(.O (g13997), .I1 (g7664), .I2 (g12900));
AN2X1 gate16184(.O (g13998), .I1 (g7972), .I2 (g12907));
AN2X1 gate16185(.O (g14006), .I1 (g7670), .I2 (g12914));
AN2X1 gate16186(.O (g14007), .I1 (g7673), .I2 (g12915));
AN2X1 gate16187(.O (g14022), .I1 (g7679), .I2 (g12921));
AN2X1 gate16188(.O (g14023), .I1 (g7682), .I2 (g12922));
AN2X1 gate16189(.O (g14039), .I1 (g7688), .I2 (g12931));
AN2X1 gate16190(.O (g14040), .I1 (g7691), .I2 (g12932));
AN2X1 gate16191(.O (g14059), .I1 (g7697), .I2 (g12934));
AN2X1 gate16192(.O (g14067), .I1 (g7703), .I2 (g12940));
AN2X1 gate16193(.O (g14097), .I1 (g7706), .I2 (g12943));
AN2X1 gate16194(.O (g14098), .I1 (g7709), .I2 (g12944));
AN2X1 gate16195(.O (g14113), .I1 (g7715), .I2 (g12950));
AN2X1 gate16196(.O (g14114), .I1 (g7718), .I2 (g12951));
AN2X1 gate16197(.O (g14130), .I1 (g7724), .I2 (g12960));
AN2X1 gate16198(.O (g14131), .I1 (g7727), .I2 (g12961));
AN2X1 gate16199(.O (g14143), .I1 (g8026), .I2 (g12965));
AN2X1 gate16200(.O (g14182), .I1 (g7733), .I2 (g12969));
AN2X1 gate16201(.O (g14212), .I1 (g7736), .I2 (g12972));
AN2X1 gate16202(.O (g14213), .I1 (g7739), .I2 (g12973));
AN2X1 gate16203(.O (g14228), .I1 (g7745), .I2 (g12979));
AN2X1 gate16204(.O (g14229), .I1 (g7748), .I2 (g12980));
AN2X1 gate16205(.O (g14297), .I1 (g7757), .I2 (g12993));
AN2X1 gate16206(.O (g14327), .I1 (g7760), .I2 (g12996));
AN2X1 gate16207(.O (g14328), .I1 (g7763), .I2 (g12997));
AN2X1 gate16208(.O (g14336), .I1 (g8099), .I2 (g12998));
AN2X1 gate16209(.O (g14419), .I1 (g7779), .I2 (g13003));
AN2X1 gate16210(.O (g14690), .I1 (g7841), .I2 (g13101));
AN2X1 gate16211(.O (g14724), .I1 (g7861), .I2 (g13117));
AN2X1 gate16212(.O (g14752), .I1 (g7891), .I2 (g13130));
AN2X1 gate16213(.O (g14767), .I1 (g13245), .I2 (g10765));
AN2X1 gate16214(.O (g14773), .I1 (g7915), .I2 (g13141));
AN2X1 gate16215(.O (g14884), .I1 (g8169), .I2 (g12548));
AN2X1 gate16216(.O (g14894), .I1 (g3940), .I2 (g13148));
AN2X1 gate16217(.O (g14956), .I1 (g11059), .I2 (g13151));
AN2X1 gate16218(.O (g14957), .I1 (g4015), .I2 (g13152));
AN2X1 gate16219(.O (g14958), .I1 (g4016), .I2 (g13153));
AN2X1 gate16220(.O (g14975), .I1 (g4047), .I2 (g13154));
AN2X1 gate16221(.O (g15020), .I1 (g8090), .I2 (g12561));
AN2X1 gate16222(.O (g15030), .I1 (g4110), .I2 (g13158));
AN2X1 gate16223(.O (g15031), .I1 (g4111), .I2 (g13159));
AN2X1 gate16224(.O (g15046), .I1 (g4142), .I2 (g13161));
AN2X1 gate16225(.O (g15047), .I1 (g4143), .I2 (g13162));
AN2X1 gate16226(.O (g15064), .I1 (g4174), .I2 (g13163));
AN2X1 gate16227(.O (g15093), .I1 (g7869), .I2 (g12601));
AN2X1 gate16228(.O (g15094), .I1 (g7872), .I2 (g12604));
AN2X1 gate16229(.O (g15104), .I1 (g4220), .I2 (g13167));
AN2X1 gate16230(.O (g15105), .I1 (g4224), .I2 (g13168));
AN2X1 gate16231(.O (g15126), .I1 (g4249), .I2 (g13169));
AN2X1 gate16232(.O (g15127), .I1 (g4250), .I2 (g13170));
AN2X1 gate16233(.O (g15142), .I1 (g4281), .I2 (g13172));
AN2X1 gate16234(.O (g15143), .I1 (g4282), .I2 (g13173));
AN2X1 gate16235(.O (g15160), .I1 (g4313), .I2 (g13174));
AN2X1 gate16236(.O (g15171), .I1 (g8015), .I2 (g12647));
AN2X1 gate16237(.O (g15172), .I1 (g4346), .I2 (g13176));
AN2X1 gate16238(.O (g15173), .I1 (g4347), .I2 (g13177));
AN2X1 gate16239(.O (g15178), .I1 (g640), .I2 (g12651));
AN2X1 gate16240(.O (g15196), .I1 (g4375), .I2 (g13178));
AN2X1 gate16241(.O (g15197), .I1 (g4379), .I2 (g13179));
AN2X1 gate16242(.O (g15218), .I1 (g4404), .I2 (g13180));
AN2X1 gate16243(.O (g15219), .I1 (g4405), .I2 (g13181));
AN2X1 gate16244(.O (g15234), .I1 (g4436), .I2 (g13183));
AN2X1 gate16245(.O (g15235), .I1 (g4437), .I2 (g13184));
AN2X1 gate16246(.O (g15243), .I1 (g7849), .I2 (g12692));
AN2X1 gate16247(.O (g15244), .I1 (g7852), .I2 (g12695));
AN2X1 gate16248(.O (g15245), .I1 (g4474), .I2 (g13185));
AN2X1 gate16249(.O (g15246), .I1 (g4475), .I2 (g13186));
AN2X1 gate16250(.O (g15247), .I1 (g4479), .I2 (g13187));
AN2X1 gate16251(.O (g15257), .I1 (g4357), .I2 (g12702));
AN2X1 gate16252(.O (g15258), .I1 (g4515), .I2 (g13188));
AN2X1 gate16253(.O (g15259), .I1 (g4516), .I2 (g13189));
AN2X1 gate16254(.O (g15264), .I1 (g1326), .I2 (g12705));
AN2X1 gate16255(.O (g15282), .I1 (g4544), .I2 (g13190));
AN2X1 gate16256(.O (g15283), .I1 (g4548), .I2 (g13191));
AN2X1 gate16257(.O (g15304), .I1 (g4573), .I2 (g13192));
AN2X1 gate16258(.O (g15305), .I1 (g4574), .I2 (g13193));
AN2X1 gate16259(.O (g15320), .I1 (g7964), .I2 (g12744));
AN2X1 gate16260(.O (g15321), .I1 (g4601), .I2 (g13195));
AN2X1 gate16261(.O (g15324), .I1 (g4609), .I2 (g13196));
AN2X1 gate16262(.O (g15325), .I1 (g4610), .I2 (g13197));
AN2X1 gate16263(.O (g15335), .I1 (g4489), .I2 (g12749));
AN2X1 gate16264(.O (g15336), .I1 (g4492), .I2 (g12752));
AN2X1 gate16265(.O (g15337), .I1 (g4650), .I2 (g13198));
AN2X1 gate16266(.O (g15338), .I1 (g4651), .I2 (g13199));
AN2X1 gate16267(.O (g15339), .I1 (g4655), .I2 (g13200));
AN2X1 gate16268(.O (g15349), .I1 (g4526), .I2 (g12759));
AN2X1 gate16269(.O (g15350), .I1 (g4691), .I2 (g13201));
AN2X1 gate16270(.O (g15351), .I1 (g4692), .I2 (g13202));
AN2X1 gate16271(.O (g15356), .I1 (g2020), .I2 (g12762));
AN2X1 gate16272(.O (g15374), .I1 (g4720), .I2 (g13203));
AN2X1 gate16273(.O (g15375), .I1 (g4724), .I2 (g13204));
AN2X1 gate16274(.O (g15388), .I1 (g7834), .I2 (g12769));
AN2X1 gate16275(.O (g15389), .I1 (g8246), .I2 (g12772));
AN2X1 gate16276(.O (g15391), .I1 (g4752), .I2 (g13205));
AN2X1 gate16277(.O (g15392), .I1 (g4753), .I2 (g13206));
AN2X1 gate16278(.O (g15402), .I1 (g4620), .I2 (g12783));
AN2X1 gate16279(.O (g15403), .I1 (g4623), .I2 (g12786));
AN2X1 gate16280(.O (g15407), .I1 (g4778), .I2 (g13207));
AN2X1 gate16281(.O (g15410), .I1 (g4786), .I2 (g13208));
AN2X1 gate16282(.O (g15411), .I1 (g4787), .I2 (g13209));
AN2X1 gate16283(.O (g15421), .I1 (g4665), .I2 (g12791));
AN2X1 gate16284(.O (g15422), .I1 (g4668), .I2 (g12794));
AN2X1 gate16285(.O (g15423), .I1 (g4827), .I2 (g13210));
AN2X1 gate16286(.O (g15424), .I1 (g4828), .I2 (g13211));
AN2X1 gate16287(.O (g15425), .I1 (g4832), .I2 (g13212));
AN2X1 gate16288(.O (g15435), .I1 (g4702), .I2 (g12801));
AN2X1 gate16289(.O (g15436), .I1 (g4868), .I2 (g13213));
AN2X1 gate16290(.O (g15437), .I1 (g4869), .I2 (g13214));
AN2X1 gate16291(.O (g15442), .I1 (g2714), .I2 (g12804));
AN2X1 gate16292(.O (g15452), .I1 (g7916), .I2 (g12808));
AN2X1 gate16293(.O (g15453), .I1 (g6898), .I2 (g12811));
AN2X1 gate16294(.O (g15459), .I1 (g4897), .I2 (g13218));
AN2X1 gate16295(.O (g15460), .I1 (g4898), .I2 (g13219));
AN2X1 gate16296(.O (g15470), .I1 (g4763), .I2 (g12816));
AN2X1 gate16297(.O (g15475), .I1 (g4928), .I2 (g13220));
AN2X1 gate16298(.O (g15476), .I1 (g4929), .I2 (g13221));
AN2X1 gate16299(.O (g15486), .I1 (g4797), .I2 (g12822));
AN2X1 gate16300(.O (g15487), .I1 (g4800), .I2 (g12825));
AN2X1 gate16301(.O (g15491), .I1 (g4954), .I2 (g13222));
AN2X1 gate16302(.O (g15494), .I1 (g4962), .I2 (g13223));
AN2X1 gate16303(.O (g15495), .I1 (g4963), .I2 (g13224));
AN2X1 gate16304(.O (g15505), .I1 (g4842), .I2 (g12830));
AN2X1 gate16305(.O (g15506), .I1 (g4845), .I2 (g12833));
AN2X1 gate16306(.O (g15507), .I1 (g5003), .I2 (g13225));
AN2X1 gate16307(.O (g15508), .I1 (g5004), .I2 (g13226));
AN2X1 gate16308(.O (g15509), .I1 (g5008), .I2 (g13227));
AN2X1 gate16309(.O (g15519), .I1 (g4879), .I2 (g12840));
AN2X1 gate16310(.O (g15520), .I1 (g8172), .I2 (g12844));
AN2X1 gate16311(.O (g15526), .I1 (g5033), .I2 (g13232));
AN2X1 gate16312(.O (g15527), .I1 (g5034), .I2 (g13233));
AN2X1 gate16313(.O (g15545), .I1 (g5056), .I2 (g13237));
AN2X1 gate16314(.O (g15546), .I1 (g5057), .I2 (g13238));
AN2X1 gate16315(.O (g15556), .I1 (g4939), .I2 (g12854));
AN2X1 gate16316(.O (g15561), .I1 (g5087), .I2 (g13239));
AN2X1 gate16317(.O (g15562), .I1 (g5088), .I2 (g13240));
AN2X1 gate16318(.O (g15572), .I1 (g4973), .I2 (g12860));
AN2X1 gate16319(.O (g15573), .I1 (g4976), .I2 (g12863));
AN2X1 gate16320(.O (g15577), .I1 (g5113), .I2 (g13241));
AN2X1 gate16321(.O (g15580), .I1 (g5121), .I2 (g13242));
AN2X1 gate16322(.O (g15581), .I1 (g5122), .I2 (g13243));
AN2X1 gate16323(.O (g15591), .I1 (g5018), .I2 (g12868));
AN2X1 gate16324(.O (g15592), .I1 (g5021), .I2 (g12871));
AN2X1 gate16325(.O (g15593), .I1 (g7897), .I2 (g13244));
AN2X1 gate16326(.O (g15594), .I1 (g5148), .I2 (g13249));
AN2X1 gate16327(.O (g15595), .I1 (g5149), .I2 (g13250));
AN2X1 gate16328(.O (g15604), .I1 (g5162), .I2 (g13255));
AN2X1 gate16329(.O (g15605), .I1 (g5163), .I2 (g13256));
AN2X1 gate16330(.O (g15623), .I1 (g5185), .I2 (g13260));
AN2X1 gate16331(.O (g15624), .I1 (g5186), .I2 (g13261));
AN2X1 gate16332(.O (g15634), .I1 (g5098), .I2 (g12895));
AN2X1 gate16333(.O (g15639), .I1 (g5216), .I2 (g13262));
AN2X1 gate16334(.O (g15640), .I1 (g5217), .I2 (g13263));
AN2X1 gate16335(.O (g15650), .I1 (g5132), .I2 (g12901));
AN2X1 gate16336(.O (g15651), .I1 (g5135), .I2 (g12904));
AN2X1 gate16337(.O (g15658), .I1 (g8177), .I2 (g13264));
AN2X1 gate16338(.O (g15666), .I1 (g5233), .I2 (g13268));
AN2X1 gate16339(.O (g15670), .I1 (g5241), .I2 (g13272));
AN2X1 gate16340(.O (g15671), .I1 (g5242), .I2 (g13273));
AN2X1 gate16341(.O (g15680), .I1 (g5255), .I2 (g13278));
AN2X1 gate16342(.O (g15681), .I1 (g5256), .I2 (g13279));
AN2X1 gate16343(.O (g15699), .I1 (g5278), .I2 (g13283));
AN2X1 gate16344(.O (g15700), .I1 (g5279), .I2 (g13284));
AN2X1 gate16345(.O (g15710), .I1 (g5227), .I2 (g12935));
AN2X1 gate16346(.O (g15717), .I1 (g7924), .I2 (g13285));
AN2X1 gate16347(.O (g15725), .I1 (g5296), .I2 (g13293));
AN2X1 gate16348(.O (g15729), .I1 (g5304), .I2 (g13297));
AN2X1 gate16349(.O (g15730), .I1 (g5305), .I2 (g13298));
AN2X1 gate16350(.O (g15739), .I1 (g5318), .I2 (g13303));
AN2X1 gate16351(.O (g15740), .I1 (g5319), .I2 (g13304));
AN2X1 gate16352(.O (g15753), .I1 (g7542), .I2 (g12962));
AN2X1 gate16353(.O (g15754), .I1 (g7837), .I2 (g13308));
AN2X1 gate16354(.O (g15755), .I1 (g8178), .I2 (g13309));
AN2X1 gate16355(.O (g15765), .I1 (g5333), .I2 (g13324));
AN2X1 gate16356(.O (g15769), .I1 (g5341), .I2 (g13328));
AN2X1 gate16357(.O (g15770), .I1 (g5342), .I2 (g13329));
AN3X1 gate16358(.O (I22028), .I1 (g13004), .I2 (g3018), .I3 (g7549));
AN3X1 gate16359(.O (g15780), .I1 (g7471), .I2 (g3032), .I3 (I22028));
AN2X1 gate16360(.O (g15781), .I1 (g7971), .I2 (g13330));
AN2X1 gate16361(.O (g15793), .I1 (g5361), .I2 (g13347));
AN2X1 gate16362(.O (g15801), .I1 (g7856), .I2 (g13351));
AN2X1 gate16363(.O (g15802), .I1 (g8253), .I2 (g13352));
AN2X1 gate16364(.O (g15817), .I1 (g8025), .I2 (g13373));
AN2X1 gate16365(.O (g15828), .I1 (g7877), .I2 (g13398));
AN2X1 gate16366(.O (g15829), .I1 (g7857), .I2 (g13400));
AN2X1 gate16367(.O (g15840), .I1 (g8098), .I2 (g11620));
AN2X1 gate16368(.O (g15852), .I1 (g7878), .I2 (g11642));
AN3X1 gate16369(.O (I22136), .I1 (g13082), .I2 (g2912), .I3 (g7522));
AN3X1 gate16370(.O (g15902), .I1 (g7607), .I2 (g2920), .I3 (I22136));
AN2X1 gate16371(.O (g15998), .I1 (g5469), .I2 (g11732));
AN2X1 gate16372(.O (g16003), .I1 (g12013), .I2 (g10826));
AN2X1 gate16373(.O (g16004), .I1 (g5587), .I2 (g11734));
AN2X1 gate16374(.O (g16008), .I1 (g5504), .I2 (g11735));
AN2X1 gate16375(.O (g16009), .I1 (g12071), .I2 (g10843));
AN2X1 gate16376(.O (g16010), .I1 (g7639), .I2 (g11736));
AN2X1 gate16377(.O (g16015), .I1 (g12013), .I2 (g10859));
AN2X1 gate16378(.O (g16016), .I1 (g5601), .I2 (g11740));
AN2X1 gate16379(.O (g16017), .I1 (g12130), .I2 (g10862));
AN2X1 gate16380(.O (g16018), .I1 (g6149), .I2 (g11741));
AN2X1 gate16381(.O (g16019), .I1 (g5507), .I2 (g11742));
AN2X1 gate16382(.O (g16028), .I1 (g5543), .I2 (g11745));
AN2X1 gate16383(.O (g16029), .I1 (g12071), .I2 (g10877));
AN2X1 gate16384(.O (g16030), .I1 (g7667), .I2 (g11746));
AN2X1 gate16385(.O (g16031), .I1 (g6227), .I2 (g11747));
AN2X1 gate16386(.O (g16032), .I1 (g12187), .I2 (g10883));
AN2X1 gate16387(.O (g16033), .I1 (g5546), .I2 (g11748));
AN2X1 gate16388(.O (g16045), .I1 (g12013), .I2 (g10892));
AN2X1 gate16389(.O (g16046), .I1 (g5618), .I2 (g11761));
AN2X1 gate16390(.O (g16047), .I1 (g12130), .I2 (g10895));
AN2X1 gate16391(.O (g16048), .I1 (g6170), .I2 (g11762));
AN2X1 gate16392(.O (g16049), .I1 (g6638), .I2 (g11763));
AN2X1 gate16393(.O (g16050), .I1 (g5590), .I2 (g11764));
AN2X1 gate16394(.O (g16051), .I1 (g12235), .I2 (g10901));
AN2X1 gate16395(.O (g16052), .I1 (g5591), .I2 (g11765));
AN2X1 gate16396(.O (g16053), .I1 (g297), .I2 (g11770));
AN2X1 gate16397(.O (g16066), .I1 (g12071), .I2 (g10912));
AN2X1 gate16398(.O (g16067), .I1 (g7700), .I2 (g11774));
AN2X1 gate16399(.O (g16068), .I1 (g6310), .I2 (g11775));
AN2X1 gate16400(.O (g16069), .I1 (g5346), .I2 (g11776));
AN2X1 gate16401(.O (g16070), .I1 (g12187), .I2 (g10921));
AN2X1 gate16402(.O (g16071), .I1 (g5604), .I2 (g11777));
AN2X1 gate16403(.O (g16072), .I1 (g12275), .I2 (g10924));
AN2X1 gate16404(.O (g16073), .I1 (g5605), .I2 (g11778));
AN2X1 gate16405(.O (g16074), .I1 (g5646), .I2 (g11782));
AN2X1 gate16406(.O (g16081), .I1 (g3304), .I2 (g11783));
AN2X1 gate16407(.O (g16089), .I1 (g984), .I2 (g11787));
AN2X1 gate16408(.O (g16100), .I1 (g12130), .I2 (g10937));
AN2X1 gate16409(.O (g16101), .I1 (g6197), .I2 (g11794));
AN2X1 gate16410(.O (g16102), .I1 (g6905), .I2 (g11795));
AN2X1 gate16411(.O (g16103), .I1 (g5621), .I2 (g11796));
AN2X1 gate16412(.O (g16104), .I1 (g12235), .I2 (g10946));
AN2X1 gate16413(.O (g16105), .I1 (g5622), .I2 (g11797));
AN2X1 gate16414(.O (g16106), .I1 (g12308), .I2 (g10949));
AN2X1 gate16415(.O (g16107), .I1 (g5666), .I2 (g11801));
AN2X1 gate16416(.O (g16108), .I1 (g5667), .I2 (g11802));
AN2X1 gate16417(.O (g16109), .I1 (g8277), .I2 (g11803));
AN2X1 gate16418(.O (g16110), .I1 (g516), .I2 (g11804));
AN2X1 gate16419(.O (g16111), .I1 (g5551), .I2 (g13215));
AN2X1 gate16420(.O (g16112), .I1 (g5684), .I2 (g11808));
AN2X1 gate16421(.O (g16119), .I1 (g3460), .I2 (g11809));
AN2X1 gate16422(.O (g16127), .I1 (g1678), .I2 (g11813));
AN2X1 gate16423(.O (g16133), .I1 (g6444), .I2 (g11817));
AN2X1 gate16424(.O (g16134), .I1 (g5363), .I2 (g11818));
AN2X1 gate16425(.O (g16135), .I1 (g12187), .I2 (g10980));
AN2X1 gate16426(.O (g16136), .I1 (g5640), .I2 (g11819));
AN2X1 gate16427(.O (g16137), .I1 (g12275), .I2 (g10983));
AN2X1 gate16428(.O (g16138), .I1 (g5641), .I2 (g11820));
AN2X1 gate16429(.O (g16139), .I1 (g5704), .I2 (g11824));
AN2X1 gate16430(.O (g16140), .I1 (g5705), .I2 (g11825));
AN2X1 gate16431(.O (g16141), .I1 (g5706), .I2 (g11826));
AN2X1 gate16432(.O (g16152), .I1 (g517), .I2 (g11829));
AN2X1 gate16433(.O (g16153), .I1 (g5592), .I2 (g13229));
AN2X1 gate16434(.O (g16158), .I1 (g5718), .I2 (g11834));
AN2X1 gate16435(.O (g16159), .I1 (g5719), .I2 (g11835));
AN2X1 gate16436(.O (g16160), .I1 (g8286), .I2 (g11836));
AN2X1 gate16437(.O (g16161), .I1 (g1202), .I2 (g11837));
AN2X1 gate16438(.O (g16162), .I1 (g5597), .I2 (g13234));
AN2X1 gate16439(.O (g16163), .I1 (g5736), .I2 (g11841));
AN2X1 gate16440(.O (g16170), .I1 (g3616), .I2 (g11842));
AN2X1 gate16441(.O (g16178), .I1 (g2372), .I2 (g11846));
AN2X1 gate16442(.O (g16182), .I1 (g7149), .I2 (g11852));
AN2X1 gate16443(.O (g16183), .I1 (g12235), .I2 (g11014));
AN2X1 gate16444(.O (g16184), .I1 (g5663), .I2 (g11853));
AN2X1 gate16445(.O (g16185), .I1 (g12308), .I2 (g11017));
AN2X1 gate16446(.O (g16186), .I1 (g5753), .I2 (g11856));
AN2X1 gate16447(.O (g16187), .I1 (g5754), .I2 (g11857));
AN2X1 gate16448(.O (g16188), .I1 (g5755), .I2 (g11858));
AN2X1 gate16449(.O (g16197), .I1 (g518), .I2 (g11862));
AN2X1 gate16450(.O (g16198), .I1 (g5762), .I2 (g11866));
AN2X1 gate16451(.O (g16199), .I1 (g5763), .I2 (g11867));
AN2X1 gate16452(.O (g16200), .I1 (g5764), .I2 (g11868));
AN2X1 gate16453(.O (g16211), .I1 (g1203), .I2 (g11871));
AN2X1 gate16454(.O (g16212), .I1 (g5609), .I2 (g13252));
AN2X1 gate16455(.O (g16217), .I1 (g5776), .I2 (g11876));
AN2X1 gate16456(.O (g16218), .I1 (g5777), .I2 (g11877));
AN2X1 gate16457(.O (g16219), .I1 (g8295), .I2 (g11878));
AN2X1 gate16458(.O (g16220), .I1 (g1896), .I2 (g11879));
AN2X1 gate16459(.O (g16221), .I1 (g5614), .I2 (g13257));
AN2X1 gate16460(.O (g16222), .I1 (g5794), .I2 (g11883));
AN2X1 gate16461(.O (g16229), .I1 (g3772), .I2 (g11884));
AN2X1 gate16462(.O (g16237), .I1 (g5379), .I2 (g11886));
AN2X1 gate16463(.O (g16238), .I1 (g12275), .I2 (g11066));
AN2X1 gate16464(.O (g16239), .I1 (g5700), .I2 (g11887));
AN2X1 gate16465(.O (g16240), .I1 (g5804), .I2 (g11891));
AN2X1 gate16466(.O (g16241), .I1 (g5805), .I2 (g11892));
AN2X1 gate16467(.O (g16242), .I1 (g5806), .I2 (g11893));
AN2X1 gate16468(.O (g16250), .I1 (g519), .I2 (g11895));
AN2X1 gate16469(.O (g16251), .I1 (g5812), .I2 (g11898));
AN2X1 gate16470(.O (g16252), .I1 (g5813), .I2 (g11899));
AN2X1 gate16471(.O (g16253), .I1 (g5814), .I2 (g11900));
AN2X1 gate16472(.O (g16262), .I1 (g1204), .I2 (g11904));
AN2X1 gate16473(.O (g16263), .I1 (g5821), .I2 (g11908));
AN2X1 gate16474(.O (g16264), .I1 (g5822), .I2 (g11909));
AN2X1 gate16475(.O (g16265), .I1 (g5823), .I2 (g11910));
AN2X1 gate16476(.O (g16276), .I1 (g1897), .I2 (g11913));
AN2X1 gate16477(.O (g16277), .I1 (g5634), .I2 (g13275));
AN2X1 gate16478(.O (g16282), .I1 (g5835), .I2 (g11918));
AN2X1 gate16479(.O (g16283), .I1 (g5836), .I2 (g11919));
AN2X1 gate16480(.O (g16284), .I1 (g8304), .I2 (g11920));
AN2X1 gate16481(.O (g16285), .I1 (g2590), .I2 (g11921));
AN2X1 gate16482(.O (g16286), .I1 (g5639), .I2 (g13280));
AN2X1 gate16483(.O (g16288), .I1 (g12308), .I2 (g11129));
AN2X1 gate16484(.O (g16289), .I1 (g5853), .I2 (g11929));
AN2X1 gate16485(.O (g16290), .I1 (g5854), .I2 (g11930));
AN2X1 gate16486(.O (g16291), .I1 (g5855), .I2 (g11931));
AN2X1 gate16487(.O (g16292), .I1 (g294), .I2 (g11932));
AN2X1 gate16488(.O (g16298), .I1 (g520), .I2 (g11936));
AN2X1 gate16489(.O (g16299), .I1 (g5860), .I2 (g11941));
AN2X1 gate16490(.O (g16300), .I1 (g5861), .I2 (g11942));
AN2X1 gate16491(.O (g16301), .I1 (g5862), .I2 (g11943));
AN2X1 gate16492(.O (g16309), .I1 (g1205), .I2 (g11945));
AN2X1 gate16493(.O (g16310), .I1 (g5868), .I2 (g11948));
AN2X1 gate16494(.O (g16311), .I1 (g5869), .I2 (g11949));
AN2X1 gate16495(.O (g16312), .I1 (g5870), .I2 (g11950));
AN2X1 gate16496(.O (g16321), .I1 (g1898), .I2 (g11954));
AN2X1 gate16497(.O (g16322), .I1 (g5877), .I2 (g11958));
AN2X1 gate16498(.O (g16323), .I1 (g5878), .I2 (g11959));
AN2X1 gate16499(.O (g16324), .I1 (g5879), .I2 (g11960));
AN2X1 gate16500(.O (g16335), .I1 (g2591), .I2 (g11963));
AN2X1 gate16501(.O (g16336), .I1 (g5662), .I2 (g13300));
AN2X1 gate16502(.O (g16342), .I1 (g5894), .I2 (g11968));
AN2X1 gate16503(.O (g16343), .I1 (g5895), .I2 (g11969));
AN2X1 gate16504(.O (g16344), .I1 (g5896), .I2 (g11970));
AN2X1 gate16505(.O (g16345), .I1 (g5897), .I2 (g11971));
AN2X1 gate16506(.O (g16346), .I1 (g295), .I2 (g11972));
AN2X1 gate16507(.O (g16347), .I1 (g5900), .I2 (g11982));
AN2X1 gate16508(.O (g16348), .I1 (g5901), .I2 (g11983));
AN2X1 gate16509(.O (g16349), .I1 (g5902), .I2 (g11984));
AN2X1 gate16510(.O (g16350), .I1 (g981), .I2 (g11985));
AN2X1 gate16511(.O (g16356), .I1 (g1206), .I2 (g11989));
AN2X1 gate16512(.O (g16357), .I1 (g5907), .I2 (g11994));
AN2X1 gate16513(.O (g16358), .I1 (g5908), .I2 (g11995));
AN2X1 gate16514(.O (g16359), .I1 (g5909), .I2 (g11996));
AN2X1 gate16515(.O (g16367), .I1 (g1899), .I2 (g11998));
AN2X1 gate16516(.O (g16368), .I1 (g5915), .I2 (g12001));
AN2X1 gate16517(.O (g16369), .I1 (g5916), .I2 (g12002));
AN2X1 gate16518(.O (g16370), .I1 (g5917), .I2 (g12003));
AN2X1 gate16519(.O (g16379), .I1 (g2592), .I2 (g12007));
AN2X1 gate16520(.O (g16380), .I1 (g5925), .I2 (g12020));
AN2X1 gate16521(.O (g16381), .I1 (g5926), .I2 (g12021));
AN2X1 gate16522(.O (g16382), .I1 (g5927), .I2 (g12022));
AN2X1 gate16523(.O (g16383), .I1 (g5928), .I2 (g12023));
AN2X1 gate16524(.O (g16384), .I1 (g296), .I2 (g12024));
AN2X1 gate16525(.O (g16385), .I1 (g5714), .I2 (g13336));
AN2X1 gate16526(.O (g16386), .I1 (g5933), .I2 (g12037));
AN2X1 gate16527(.O (g16387), .I1 (g5934), .I2 (g12038));
AN2X1 gate16528(.O (g16388), .I1 (g5935), .I2 (g12039));
AN2X1 gate16529(.O (g16389), .I1 (g5936), .I2 (g12040));
AN2X1 gate16530(.O (g16390), .I1 (g982), .I2 (g12041));
AN2X1 gate16531(.O (g16391), .I1 (g5939), .I2 (g12051));
AN2X1 gate16532(.O (g16392), .I1 (g5940), .I2 (g12052));
AN2X1 gate16533(.O (g16393), .I1 (g5941), .I2 (g12053));
AN2X1 gate16534(.O (g16394), .I1 (g1675), .I2 (g12054));
AN2X1 gate16535(.O (g16400), .I1 (g1900), .I2 (g12058));
AN2X1 gate16536(.O (g16401), .I1 (g5946), .I2 (g12063));
AN2X1 gate16537(.O (g16402), .I1 (g5947), .I2 (g12064));
AN2X1 gate16538(.O (g16403), .I1 (g5948), .I2 (g12065));
AN2X1 gate16539(.O (g16411), .I1 (g2593), .I2 (g12067));
AN2X1 gate16540(.O (g16413), .I1 (g5954), .I2 (g12075));
AN2X1 gate16541(.O (g16414), .I1 (g5955), .I2 (g12076));
AN2X1 gate16542(.O (g16415), .I1 (g5956), .I2 (g12077));
AN2X1 gate16543(.O (g16416), .I1 (g5957), .I2 (g12078));
AN2X1 gate16544(.O (g16417), .I1 (g5759), .I2 (g13356));
AN2X1 gate16545(.O (g16418), .I1 (g5959), .I2 (g12084));
AN2X1 gate16546(.O (g16419), .I1 (g5960), .I2 (g12085));
AN2X1 gate16547(.O (g16420), .I1 (g5961), .I2 (g12086));
AN2X1 gate16548(.O (g16421), .I1 (g5962), .I2 (g12087));
AN2X1 gate16549(.O (g16422), .I1 (g983), .I2 (g12088));
AN2X1 gate16550(.O (g16423), .I1 (g5772), .I2 (g13361));
AN2X1 gate16551(.O (g16424), .I1 (g5967), .I2 (g12101));
AN2X1 gate16552(.O (g16425), .I1 (g5968), .I2 (g12102));
AN2X1 gate16553(.O (g16426), .I1 (g5969), .I2 (g12103));
AN2X1 gate16554(.O (g16427), .I1 (g5970), .I2 (g12104));
AN2X1 gate16555(.O (g16428), .I1 (g1676), .I2 (g12105));
AN2X1 gate16556(.O (g16429), .I1 (g5973), .I2 (g12115));
AN2X1 gate16557(.O (g16430), .I1 (g5974), .I2 (g12116));
AN2X1 gate16558(.O (g16431), .I1 (g5975), .I2 (g12117));
AN2X1 gate16559(.O (g16432), .I1 (g2369), .I2 (g12118));
AN2X1 gate16560(.O (g16438), .I1 (g2594), .I2 (g12122));
AN2X1 gate16561(.O (g16443), .I1 (g5980), .I2 (g12134));
AN2X1 gate16562(.O (g16444), .I1 (g5981), .I2 (g12135));
AN2X1 gate16563(.O (g16445), .I1 (g5808), .I2 (g13381));
AN2X1 gate16564(.O (g16447), .I1 (g5983), .I2 (g12147));
AN2X1 gate16565(.O (g16448), .I1 (g5984), .I2 (g12148));
AN2X1 gate16566(.O (g16449), .I1 (g5985), .I2 (g12149));
AN2X1 gate16567(.O (g16450), .I1 (g5986), .I2 (g12150));
AN2X1 gate16568(.O (g16451), .I1 (g5818), .I2 (g13386));
AN2X1 gate16569(.O (g16452), .I1 (g5988), .I2 (g12156));
AN2X1 gate16570(.O (g16453), .I1 (g5989), .I2 (g12157));
AN2X1 gate16571(.O (g16454), .I1 (g5990), .I2 (g12158));
AN2X1 gate16572(.O (g16455), .I1 (g5991), .I2 (g12159));
AN2X1 gate16573(.O (g16456), .I1 (g1677), .I2 (g12160));
AN2X1 gate16574(.O (g16457), .I1 (g5831), .I2 (g13391));
AN2X1 gate16575(.O (g16458), .I1 (g5996), .I2 (g12173));
AN2X1 gate16576(.O (g16459), .I1 (g5997), .I2 (g12174));
AN2X1 gate16577(.O (g16460), .I1 (g5998), .I2 (g12175));
AN2X1 gate16578(.O (g16461), .I1 (g5999), .I2 (g12176));
AN2X1 gate16579(.O (g16462), .I1 (g2370), .I2 (g12177));
AN4X1 gate16580(.O (g16505), .I1 (g14776), .I2 (g14797), .I3 (g16142), .I4 (g16243));
AN4X1 gate16581(.O (g16513), .I1 (g15065), .I2 (g13724), .I3 (g13764), .I4 (g13797));
AN4X1 gate16582(.O (g16527), .I1 (g14811), .I2 (g14849), .I3 (g16201), .I4 (g16302));
AN4X1 gate16583(.O (g16535), .I1 (g15161), .I2 (g13774), .I3 (g13805), .I4 (g13825));
AN4X1 gate16584(.O (g16558), .I1 (g14863), .I2 (g14922), .I3 (g16266), .I4 (g16360));
AN4X1 gate16585(.O (g16590), .I1 (g14936), .I2 (g15003), .I3 (g16325), .I4 (g16404));
AN2X1 gate16586(.O (g16607), .I1 (g15022), .I2 (g15096));
AN2X1 gate16587(.O (g16625), .I1 (g15118), .I2 (g15188));
AN2X1 gate16588(.O (g16639), .I1 (g15210), .I2 (g15274));
AN2X1 gate16589(.O (g16650), .I1 (g15296), .I2 (g15366));
AN2X1 gate16590(.O (g16850), .I1 (g6226), .I2 (g14764));
AN2X1 gate16591(.O (g16855), .I1 (g15722), .I2 (g8646));
AN2X1 gate16592(.O (g16856), .I1 (g6443), .I2 (g14794));
AN2X1 gate16593(.O (g16859), .I1 (g15762), .I2 (g8662));
AN2X1 gate16594(.O (g16864), .I1 (g15790), .I2 (g8681));
AN2X1 gate16595(.O (g16865), .I1 (g6896), .I2 (g14881));
AN2X1 gate16596(.O (g16879), .I1 (g15813), .I2 (g8693));
AN2X1 gate16597(.O (g16894), .I1 (g7156), .I2 (g14959));
AN2X1 gate16598(.O (g16907), .I1 (g7335), .I2 (g15017));
AN2X1 gate16599(.O (g16908), .I1 (g7838), .I2 (g15032));
AN2X1 gate16600(.O (g16909), .I1 (g6908), .I2 (g15033));
AN2X1 gate16601(.O (g16923), .I1 (g7352), .I2 (g15048));
AN2X1 gate16602(.O (g16938), .I1 (g7858), .I2 (g15128));
AN2X1 gate16603(.O (g16939), .I1 (g7158), .I2 (g15129));
AN2X1 gate16604(.O (g16953), .I1 (g7482), .I2 (g15144));
AN2X1 gate16605(.O (g16964), .I1 (g7520), .I2 (g15170));
AN2X1 gate16606(.O (g16966), .I1 (g7529), .I2 (g15174));
AN2X1 gate16607(.O (g16967), .I1 (g7827), .I2 (g15175));
AN2X1 gate16608(.O (g16968), .I1 (g6672), .I2 (g15176));
AN2X1 gate16609(.O (g16969), .I1 (g7888), .I2 (g15220));
AN2X1 gate16610(.O (g16970), .I1 (g7354), .I2 (g15221));
AN2X1 gate16611(.O (g16984), .I1 (g7538), .I2 (g15236));
AN2X1 gate16612(.O (g16987), .I1 (g7555), .I2 (g15260));
AN2X1 gate16613(.O (g16988), .I1 (g7842), .I2 (g15261));
AN2X1 gate16614(.O (g16989), .I1 (g6974), .I2 (g15262));
AN2X1 gate16615(.O (g16990), .I1 (g7912), .I2 (g15306));
AN2X1 gate16616(.O (g16991), .I1 (g7484), .I2 (g15307));
AN2X1 gate16617(.O (g16993), .I1 (g7576), .I2 (g15322));
AN2X1 gate16618(.O (g16994), .I1 (g7819), .I2 (g15323));
AN2X1 gate16619(.O (g16997), .I1 (g7578), .I2 (g15352));
AN2X1 gate16620(.O (g16998), .I1 (g7862), .I2 (g15353));
AN2X1 gate16621(.O (g16999), .I1 (g7224), .I2 (g15354));
AN3X1 gate16622(.O (g17001), .I1 (g3254), .I2 (g10694), .I3 (g14144));
AN2X1 gate16623(.O (g17015), .I1 (g7996), .I2 (g15390));
AN2X1 gate16624(.O (g17017), .I1 (g7590), .I2 (g15408));
AN2X1 gate16625(.O (g17018), .I1 (g7830), .I2 (g15409));
AN2X1 gate16626(.O (g17021), .I1 (g7592), .I2 (g15438));
AN2X1 gate16627(.O (g17022), .I1 (g7892), .I2 (g15439));
AN2X1 gate16628(.O (g17023), .I1 (g7420), .I2 (g15440));
AN2X1 gate16629(.O (g17028), .I1 (g7604), .I2 (g15458));
AN3X1 gate16630(.O (g17031), .I1 (g3410), .I2 (g10714), .I3 (g14259));
AN2X1 gate16631(.O (g17045), .I1 (g8071), .I2 (g15474));
AN2X1 gate16632(.O (g17047), .I1 (g7605), .I2 (g15492));
AN2X1 gate16633(.O (g17048), .I1 (g7845), .I2 (g15493));
AN2X1 gate16634(.O (g17055), .I1 (g7153), .I2 (g15524));
AN2X1 gate16635(.O (g17056), .I1 (g7953), .I2 (g15525));
AN2X1 gate16636(.O (g17062), .I1 (g7613), .I2 (g15544));
AN3X1 gate16637(.O (g17065), .I1 (g3566), .I2 (g10735), .I3 (g14381));
AN2X1 gate16638(.O (g17079), .I1 (g8156), .I2 (g15560));
AN2X1 gate16639(.O (g17081), .I1 (g7614), .I2 (g15578));
AN2X1 gate16640(.O (g17082), .I1 (g7865), .I2 (g15579));
AN2X1 gate16641(.O (g17084), .I1 (g7629), .I2 (g13954));
AN2X1 gate16642(.O (g17090), .I1 (g7349), .I2 (g15602));
AN2X1 gate16643(.O (g17091), .I1 (g8004), .I2 (g15603));
AN2X1 gate16644(.O (g17097), .I1 (g7622), .I2 (g15622));
AN3X1 gate16645(.O (g17100), .I1 (g3722), .I2 (g10754), .I3 (g14493));
AN2X1 gate16646(.O (g17114), .I1 (g8242), .I2 (g15638));
AN2X1 gate16647(.O (g17116), .I1 (g7649), .I2 (g14008));
AN2X1 gate16648(.O (g17117), .I1 (g7906), .I2 (g15665));
AN2X1 gate16649(.O (g17122), .I1 (g7658), .I2 (g14024));
AN2X1 gate16650(.O (g17128), .I1 (g7479), .I2 (g15678));
AN2X1 gate16651(.O (g17129), .I1 (g8079), .I2 (g15679));
AN2X1 gate16652(.O (g17135), .I1 (g7638), .I2 (g15698));
AN2X1 gate16653(.O (g17138), .I1 (g7676), .I2 (g14068));
AN2X1 gate16654(.O (g17143), .I1 (g7685), .I2 (g14099));
AN2X1 gate16655(.O (g17144), .I1 (g7958), .I2 (g15724));
AN2X1 gate16656(.O (g17149), .I1 (g7694), .I2 (g14115));
AN2X1 gate16657(.O (g17155), .I1 (g7535), .I2 (g15737));
AN2X1 gate16658(.O (g17156), .I1 (g8164), .I2 (g15738));
AN2X1 gate16659(.O (g17161), .I1 (g7712), .I2 (g14183));
AN2X1 gate16660(.O (g17166), .I1 (g7721), .I2 (g14214));
AN2X1 gate16661(.O (g17167), .I1 (g8009), .I2 (g15764));
AN2X1 gate16662(.O (g17172), .I1 (g7730), .I2 (g14230));
AN2X1 gate16663(.O (g17176), .I1 (g7742), .I2 (g14298));
AN2X1 gate16664(.O (g17181), .I1 (g7751), .I2 (g14329));
AN2X1 gate16665(.O (g17182), .I1 (g8084), .I2 (g15792));
AN2X1 gate16666(.O (g17193), .I1 (g7766), .I2 (g14420));
AN2X1 gate16667(.O (g17268), .I1 (g8024), .I2 (g15991));
AN2X1 gate16668(.O (g17301), .I1 (g8097), .I2 (g15994));
AN2X1 gate16669(.O (g17339), .I1 (g8176), .I2 (g15997));
AN2X1 gate16670(.O (g17352), .I1 (g3942), .I2 (g14960));
AN2X1 gate16671(.O (g17353), .I1 (g3945), .I2 (g14963));
AN2X1 gate16672(.O (g17381), .I1 (g8250), .I2 (g16001));
AN2X1 gate16673(.O (g17382), .I1 (g8252), .I2 (g16002));
AN2X1 gate16674(.O (g17393), .I1 (g3941), .I2 (g16005));
AN2X1 gate16675(.O (g17395), .I1 (g6177), .I2 (g15034));
AN2X1 gate16676(.O (g17396), .I1 (g4020), .I2 (g15037));
AN2X1 gate16677(.O (g17397), .I1 (g4023), .I2 (g15040));
AN2X1 gate16678(.O (g17398), .I1 (g4026), .I2 (g15043));
AN2X1 gate16679(.O (g17408), .I1 (g4049), .I2 (g15049));
AN2X1 gate16680(.O (g17409), .I1 (g4052), .I2 (g15052));
AN2X1 gate16681(.O (g17428), .I1 (g3994), .I2 (g16007));
AN2X1 gate16682(.O (g17446), .I1 (g6284), .I2 (g16011));
AN2X1 gate16683(.O (g17447), .I1 (g4115), .I2 (g15106));
AN2X1 gate16684(.O (g17448), .I1 (g4118), .I2 (g15109));
AN2X1 gate16685(.O (g17449), .I1 (g4121), .I2 (g15112));
AN2X1 gate16686(.O (g17450), .I1 (g4124), .I2 (g15115));
AN2X1 gate16687(.O (g17460), .I1 (g4048), .I2 (g16012));
AN2X1 gate16688(.O (g17461), .I1 (g6209), .I2 (g15130));
AN2X1 gate16689(.O (g17462), .I1 (g4147), .I2 (g15133));
AN2X1 gate16690(.O (g17463), .I1 (g4150), .I2 (g15136));
AN2X1 gate16691(.O (g17464), .I1 (g4153), .I2 (g15139));
AN2X1 gate16692(.O (g17474), .I1 (g4176), .I2 (g15145));
AN2X1 gate16693(.O (g17475), .I1 (g4179), .I2 (g15148));
AN2X1 gate16694(.O (g17485), .I1 (g4089), .I2 (g16013));
AN2X1 gate16695(.O (g17486), .I1 (g4091), .I2 (g16014));
AN2X1 gate16696(.O (g17506), .I1 (g6675), .I2 (g16023));
AN2X1 gate16697(.O (g17508), .I1 (g4225), .I2 (g15179));
AN2X1 gate16698(.O (g17509), .I1 (g4228), .I2 (g15182));
AN2X1 gate16699(.O (g17510), .I1 (g4231), .I2 (g15185));
AN2X1 gate16700(.O (g17526), .I1 (g6421), .I2 (g16025));
AN2X1 gate16701(.O (g17527), .I1 (g4254), .I2 (g15198));
AN2X1 gate16702(.O (g17528), .I1 (g4257), .I2 (g15201));
AN2X1 gate16703(.O (g17529), .I1 (g4260), .I2 (g15204));
AN2X1 gate16704(.O (g17530), .I1 (g4263), .I2 (g15207));
AN2X1 gate16705(.O (g17540), .I1 (g4175), .I2 (g16026));
AN2X1 gate16706(.O (g17541), .I1 (g6298), .I2 (g15222));
AN2X1 gate16707(.O (g17542), .I1 (g4286), .I2 (g15225));
AN2X1 gate16708(.O (g17543), .I1 (g4289), .I2 (g15228));
AN2X1 gate16709(.O (g17544), .I1 (g4292), .I2 (g15231));
AN2X1 gate16710(.O (g17554), .I1 (g4315), .I2 (g15237));
AN2X1 gate16711(.O (g17555), .I1 (g4318), .I2 (g15240));
AN2X1 gate16712(.O (g17556), .I1 (g4201), .I2 (g16027));
AN2X1 gate16713(.O (g17576), .I1 (g4348), .I2 (g15248));
AN2X1 gate16714(.O (g17577), .I1 (g4351), .I2 (g15251));
AN2X1 gate16715(.O (g17578), .I1 (g4354), .I2 (g15254));
AN2X1 gate16716(.O (g17597), .I1 (g6977), .I2 (g16039));
AN2X1 gate16717(.O (g17598), .I1 (g4380), .I2 (g15265));
AN2X1 gate16718(.O (g17599), .I1 (g4383), .I2 (g15268));
AN2X1 gate16719(.O (g17600), .I1 (g4386), .I2 (g15271));
AN2X1 gate16720(.O (g17616), .I1 (g6626), .I2 (g16041));
AN2X1 gate16721(.O (g17617), .I1 (g4409), .I2 (g15284));
AN2X1 gate16722(.O (g17618), .I1 (g4412), .I2 (g15287));
AN2X1 gate16723(.O (g17619), .I1 (g4415), .I2 (g15290));
AN2X1 gate16724(.O (g17620), .I1 (g4418), .I2 (g15293));
AN2X1 gate16725(.O (g17630), .I1 (g4314), .I2 (g16042));
AN2X1 gate16726(.O (g17631), .I1 (g6435), .I2 (g15308));
AN2X1 gate16727(.O (g17632), .I1 (g4441), .I2 (g15311));
AN2X1 gate16728(.O (g17633), .I1 (g4444), .I2 (g15314));
AN2X1 gate16729(.O (g17634), .I1 (g4447), .I2 (g15317));
AN2X1 gate16730(.O (g17635), .I1 (g4322), .I2 (g16043));
AN2X1 gate16731(.O (g17636), .I1 (g4324), .I2 (g16044));
AN2X1 gate16732(.O (g17652), .I1 (g4480), .I2 (g15326));
AN2X1 gate16733(.O (g17653), .I1 (g4483), .I2 (g15329));
AN2X1 gate16734(.O (g17654), .I1 (g4486), .I2 (g15332));
AN2X1 gate16735(.O (g17673), .I1 (g4517), .I2 (g15340));
AN2X1 gate16736(.O (g17674), .I1 (g4520), .I2 (g15343));
AN2X1 gate16737(.O (g17675), .I1 (g4523), .I2 (g15346));
AN2X1 gate16738(.O (g17694), .I1 (g7227), .I2 (g16061));
AN2X1 gate16739(.O (g17695), .I1 (g4549), .I2 (g15357));
AN2X1 gate16740(.O (g17696), .I1 (g4552), .I2 (g15360));
AN2X1 gate16741(.O (g17697), .I1 (g4555), .I2 (g15363));
AN2X1 gate16742(.O (g17713), .I1 (g6890), .I2 (g16063));
AN2X1 gate16743(.O (g17714), .I1 (g4578), .I2 (g15376));
AN2X1 gate16744(.O (g17715), .I1 (g4581), .I2 (g15379));
AN2X1 gate16745(.O (g17716), .I1 (g4584), .I2 (g15382));
AN2X1 gate16746(.O (g17717), .I1 (g4587), .I2 (g15385));
AN2X1 gate16747(.O (g17718), .I1 (g4451), .I2 (g16064));
AN2X1 gate16748(.O (g17719), .I1 (g2993), .I2 (g16065));
AN2X1 gate16749(.O (g17734), .I1 (g4611), .I2 (g15393));
AN2X1 gate16750(.O (g17735), .I1 (g4614), .I2 (g15396));
AN2X1 gate16751(.O (g17736), .I1 (g4617), .I2 (g15399));
AN2X1 gate16752(.O (g17737), .I1 (g4626), .I2 (g15404));
AN2X1 gate16753(.O (g17752), .I1 (g4656), .I2 (g15412));
AN2X1 gate16754(.O (g17753), .I1 (g4659), .I2 (g15415));
AN2X1 gate16755(.O (g17754), .I1 (g4662), .I2 (g15418));
AN2X1 gate16756(.O (g17773), .I1 (g4693), .I2 (g15426));
AN2X1 gate16757(.O (g17774), .I1 (g4696), .I2 (g15429));
AN2X1 gate16758(.O (g17775), .I1 (g4699), .I2 (g15432));
AN2X1 gate16759(.O (g17794), .I1 (g7423), .I2 (g16097));
AN2X1 gate16760(.O (g17795), .I1 (g4725), .I2 (g15443));
AN2X1 gate16761(.O (g17796), .I1 (g4728), .I2 (g15446));
AN2X1 gate16762(.O (g17797), .I1 (g4731), .I2 (g15449));
AN2X1 gate16763(.O (g17798), .I1 (g4591), .I2 (g16099));
AN2X1 gate16764(.O (g17812), .I1 (g4754), .I2 (g15461));
AN2X1 gate16765(.O (g17813), .I1 (g4757), .I2 (g15464));
AN2X1 gate16766(.O (g17814), .I1 (g4760), .I2 (g15467));
AN2X1 gate16767(.O (g17824), .I1 (g4766), .I2 (g15471));
AN2X1 gate16768(.O (g17835), .I1 (g4788), .I2 (g15477));
AN2X1 gate16769(.O (g17836), .I1 (g4791), .I2 (g15480));
AN2X1 gate16770(.O (g17837), .I1 (g4794), .I2 (g15483));
AN2X1 gate16771(.O (g17838), .I1 (g4803), .I2 (g15488));
AN2X1 gate16772(.O (g17853), .I1 (g4833), .I2 (g15496));
AN2X1 gate16773(.O (g17854), .I1 (g4836), .I2 (g15499));
AN2X1 gate16774(.O (g17855), .I1 (g4839), .I2 (g15502));
AN2X1 gate16775(.O (g17874), .I1 (g4870), .I2 (g15510));
AN2X1 gate16776(.O (g17875), .I1 (g4873), .I2 (g15513));
AN2X1 gate16777(.O (g17876), .I1 (g4876), .I2 (g15516));
AN2X1 gate16778(.O (g17877), .I1 (g2998), .I2 (g15521));
AN2X1 gate16779(.O (g17900), .I1 (g4899), .I2 (g15528));
AN2X1 gate16780(.O (g17901), .I1 (g4902), .I2 (g15531));
AN2X1 gate16781(.O (g17902), .I1 (g4905), .I2 (g15534));
AN2X1 gate16782(.O (g17912), .I1 (g4908), .I2 (g15537));
AN2X1 gate16783(.O (g17924), .I1 (g4930), .I2 (g15547));
AN2X1 gate16784(.O (g17925), .I1 (g4933), .I2 (g15550));
AN2X1 gate16785(.O (g17926), .I1 (g4936), .I2 (g15553));
AN2X1 gate16786(.O (g17936), .I1 (g4942), .I2 (g15557));
AN2X1 gate16787(.O (g17947), .I1 (g4964), .I2 (g15563));
AN2X1 gate16788(.O (g17948), .I1 (g4967), .I2 (g15566));
AN2X1 gate16789(.O (g17949), .I1 (g4970), .I2 (g15569));
AN2X1 gate16790(.O (g17950), .I1 (g4979), .I2 (g15574));
AN2X1 gate16791(.O (g17965), .I1 (g5009), .I2 (g15582));
AN2X1 gate16792(.O (g17966), .I1 (g5012), .I2 (g15585));
AN2X1 gate16793(.O (g17967), .I1 (g5015), .I2 (g15588));
AN2X1 gate16794(.O (g17989), .I1 (g5035), .I2 (g15596));
AN2X1 gate16795(.O (g17990), .I1 (g5038), .I2 (g15599));
AN2X1 gate16796(.O (g18011), .I1 (g5058), .I2 (g15606));
AN2X1 gate16797(.O (g18012), .I1 (g5061), .I2 (g15609));
AN2X1 gate16798(.O (g18013), .I1 (g5064), .I2 (g15612));
AN2X1 gate16799(.O (g18023), .I1 (g5067), .I2 (g15615));
AN2X1 gate16800(.O (g18035), .I1 (g5089), .I2 (g15625));
AN2X1 gate16801(.O (g18036), .I1 (g5092), .I2 (g15628));
AN2X1 gate16802(.O (g18037), .I1 (g5095), .I2 (g15631));
AN2X1 gate16803(.O (g18047), .I1 (g5101), .I2 (g15635));
AN2X1 gate16804(.O (g18058), .I1 (g5123), .I2 (g15641));
AN2X1 gate16805(.O (g18059), .I1 (g5126), .I2 (g15644));
AN2X1 gate16806(.O (g18060), .I1 (g5129), .I2 (g15647));
AN2X1 gate16807(.O (g18061), .I1 (g5138), .I2 (g15652));
AN2X1 gate16808(.O (g18062), .I1 (g7462), .I2 (g15655));
AN2X1 gate16809(.O (g18088), .I1 (g5150), .I2 (g15667));
AN2X1 gate16810(.O (g18106), .I1 (g5164), .I2 (g15672));
AN2X1 gate16811(.O (g18107), .I1 (g5167), .I2 (g15675));
AN2X1 gate16812(.O (g18128), .I1 (g5187), .I2 (g15682));
AN2X1 gate16813(.O (g18129), .I1 (g5190), .I2 (g15685));
AN2X1 gate16814(.O (g18130), .I1 (g5193), .I2 (g15688));
AN2X1 gate16815(.O (g18140), .I1 (g5196), .I2 (g15691));
AN2X1 gate16816(.O (g18152), .I1 (g5218), .I2 (g15701));
AN2X1 gate16817(.O (g18153), .I1 (g5221), .I2 (g15704));
AN2X1 gate16818(.O (g18154), .I1 (g5224), .I2 (g15707));
AN2X1 gate16819(.O (g18164), .I1 (g5230), .I2 (g15711));
AN2X1 gate16820(.O (g18165), .I1 (g2883), .I2 (g16287));
AN2X1 gate16821(.O (g18169), .I1 (g7527), .I2 (g15714));
AN2X1 gate16822(.O (g18204), .I1 (g5243), .I2 (g15726));
AN2X1 gate16823(.O (g18222), .I1 (g5257), .I2 (g15731));
AN2X1 gate16824(.O (g18223), .I1 (g5260), .I2 (g15734));
AN2X1 gate16825(.O (g18244), .I1 (g5280), .I2 (g15741));
AN2X1 gate16826(.O (g18245), .I1 (g5283), .I2 (g15744));
AN2X1 gate16827(.O (g18246), .I1 (g5286), .I2 (g15747));
AN2X1 gate16828(.O (g18256), .I1 (g5289), .I2 (g15750));
AN2X1 gate16829(.O (g18311), .I1 (g5306), .I2 (g15766));
AN2X1 gate16830(.O (g18329), .I1 (g5320), .I2 (g15771));
AN2X1 gate16831(.O (g18330), .I1 (g5323), .I2 (g15774));
AN2X1 gate16832(.O (g18333), .I1 (g2888), .I2 (g15777));
AN2X1 gate16833(.O (g18404), .I1 (g5343), .I2 (g15794));
AN3X1 gate16834(.O (I24619), .I1 (g14776), .I2 (g14837), .I3 (g16142));
AN3X1 gate16835(.O (g18547), .I1 (g13677), .I2 (g13750), .I3 (I24619));
AN3X1 gate16836(.O (I24689), .I1 (g14811), .I2 (g14910), .I3 (g16201));
AN3X1 gate16837(.O (g18597), .I1 (g13714), .I2 (g13791), .I3 (I24689));
AN3X1 gate16838(.O (I24738), .I1 (g14863), .I2 (g14991), .I3 (g16266));
AN3X1 gate16839(.O (g18629), .I1 (g13764), .I2 (g13819), .I3 (I24738));
AN3X1 gate16840(.O (I24758), .I1 (g14936), .I2 (g15080), .I3 (g16325));
AN3X1 gate16841(.O (g18638), .I1 (g13805), .I2 (g13840), .I3 (I24758));
AN4X1 gate16842(.O (g18645), .I1 (g14776), .I2 (g14895), .I3 (g16142), .I4 (g13750));
AN3X1 gate16843(.O (g18647), .I1 (g14895), .I2 (g16142), .I3 (g16243));
AN4X1 gate16844(.O (g18648), .I1 (g14811), .I2 (g14976), .I3 (g16201), .I4 (g13791));
AN4X1 gate16845(.O (g18649), .I1 (g14776), .I2 (g14837), .I3 (g13657), .I4 (g16189));
AN3X1 gate16846(.O (g18650), .I1 (g14976), .I2 (g16201), .I3 (g16302));
AN4X1 gate16847(.O (g18651), .I1 (g14863), .I2 (g15065), .I3 (g16266), .I4 (g13819));
AN4X1 gate16848(.O (g18652), .I1 (g14797), .I2 (g13657), .I3 (g13677), .I4 (g16243));
AN4X1 gate16849(.O (g18653), .I1 (g14811), .I2 (g14910), .I3 (g13687), .I4 (g16254));
AN3X1 gate16850(.O (g18654), .I1 (g15065), .I2 (g16266), .I3 (g16360));
AN4X1 gate16851(.O (g18655), .I1 (g14936), .I2 (g15161), .I3 (g16325), .I4 (g13840));
AN4X1 gate16852(.O (g18665), .I1 (g14776), .I2 (g14837), .I3 (g16189), .I4 (g13706));
AN4X1 gate16853(.O (g18666), .I1 (g14849), .I2 (g13687), .I3 (g13714), .I4 (g16302));
AN4X1 gate16854(.O (g18667), .I1 (g14863), .I2 (g14991), .I3 (g13724), .I4 (g16313));
AN3X1 gate16855(.O (g18668), .I1 (g15161), .I2 (g16325), .I3 (g16404));
AN4X1 gate16856(.O (g18688), .I1 (g14811), .I2 (g14910), .I3 (g16254), .I4 (g13756));
AN4X1 gate16857(.O (g18689), .I1 (g14922), .I2 (g13724), .I3 (g13764), .I4 (g16360));
AN4X1 gate16858(.O (g18690), .I1 (g14936), .I2 (g15080), .I3 (g13774), .I4 (g16371));
AN4X1 gate16859(.O (g18717), .I1 (g14863), .I2 (g14991), .I3 (g16313), .I4 (g13797));
AN4X1 gate16860(.O (g18718), .I1 (g15003), .I2 (g13774), .I3 (g13805), .I4 (g16404));
AN4X1 gate16861(.O (g18753), .I1 (g14936), .I2 (g15080), .I3 (g16371), .I4 (g13825));
AN2X1 gate16862(.O (g18982), .I1 (g13519), .I2 (g16154));
AN2X1 gate16863(.O (g18990), .I1 (g13530), .I2 (g16213));
AN4X1 gate16864(.O (g18994), .I1 (g14895), .I2 (g13657), .I3 (g13677), .I4 (g13706));
AN2X1 gate16865(.O (g18997), .I1 (g13541), .I2 (g16278));
AN4X1 gate16866(.O (g19007), .I1 (g14976), .I2 (g13687), .I3 (g13714), .I4 (g13756));
AN2X1 gate16867(.O (g19010), .I1 (g13552), .I2 (g16337));
AN4X1 gate16868(.O (g19063), .I1 (g18679), .I2 (g14910), .I3 (g13687), .I4 (g16254));
AN4X1 gate16869(.O (g19079), .I1 (g14797), .I2 (g18692), .I3 (g16142), .I4 (g16189));
AN4X1 gate16870(.O (g19080), .I1 (g18708), .I2 (g14991), .I3 (g13724), .I4 (g16313));
AN2X1 gate16871(.O (g19087), .I1 (g17215), .I2 (g16540));
AN4X1 gate16872(.O (g19088), .I1 (g18656), .I2 (g14797), .I3 (g16189), .I4 (g13706));
AN4X1 gate16873(.O (g19089), .I1 (g14849), .I2 (g18728), .I3 (g16201), .I4 (g16254));
AN4X1 gate16874(.O (g19090), .I1 (g18744), .I2 (g15080), .I3 (g13774), .I4 (g16371));
AN4X1 gate16875(.O (g19092), .I1 (g14776), .I2 (g18670), .I3 (g18692), .I4 (g16293));
AN2X1 gate16876(.O (g19093), .I1 (g17218), .I2 (g16572));
AN4X1 gate16877(.O (g19094), .I1 (g18679), .I2 (g14849), .I3 (g16254), .I4 (g13756));
AN4X1 gate16878(.O (g19095), .I1 (g14922), .I2 (g18765), .I3 (g16266), .I4 (g16313));
AN3X1 gate16879(.O (I25280), .I1 (g18656), .I2 (g18670), .I3 (g18720));
AN3X1 gate16880(.O (g19097), .I1 (g13657), .I2 (g16243), .I3 (I25280));
AN4X1 gate16881(.O (g19099), .I1 (g14811), .I2 (g18699), .I3 (g18728), .I4 (g16351));
AN2X1 gate16882(.O (g19100), .I1 (g17220), .I2 (g16596));
AN4X1 gate16883(.O (g19101), .I1 (g18708), .I2 (g14922), .I3 (g16313), .I4 (g13797));
AN4X1 gate16884(.O (g19102), .I1 (g15003), .I2 (g18796), .I3 (g16325), .I4 (g16371));
AN3X1 gate16885(.O (I25291), .I1 (g18679), .I2 (g18699), .I3 (g18758));
AN3X1 gate16886(.O (g19104), .I1 (g13687), .I2 (g16302), .I3 (I25291));
AN4X1 gate16887(.O (g19106), .I1 (g14863), .I2 (g18735), .I3 (g18765), .I4 (g16395));
AN2X1 gate16888(.O (g19107), .I1 (g17223), .I2 (g16616));
AN4X1 gate16889(.O (g19108), .I1 (g18744), .I2 (g15003), .I3 (g16371), .I4 (g13825));
AN3X1 gate16890(.O (I25300), .I1 (g18708), .I2 (g18735), .I3 (g18789));
AN3X1 gate16891(.O (g19109), .I1 (g13724), .I2 (g16360), .I3 (I25300));
AN4X1 gate16892(.O (g19111), .I1 (g14936), .I2 (g18772), .I3 (g18796), .I4 (g16433));
AN2X1 gate16893(.O (g19112), .I1 (g14657), .I2 (g16633));
AN3X1 gate16894(.O (I25311), .I1 (g18744), .I2 (g18772), .I3 (g18815));
AN3X1 gate16895(.O (g19116), .I1 (g13774), .I2 (g16404), .I3 (I25311));
AN2X1 gate16896(.O (g19117), .I1 (g14691), .I2 (g16644));
AN2X1 gate16897(.O (g19124), .I1 (g14725), .I2 (g16656));
AN2X1 gate16898(.O (g19131), .I1 (g14753), .I2 (g16673));
AN2X1 gate16899(.O (g19142), .I1 (g17159), .I2 (g16719));
AN2X1 gate16900(.O (g19143), .I1 (g17174), .I2 (g16761));
AN2X1 gate16901(.O (g19146), .I1 (g17191), .I2 (g16788));
AN2X1 gate16902(.O (g19148), .I1 (g17202), .I2 (g16817));
AN2X1 gate16903(.O (g19150), .I1 (g17189), .I2 (g8602));
AN2X1 gate16904(.O (g19155), .I1 (g17200), .I2 (g8614));
AN2X1 gate16905(.O (g19161), .I1 (g17207), .I2 (g8627));
AN2X1 gate16906(.O (g19166), .I1 (g17212), .I2 (g8637));
AN2X1 gate16907(.O (g19228), .I1 (g16662), .I2 (g12125));
AN2X1 gate16908(.O (g19236), .I1 (g16935), .I2 (g8802));
AN3X1 gate16909(.O (g19241), .I1 (g16867), .I2 (g14158), .I3 (g14071));
AN2X1 gate16910(.O (g19248), .I1 (g16662), .I2 (g8817));
AN2X1 gate16911(.O (g19252), .I1 (g18725), .I2 (g9527));
AN3X1 gate16912(.O (g19254), .I1 (g16895), .I2 (g14273), .I3 (g14186));
AN2X1 gate16913(.O (g19260), .I1 (g16749), .I2 (g3124));
AN3X1 gate16914(.O (g19267), .I1 (g16924), .I2 (g14395), .I3 (g14301));
AN3X1 gate16915(.O (g19282), .I1 (g16954), .I2 (g14507), .I3 (g14423));
AN2X1 gate16916(.O (g19284), .I1 (g18063), .I2 (g3111));
AN2X1 gate16917(.O (g19285), .I1 (g16749), .I2 (g7642));
AN2X1 gate16918(.O (g19289), .I1 (g17029), .I2 (g8580));
AN3X1 gate16919(.O (g19303), .I1 (g16867), .I2 (g16543), .I3 (g14071));
AN2X1 gate16920(.O (g19307), .I1 (g17063), .I2 (g8587));
AN2X1 gate16921(.O (g19316), .I1 (g18063), .I2 (g3110));
AN2X1 gate16922(.O (g19317), .I1 (g16749), .I2 (g3126));
AN3X1 gate16923(.O (g19320), .I1 (g16867), .I2 (g16515), .I3 (g14158));
AN3X1 gate16924(.O (g19324), .I1 (g16895), .I2 (g16575), .I3 (g14186));
AN2X1 gate16925(.O (g19328), .I1 (g17098), .I2 (g8594));
AN3X1 gate16926(.O (g19347), .I1 (g16895), .I2 (g16546), .I3 (g14273));
AN3X1 gate16927(.O (g19351), .I1 (g16924), .I2 (g16599), .I3 (g14301));
AN2X1 gate16928(.O (g19355), .I1 (g17136), .I2 (g8605));
AN2X1 gate16929(.O (g19356), .I1 (g18063), .I2 (g3112));
AN3X1 gate16930(.O (g19381), .I1 (g16924), .I2 (g16578), .I3 (g14395));
AN3X1 gate16931(.O (g19385), .I1 (g16954), .I2 (g16619), .I3 (g14423));
AN3X1 gate16932(.O (g19413), .I1 (g16954), .I2 (g16602), .I3 (g14507));
AN3X1 gate16933(.O (g19449), .I1 (g16884), .I2 (g14797), .I3 (g14776));
AN3X1 gate16934(.O (g19476), .I1 (g16913), .I2 (g14849), .I3 (g14811));
AN3X1 gate16935(.O (g19499), .I1 (g16943), .I2 (g14922), .I3 (g14863));
AN3X1 gate16936(.O (g19520), .I1 (g16974), .I2 (g15003), .I3 (g14936));
AN3X1 gate16937(.O (g19531), .I1 (g16884), .I2 (g16722), .I3 (g14776));
AN3X1 gate16938(.O (g19540), .I1 (g16884), .I2 (g16697), .I3 (g14797));
AN3X1 gate16939(.O (g19541), .I1 (g16913), .I2 (g16764), .I3 (g14811));
AN3X1 gate16940(.O (g19544), .I1 (g16913), .I2 (g16728), .I3 (g14849));
AN3X1 gate16941(.O (g19545), .I1 (g16943), .I2 (g16791), .I3 (g14863));
AN3X1 gate16942(.O (g19547), .I1 (g16943), .I2 (g16770), .I3 (g14922));
AN3X1 gate16943(.O (g19548), .I1 (g16974), .I2 (g16820), .I3 (g14936));
AN2X1 gate16944(.O (g19549), .I1 (g7950), .I2 (g17230));
AN3X1 gate16945(.O (g19551), .I1 (g16974), .I2 (g16797), .I3 (g15003));
AN2X1 gate16946(.O (g19552), .I1 (g16829), .I2 (g6048));
AN2X1 gate16947(.O (g19553), .I1 (g7990), .I2 (g17237));
AN2X1 gate16948(.O (g19554), .I1 (g7993), .I2 (g17240));
AN2X1 gate16949(.O (g19555), .I1 (g8001), .I2 (g17243));
AN2X1 gate16950(.O (g19557), .I1 (g8053), .I2 (g17249));
AN2X1 gate16951(.O (g19558), .I1 (g8056), .I2 (g17252));
AN2X1 gate16952(.O (g19559), .I1 (g8059), .I2 (g17255));
AN2X1 gate16953(.O (g19560), .I1 (g8065), .I2 (g17259));
AN2X1 gate16954(.O (g19561), .I1 (g8068), .I2 (g17262));
AN2X1 gate16955(.O (g19562), .I1 (g8076), .I2 (g17265));
AN2X1 gate16956(.O (g19564), .I1 (g8123), .I2 (g17272));
AN2X1 gate16957(.O (g19565), .I1 (g8126), .I2 (g17275));
AN2X1 gate16958(.O (g19566), .I1 (g8129), .I2 (g17278));
AN2X1 gate16959(.O (g19567), .I1 (g8138), .I2 (g17282));
AN2X1 gate16960(.O (g19568), .I1 (g8141), .I2 (g17285));
AN2X1 gate16961(.O (g19569), .I1 (g8144), .I2 (g17288));
AN2X1 gate16962(.O (g19570), .I1 (g8150), .I2 (g17291));
AN2X1 gate16963(.O (g19571), .I1 (g8153), .I2 (g17294));
AN2X1 gate16964(.O (g19572), .I1 (g8161), .I2 (g17297));
AN2X1 gate16965(.O (g19574), .I1 (g8191), .I2 (g17304));
AN2X1 gate16966(.O (g19575), .I1 (g8194), .I2 (g17307));
AN2X1 gate16967(.O (g19576), .I1 (g8197), .I2 (g17310));
AN2X1 gate16968(.O (g19584), .I1 (g640), .I2 (g18756));
AN2X1 gate16969(.O (g19585), .I1 (g692), .I2 (g18757));
AN2X1 gate16970(.O (g19586), .I1 (g8209), .I2 (g17315));
AN2X1 gate16971(.O (g19587), .I1 (g8212), .I2 (g17318));
AN2X1 gate16972(.O (g19588), .I1 (g8215), .I2 (g17321));
AN2X1 gate16973(.O (g19589), .I1 (g8224), .I2 (g17324));
AN2X1 gate16974(.O (g19590), .I1 (g8227), .I2 (g17327));
AN2X1 gate16975(.O (g19591), .I1 (g8230), .I2 (g17330));
AN2X1 gate16976(.O (g19592), .I1 (g8236), .I2 (g17333));
AN2X1 gate16977(.O (g19593), .I1 (g8239), .I2 (g17336));
AN2X1 gate16978(.O (g19594), .I1 (g16935), .I2 (g12555));
AN2X1 gate16979(.O (g19597), .I1 (g3922), .I2 (g17342));
AN2X1 gate16980(.O (g19598), .I1 (g3925), .I2 (g17345));
AN2X1 gate16981(.O (g19599), .I1 (g3928), .I2 (g17348));
AN2X1 gate16982(.O (g19600), .I1 (g633), .I2 (g18783));
AN2X1 gate16983(.O (g19601), .I1 (g640), .I2 (g18784));
AN2X1 gate16984(.O (g19602), .I1 (g633), .I2 (g18785));
AN2X1 gate16985(.O (g19603), .I1 (g692), .I2 (g18786));
AN2X1 gate16986(.O (g19604), .I1 (g3948), .I2 (g17354));
AN2X1 gate16987(.O (g19605), .I1 (g3951), .I2 (g17357));
AN2X1 gate16988(.O (g19606), .I1 (g3954), .I2 (g17360));
AN2X1 gate16989(.O (g19614), .I1 (g1326), .I2 (g18787));
AN2X1 gate16990(.O (g19615), .I1 (g1378), .I2 (g18788));
AN2X1 gate16991(.O (g19616), .I1 (g3966), .I2 (g17363));
AN2X1 gate16992(.O (g19617), .I1 (g3969), .I2 (g17366));
AN2X1 gate16993(.O (g19618), .I1 (g3972), .I2 (g17369));
AN2X1 gate16994(.O (g19619), .I1 (g3981), .I2 (g17372));
AN2X1 gate16995(.O (g19620), .I1 (g3984), .I2 (g17375));
AN2X1 gate16996(.O (g19621), .I1 (g3987), .I2 (g17378));
AN2X1 gate16997(.O (g19623), .I1 (g4000), .I2 (g17384));
AN2X1 gate16998(.O (g19624), .I1 (g4003), .I2 (g17387));
AN2X1 gate16999(.O (g19625), .I1 (g4006), .I2 (g17390));
AN2X1 gate17000(.O (g19626), .I1 (g640), .I2 (g18805));
AN2X1 gate17001(.O (g19627), .I1 (g633), .I2 (g18806));
AN2X1 gate17002(.O (g19628), .I1 (g653), .I2 (g18807));
AN2X1 gate17003(.O (g19629), .I1 (g692), .I2 (g18808));
AN2X1 gate17004(.O (g19630), .I1 (g4029), .I2 (g17399));
AN2X1 gate17005(.O (g19631), .I1 (g4032), .I2 (g17402));
AN2X1 gate17006(.O (g19632), .I1 (g4035), .I2 (g17405));
AN2X1 gate17007(.O (g19633), .I1 (g1319), .I2 (g18809));
AN2X1 gate17008(.O (g19634), .I1 (g1326), .I2 (g18810));
AN2X1 gate17009(.O (g19635), .I1 (g1319), .I2 (g18811));
AN2X1 gate17010(.O (g19636), .I1 (g1378), .I2 (g18812));
AN2X1 gate17011(.O (g19637), .I1 (g4055), .I2 (g17410));
AN2X1 gate17012(.O (g19638), .I1 (g4058), .I2 (g17413));
AN2X1 gate17013(.O (g19639), .I1 (g4061), .I2 (g17416));
AN2X1 gate17014(.O (g19647), .I1 (g2020), .I2 (g18813));
AN2X1 gate17015(.O (g19648), .I1 (g2072), .I2 (g18814));
AN2X1 gate17016(.O (g19649), .I1 (g4073), .I2 (g17419));
AN2X1 gate17017(.O (g19650), .I1 (g4076), .I2 (g17422));
AN2X1 gate17018(.O (g19651), .I1 (g4079), .I2 (g17425));
AN2X1 gate17019(.O (g19653), .I1 (g4095), .I2 (g17430));
AN2X1 gate17020(.O (g19654), .I1 (g4098), .I2 (g17433));
AN2X1 gate17021(.O (g19655), .I1 (g4101), .I2 (g17436));
AN2X1 gate17022(.O (g19656), .I1 (g4104), .I2 (g17439));
AN2X1 gate17023(.O (g19660), .I1 (g633), .I2 (g18822));
AN2X1 gate17024(.O (g19661), .I1 (g653), .I2 (g18823));
AN2X1 gate17025(.O (g19662), .I1 (g646), .I2 (g18824));
AN2X1 gate17026(.O (g19663), .I1 (g4127), .I2 (g17451));
AN2X1 gate17027(.O (g19664), .I1 (g4130), .I2 (g17454));
AN2X1 gate17028(.O (g19665), .I1 (g4133), .I2 (g17457));
AN2X1 gate17029(.O (g19666), .I1 (g1326), .I2 (g18825));
AN2X1 gate17030(.O (g19667), .I1 (g1319), .I2 (g18826));
AN2X1 gate17031(.O (g19668), .I1 (g1339), .I2 (g18827));
AN2X1 gate17032(.O (g19669), .I1 (g1378), .I2 (g18828));
AN2X1 gate17033(.O (g19670), .I1 (g4156), .I2 (g17465));
AN2X1 gate17034(.O (g19671), .I1 (g4159), .I2 (g17468));
AN2X1 gate17035(.O (g19672), .I1 (g4162), .I2 (g17471));
AN2X1 gate17036(.O (g19673), .I1 (g2013), .I2 (g18829));
AN2X1 gate17037(.O (g19674), .I1 (g2020), .I2 (g18830));
AN2X1 gate17038(.O (g19675), .I1 (g2013), .I2 (g18831));
AN2X1 gate17039(.O (g19676), .I1 (g2072), .I2 (g18832));
AN2X1 gate17040(.O (g19677), .I1 (g4182), .I2 (g17476));
AN2X1 gate17041(.O (g19678), .I1 (g4185), .I2 (g17479));
AN2X1 gate17042(.O (g19679), .I1 (g4188), .I2 (g17482));
AN2X1 gate17043(.O (g19687), .I1 (g2714), .I2 (g18833));
AN2X1 gate17044(.O (g19688), .I1 (g2766), .I2 (g18834));
AN2X1 gate17045(.O (g19691), .I1 (g16841), .I2 (g10865));
AN2X1 gate17046(.O (g19692), .I1 (g4205), .I2 (g17487));
AN2X1 gate17047(.O (g19693), .I1 (g4208), .I2 (g17490));
AN2X1 gate17048(.O (g19694), .I1 (g4211), .I2 (g17493));
AN2X1 gate17049(.O (g19695), .I1 (g4214), .I2 (g17496));
AN2X1 gate17050(.O (g19697), .I1 (g653), .I2 (g18838));
AN2X1 gate17051(.O (g19698), .I1 (g646), .I2 (g18839));
AN2X1 gate17052(.O (g19699), .I1 (g660), .I2 (g18840));
AN2X1 gate17053(.O (g19700), .I1 (g17815), .I2 (g16024));
AN2X1 gate17054(.O (g19701), .I1 (g4234), .I2 (g17511));
AN2X1 gate17055(.O (g19702), .I1 (g4237), .I2 (g17514));
AN2X1 gate17056(.O (g19703), .I1 (g4240), .I2 (g17517));
AN2X1 gate17057(.O (g19704), .I1 (g4243), .I2 (g17520));
AN2X1 gate17058(.O (g19708), .I1 (g1319), .I2 (g18841));
AN2X1 gate17059(.O (g19709), .I1 (g1339), .I2 (g18842));
AN2X1 gate17060(.O (g19710), .I1 (g1332), .I2 (g18843));
AN2X1 gate17061(.O (g19711), .I1 (g4266), .I2 (g17531));
AN2X1 gate17062(.O (g19712), .I1 (g4269), .I2 (g17534));
AN2X1 gate17063(.O (g19713), .I1 (g4272), .I2 (g17537));
AN2X1 gate17064(.O (g19714), .I1 (g2020), .I2 (g18844));
AN2X1 gate17065(.O (g19715), .I1 (g2013), .I2 (g18845));
AN2X1 gate17066(.O (g19716), .I1 (g2033), .I2 (g18846));
AN2X1 gate17067(.O (g19717), .I1 (g2072), .I2 (g18847));
AN2X1 gate17068(.O (g19718), .I1 (g4295), .I2 (g17545));
AN2X1 gate17069(.O (g19719), .I1 (g4298), .I2 (g17548));
AN2X1 gate17070(.O (g19720), .I1 (g4301), .I2 (g17551));
AN2X1 gate17071(.O (g19721), .I1 (g2707), .I2 (g18848));
AN2X1 gate17072(.O (g19722), .I1 (g2714), .I2 (g18849));
AN2X1 gate17073(.O (g19723), .I1 (g2707), .I2 (g18850));
AN2X1 gate17074(.O (g19724), .I1 (g2766), .I2 (g18851));
AN2X1 gate17075(.O (g19726), .I1 (g16847), .I2 (g6131));
AN2X1 gate17076(.O (g19727), .I1 (g4329), .I2 (g17557));
AN2X1 gate17077(.O (g19728), .I1 (g4332), .I2 (g17560));
AN2X1 gate17078(.O (g19729), .I1 (g4335), .I2 (g17563));
AN2X1 gate17079(.O (g19730), .I1 (g653), .I2 (g17573));
AN2X1 gate17080(.O (g19731), .I1 (g646), .I2 (g18853));
AN2X1 gate17081(.O (g19732), .I1 (g660), .I2 (g18854));
AN2X1 gate17082(.O (g19733), .I1 (g672), .I2 (g18855));
AN2X1 gate17083(.O (g19734), .I1 (g17815), .I2 (g16034));
AN2X1 gate17084(.O (g19735), .I1 (g17903), .I2 (g16035));
AN2X1 gate17085(.O (g19736), .I1 (g4360), .I2 (g17579));
AN2X1 gate17086(.O (g19737), .I1 (g4363), .I2 (g17582));
AN2X1 gate17087(.O (g19738), .I1 (g4366), .I2 (g17585));
AN2X1 gate17088(.O (g19739), .I1 (g4369), .I2 (g17588));
AN2X1 gate17089(.O (g19741), .I1 (g1339), .I2 (g18856));
AN2X1 gate17090(.O (g19742), .I1 (g1332), .I2 (g18857));
AN2X1 gate17091(.O (g19743), .I1 (g1346), .I2 (g18858));
AN2X1 gate17092(.O (g19744), .I1 (g17927), .I2 (g16040));
AN2X1 gate17093(.O (g19745), .I1 (g4389), .I2 (g17601));
AN2X1 gate17094(.O (g19746), .I1 (g4392), .I2 (g17604));
AN2X1 gate17095(.O (g19747), .I1 (g4395), .I2 (g17607));
AN2X1 gate17096(.O (g19748), .I1 (g4398), .I2 (g17610));
AN2X1 gate17097(.O (g19752), .I1 (g2013), .I2 (g18859));
AN2X1 gate17098(.O (g19753), .I1 (g2033), .I2 (g18860));
AN2X1 gate17099(.O (g19754), .I1 (g2026), .I2 (g18861));
AN2X1 gate17100(.O (g19755), .I1 (g4421), .I2 (g17621));
AN2X1 gate17101(.O (g19756), .I1 (g4424), .I2 (g17624));
AN2X1 gate17102(.O (g19757), .I1 (g4427), .I2 (g17627));
AN2X1 gate17103(.O (g19758), .I1 (g2714), .I2 (g18862));
AN2X1 gate17104(.O (g19759), .I1 (g2707), .I2 (g18863));
AN2X1 gate17105(.O (g19760), .I1 (g2727), .I2 (g18864));
AN2X1 gate17106(.O (g19761), .I1 (g2766), .I2 (g18865));
AN2X1 gate17107(.O (g19764), .I1 (g4453), .I2 (g17637));
AN2X1 gate17108(.O (g19765), .I1 (g660), .I2 (g18870));
AN2X1 gate17109(.O (g19766), .I1 (g672), .I2 (g18871));
AN2X1 gate17110(.O (g19767), .I1 (g666), .I2 (g18872));
AN2X1 gate17111(.O (g19768), .I1 (g17815), .I2 (g16054));
AN2X1 gate17112(.O (g19769), .I1 (g17903), .I2 (g16055));
AN2X1 gate17113(.O (g19770), .I1 (g4498), .I2 (g17655));
AN2X1 gate17114(.O (g19771), .I1 (g4501), .I2 (g17658));
AN2X1 gate17115(.O (g19772), .I1 (g4504), .I2 (g17661));
AN2X1 gate17116(.O (g19773), .I1 (g1339), .I2 (g17670));
AN2X1 gate17117(.O (g19774), .I1 (g1332), .I2 (g18874));
AN2X1 gate17118(.O (g19775), .I1 (g1346), .I2 (g18875));
AN2X1 gate17119(.O (g19776), .I1 (g1358), .I2 (g18876));
AN2X1 gate17120(.O (g19777), .I1 (g17927), .I2 (g16056));
AN2X1 gate17121(.O (g19778), .I1 (g18014), .I2 (g16057));
AN2X1 gate17122(.O (g19779), .I1 (g4529), .I2 (g17676));
AN2X1 gate17123(.O (g19780), .I1 (g4532), .I2 (g17679));
AN2X1 gate17124(.O (g19781), .I1 (g4535), .I2 (g17682));
AN2X1 gate17125(.O (g19782), .I1 (g4538), .I2 (g17685));
AN2X1 gate17126(.O (g19784), .I1 (g2033), .I2 (g18877));
AN2X1 gate17127(.O (g19785), .I1 (g2026), .I2 (g18878));
AN2X1 gate17128(.O (g19786), .I1 (g2040), .I2 (g18879));
AN2X1 gate17129(.O (g19787), .I1 (g18038), .I2 (g16062));
AN2X1 gate17130(.O (g19788), .I1 (g4558), .I2 (g17698));
AN2X1 gate17131(.O (g19789), .I1 (g4561), .I2 (g17701));
AN2X1 gate17132(.O (g19790), .I1 (g4564), .I2 (g17704));
AN2X1 gate17133(.O (g19791), .I1 (g4567), .I2 (g17707));
AN2X1 gate17134(.O (g19795), .I1 (g2707), .I2 (g18880));
AN2X1 gate17135(.O (g19796), .I1 (g2727), .I2 (g18881));
AN2X1 gate17136(.O (g19797), .I1 (g2720), .I2 (g18882));
AN3X1 gate17137(.O (I26240), .I1 (g18174), .I2 (g18341), .I3 (g17974));
AN3X1 gate17138(.O (g19799), .I1 (g17640), .I2 (g18074), .I3 (I26240));
AN2X1 gate17139(.O (g19802), .I1 (g672), .I2 (g18891));
AN2X1 gate17140(.O (g19803), .I1 (g666), .I2 (g18892));
AN2X1 gate17141(.O (g19804), .I1 (g679), .I2 (g18893));
AN2X1 gate17142(.O (g19805), .I1 (g17903), .I2 (g16088));
AN2X1 gate17143(.O (g19806), .I1 (g4629), .I2 (g17738));
AN2X1 gate17144(.O (g19807), .I1 (g1346), .I2 (g18896));
AN2X1 gate17145(.O (g19808), .I1 (g1358), .I2 (g18897));
AN2X1 gate17146(.O (g19809), .I1 (g1352), .I2 (g18898));
AN2X1 gate17147(.O (g19810), .I1 (g17927), .I2 (g16090));
AN2X1 gate17148(.O (g19811), .I1 (g18014), .I2 (g16091));
AN2X1 gate17149(.O (g19812), .I1 (g4674), .I2 (g17755));
AN2X1 gate17150(.O (g19813), .I1 (g4677), .I2 (g17758));
AN2X1 gate17151(.O (g19814), .I1 (g4680), .I2 (g17761));
AN2X1 gate17152(.O (g19815), .I1 (g2033), .I2 (g17770));
AN2X1 gate17153(.O (g19816), .I1 (g2026), .I2 (g18900));
AN2X1 gate17154(.O (g19817), .I1 (g2040), .I2 (g18901));
AN2X1 gate17155(.O (g19818), .I1 (g2052), .I2 (g18902));
AN2X1 gate17156(.O (g19819), .I1 (g18038), .I2 (g16092));
AN2X1 gate17157(.O (g19820), .I1 (g18131), .I2 (g16093));
AN2X1 gate17158(.O (g19821), .I1 (g4705), .I2 (g17776));
AN2X1 gate17159(.O (g19822), .I1 (g4708), .I2 (g17779));
AN2X1 gate17160(.O (g19823), .I1 (g4711), .I2 (g17782));
AN2X1 gate17161(.O (g19824), .I1 (g4714), .I2 (g17785));
AN2X1 gate17162(.O (g19826), .I1 (g2727), .I2 (g18903));
AN2X1 gate17163(.O (g19827), .I1 (g2720), .I2 (g18904));
AN2X1 gate17164(.O (g19828), .I1 (g2734), .I2 (g18905));
AN2X1 gate17165(.O (g19829), .I1 (g18155), .I2 (g16098));
AN2X1 gate17166(.O (g19836), .I1 (g7143), .I2 (g18908));
AN2X1 gate17167(.O (g19837), .I1 (g6901), .I2 (g17799));
AN2X1 gate17168(.O (g19839), .I1 (g666), .I2 (g18909));
AN2X1 gate17169(.O (g19840), .I1 (g679), .I2 (g18910));
AN2X1 gate17170(.O (g19841), .I1 (g686), .I2 (g18911));
AN3X1 gate17171(.O (I26282), .I1 (g18188), .I2 (g18089), .I3 (g17991));
AN3X1 gate17172(.O (g19842), .I1 (g14525), .I2 (g13922), .I3 (I26282));
AN3X1 gate17173(.O (I26285), .I1 (g18281), .I2 (g18436), .I3 (g18091));
AN3X1 gate17174(.O (g19843), .I1 (g17741), .I2 (g18190), .I3 (I26285));
AN2X1 gate17175(.O (g19846), .I1 (g1358), .I2 (g18914));
AN2X1 gate17176(.O (g19847), .I1 (g1352), .I2 (g18915));
AN2X1 gate17177(.O (g19848), .I1 (g1365), .I2 (g18916));
AN2X1 gate17178(.O (g19849), .I1 (g18014), .I2 (g16126));
AN2X1 gate17179(.O (g19850), .I1 (g4806), .I2 (g17839));
AN2X1 gate17180(.O (g19851), .I1 (g2040), .I2 (g18919));
AN2X1 gate17181(.O (g19852), .I1 (g2052), .I2 (g18920));
AN2X1 gate17182(.O (g19853), .I1 (g2046), .I2 (g18921));
AN2X1 gate17183(.O (g19854), .I1 (g18038), .I2 (g16128));
AN2X1 gate17184(.O (g19855), .I1 (g18131), .I2 (g16129));
AN2X1 gate17185(.O (g19856), .I1 (g4851), .I2 (g17856));
AN2X1 gate17186(.O (g19857), .I1 (g4854), .I2 (g17859));
AN2X1 gate17187(.O (g19858), .I1 (g4857), .I2 (g17862));
AN2X1 gate17188(.O (g19859), .I1 (g2727), .I2 (g17871));
AN2X1 gate17189(.O (g19860), .I1 (g2720), .I2 (g18923));
AN2X1 gate17190(.O (g19861), .I1 (g2734), .I2 (g18924));
AN2X1 gate17191(.O (g19862), .I1 (g2746), .I2 (g18925));
AN2X1 gate17192(.O (g19863), .I1 (g18155), .I2 (g16130));
AN2X1 gate17193(.O (g19864), .I1 (g18247), .I2 (g16131));
AN3X1 gate17194(.O (g19868), .I1 (g16498), .I2 (g16867), .I3 (g19001));
AN2X1 gate17195(.O (g19869), .I1 (g679), .I2 (g18926));
AN2X1 gate17196(.O (g19870), .I1 (g686), .I2 (g18927));
AN3X1 gate17197(.O (I26311), .I1 (g18353), .I2 (g13958), .I3 (g14011));
AN3X1 gate17198(.O (g19871), .I1 (g14086), .I2 (g18275), .I3 (I26311));
AN2X1 gate17199(.O (g19872), .I1 (g1352), .I2 (g18928));
AN2X1 gate17200(.O (g19873), .I1 (g1365), .I2 (g18929));
AN2X1 gate17201(.O (g19874), .I1 (g1372), .I2 (g18930));
AN3X1 gate17202(.O (I26317), .I1 (g18295), .I2 (g18205), .I3 (g18108));
AN3X1 gate17203(.O (g19875), .I1 (g14580), .I2 (g13978), .I3 (I26317));
AN3X1 gate17204(.O (I26320), .I1 (g18374), .I2 (g18509), .I3 (g18207));
AN3X1 gate17205(.O (g19876), .I1 (g17842), .I2 (g18297), .I3 (I26320));
AN2X1 gate17206(.O (g19879), .I1 (g2052), .I2 (g18933));
AN2X1 gate17207(.O (g19880), .I1 (g2046), .I2 (g18934));
AN2X1 gate17208(.O (g19881), .I1 (g2059), .I2 (g18935));
AN2X1 gate17209(.O (g19882), .I1 (g18131), .I2 (g16177));
AN2X1 gate17210(.O (g19883), .I1 (g4982), .I2 (g17951));
AN2X1 gate17211(.O (g19884), .I1 (g2734), .I2 (g18938));
AN2X1 gate17212(.O (g19885), .I1 (g2746), .I2 (g18939));
AN2X1 gate17213(.O (g19886), .I1 (g2740), .I2 (g18940));
AN2X1 gate17214(.O (g19887), .I1 (g18155), .I2 (g16179));
AN2X1 gate17215(.O (g19888), .I1 (g18247), .I2 (g16180));
AN2X1 gate17216(.O (g19889), .I1 (g2912), .I2 (g18943));
AN2X1 gate17217(.O (g19895), .I1 (g686), .I2 (g18945));
AN3X1 gate17218(.O (g19899), .I1 (g16520), .I2 (g16895), .I3 (g16507));
AN2X1 gate17219(.O (g19900), .I1 (g1365), .I2 (g18946));
AN2X1 gate17220(.O (g19901), .I1 (g1372), .I2 (g18947));
AN3X1 gate17221(.O (I26348), .I1 (g18448), .I2 (g14028), .I3 (g14102));
AN3X1 gate17222(.O (g19902), .I1 (g14201), .I2 (g18368), .I3 (I26348));
AN2X1 gate17223(.O (g19903), .I1 (g2046), .I2 (g18948));
AN2X1 gate17224(.O (g19904), .I1 (g2059), .I2 (g18949));
AN2X1 gate17225(.O (g19905), .I1 (g2066), .I2 (g18950));
AN3X1 gate17226(.O (I26354), .I1 (g18388), .I2 (g18312), .I3 (g18224));
AN3X1 gate17227(.O (g19906), .I1 (g14614), .I2 (g14048), .I3 (I26354));
AN3X1 gate17228(.O (I26357), .I1 (g18469), .I2 (g18573), .I3 (g18314));
AN3X1 gate17229(.O (g19907), .I1 (g17954), .I2 (g18390), .I3 (I26357));
AN2X1 gate17230(.O (g19910), .I1 (g2746), .I2 (g18953));
AN2X1 gate17231(.O (g19911), .I1 (g2740), .I2 (g18954));
AN2X1 gate17232(.O (g19912), .I1 (g2753), .I2 (g18955));
AN2X1 gate17233(.O (g19913), .I1 (g18247), .I2 (g16236));
AN2X1 gate17234(.O (g19914), .I1 (g3018), .I2 (g18958));
AN2X1 gate17235(.O (g19920), .I1 (g1372), .I2 (g18961));
AN3X1 gate17236(.O (g19924), .I1 (g16551), .I2 (g16924), .I3 (g16529));
AN2X1 gate17237(.O (g19925), .I1 (g2059), .I2 (g18962));
AN2X1 gate17238(.O (g19926), .I1 (g2066), .I2 (g18963));
AN3X1 gate17239(.O (I26377), .I1 (g18521), .I2 (g14119), .I3 (g14217));
AN3X1 gate17240(.O (g19927), .I1 (g14316), .I2 (g18463), .I3 (I26377));
AN2X1 gate17241(.O (g19928), .I1 (g2740), .I2 (g18964));
AN2X1 gate17242(.O (g19929), .I1 (g2753), .I2 (g18965));
AN2X1 gate17243(.O (g19930), .I1 (g2760), .I2 (g18966));
AN3X1 gate17244(.O (I26383), .I1 (g18483), .I2 (g18405), .I3 (g18331));
AN3X1 gate17245(.O (g19931), .I1 (g14637), .I2 (g14139), .I3 (I26383));
AN2X1 gate17246(.O (g19932), .I1 (g2917), .I2 (g18166));
AN2X1 gate17247(.O (g19935), .I1 (g2066), .I2 (g18972));
AN3X1 gate17248(.O (g19939), .I1 (g16583), .I2 (g16954), .I3 (g16560));
AN2X1 gate17249(.O (g19940), .I1 (g2753), .I2 (g18973));
AN2X1 gate17250(.O (g19941), .I1 (g2760), .I2 (g18974));
AN3X1 gate17251(.O (I26396), .I1 (g18585), .I2 (g14234), .I3 (g14332));
AN3X1 gate17252(.O (g19942), .I1 (g14438), .I2 (g18536), .I3 (I26396));
AN2X1 gate17253(.O (g19943), .I1 (g7562), .I2 (g18976));
AN2X1 gate17254(.O (g19944), .I1 (g3028), .I2 (g18258));
AN2X1 gate17255(.O (g19949), .I1 (g5293), .I2 (g18278));
AN2X1 gate17256(.O (g19952), .I1 (g2760), .I2 (g18987));
AN2X1 gate17257(.O (g19953), .I1 (g7566), .I2 (g18334));
AN3X1 gate17258(.O (I26416), .I1 (g18553), .I2 (g18491), .I3 (g18431));
AN3X1 gate17259(.O (g19970), .I1 (g18354), .I2 (g18276), .I3 (I26416));
AN2X1 gate17260(.O (g19971), .I1 (g5327), .I2 (g18355));
AN2X1 gate17261(.O (g19976), .I1 (g5330), .I2 (g18371));
AN3X1 gate17262(.O (I26432), .I1 (g18277), .I2 (g18189), .I3 (g18090));
AN3X1 gate17263(.O (g19982), .I1 (g17992), .I2 (g17913), .I3 (I26432));
AN2X1 gate17264(.O (g19983), .I1 (g5352), .I2 (g18432));
AN3X1 gate17265(.O (I26440), .I1 (g18603), .I2 (g18555), .I3 (g18504));
AN3X1 gate17266(.O (g20000), .I1 (g18449), .I2 (g18369), .I3 (I26440));
AN2X1 gate17267(.O (g20001), .I1 (g5355), .I2 (g18450));
AN2X1 gate17268(.O (g20006), .I1 (g5358), .I2 (g18466));
AN2X1 gate17269(.O (g20011), .I1 (g18063), .I2 (g3113));
AN2X1 gate17270(.O (g20012), .I1 (g16804), .I2 (g3135));
AN2X1 gate17271(.O (g20013), .I1 (g17720), .I2 (g12848));
AN2X1 gate17272(.O (g20014), .I1 (g7615), .I2 (g16749));
AN3X1 gate17273(.O (I26464), .I1 (g18370), .I2 (g18296), .I3 (g18206));
AN3X1 gate17274(.O (g20020), .I1 (g18109), .I2 (g18024), .I3 (I26464));
AN2X1 gate17275(.O (g20021), .I1 (g5369), .I2 (g18505));
AN3X1 gate17276(.O (I26472), .I1 (g18635), .I2 (g18605), .I3 (g18568));
AN3X1 gate17277(.O (g20038), .I1 (g18522), .I2 (g18464), .I3 (I26472));
AN2X1 gate17278(.O (g20039), .I1 (g5372), .I2 (g18523));
AN2X1 gate17279(.O (g20044), .I1 (g5375), .I2 (g18539));
AN2X1 gate17280(.O (g20048), .I1 (g16749), .I2 (g3127));
AN2X1 gate17281(.O (g20049), .I1 (g17878), .I2 (g3155));
AN2X1 gate17282(.O (g20050), .I1 (g18070), .I2 (g3161));
AN2X1 gate17283(.O (g20051), .I1 (g18063), .I2 (g3114));
AN2X1 gate17284(.O (g20052), .I1 (g16804), .I2 (g3134));
AN2X1 gate17285(.O (g20053), .I1 (g17720), .I2 (g12875));
AN3X1 gate17286(.O (I26500), .I1 (g18465), .I2 (g18389), .I3 (g18313));
AN3X1 gate17287(.O (g20062), .I1 (g18225), .I2 (g18141), .I3 (I26500));
AN2X1 gate17288(.O (g20063), .I1 (g5382), .I2 (g18569));
AN3X1 gate17289(.O (I26508), .I1 (g18644), .I2 (g18637), .I3 (g18618));
AN3X1 gate17290(.O (g20080), .I1 (g18586), .I2 (g18537), .I3 (I26508));
AN2X1 gate17291(.O (g20081), .I1 (g5385), .I2 (g18587));
AN2X1 gate17292(.O (g20084), .I1 (g17969), .I2 (g3158));
AN2X1 gate17293(.O (g20085), .I1 (g18170), .I2 (g3164));
AN2X1 gate17294(.O (g20086), .I1 (g18337), .I2 (g3170));
AN2X1 gate17295(.O (g20087), .I1 (g16749), .I2 (g7574));
AN2X1 gate17296(.O (g20088), .I1 (g16836), .I2 (g3147));
AN2X1 gate17297(.O (g20089), .I1 (g17969), .I2 (g9160));
AN2X1 gate17298(.O (g20090), .I1 (g18063), .I2 (g3120));
AN2X1 gate17299(.O (g20091), .I1 (g16804), .I2 (g3136));
AN2X1 gate17300(.O (g20092), .I1 (g16749), .I2 (g7603));
AN3X1 gate17301(.O (I26525), .I1 (g18656), .I2 (g18670), .I3 (g18692));
AN4X1 gate17302(.O (g20093), .I1 (g13657), .I2 (g13677), .I3 (g13750), .I4 (I26525));
AN3X1 gate17303(.O (I26528), .I1 (g18656), .I2 (g14837), .I3 (g13657));
AN3X1 gate17304(.O (g20094), .I1 (g13677), .I2 (g13706), .I3 (I26528));
AN3X1 gate17305(.O (I26541), .I1 (g18538), .I2 (g18484), .I3 (g18406));
AN3X1 gate17306(.O (g20103), .I1 (g18332), .I2 (g18257), .I3 (I26541));
AN2X1 gate17307(.O (g20104), .I1 (g5391), .I2 (g18619));
AN2X1 gate17308(.O (g20106), .I1 (g18261), .I2 (g3167));
AN2X1 gate17309(.O (g20107), .I1 (g18415), .I2 (g3173));
AN2X1 gate17310(.O (g20108), .I1 (g18543), .I2 (g3179));
AN2X1 gate17311(.O (g20109), .I1 (g17878), .I2 (g9504));
AN2X1 gate17312(.O (g20110), .I1 (g18070), .I2 (g9286));
AN2X1 gate17313(.O (g20111), .I1 (g18261), .I2 (g9884));
AN2X1 gate17314(.O (g20112), .I1 (g16749), .I2 (g3132));
AN2X1 gate17315(.O (g20113), .I1 (g16836), .I2 (g3142));
AN2X1 gate17316(.O (g20114), .I1 (g17969), .I2 (g9755));
AN2X1 gate17317(.O (g20115), .I1 (g16804), .I2 (g3139));
AN3X1 gate17318(.O (I26558), .I1 (g14776), .I2 (g18670), .I3 (g18720));
AN4X1 gate17319(.O (g20116), .I1 (g16142), .I2 (g13677), .I3 (g13706), .I4 (I26558));
AN3X1 gate17320(.O (I26561), .I1 (g14776), .I2 (g18720), .I3 (g13657));
AN3X1 gate17321(.O (g20117), .I1 (g16189), .I2 (g13706), .I3 (I26561));
AN3X1 gate17322(.O (I26564), .I1 (g18679), .I2 (g18699), .I3 (g18728));
AN4X1 gate17323(.O (g20118), .I1 (g13687), .I2 (g13714), .I3 (g13791), .I4 (I26564));
AN3X1 gate17324(.O (I26567), .I1 (g18679), .I2 (g14910), .I3 (g13687));
AN3X1 gate17325(.O (g20119), .I1 (g13714), .I2 (g13756), .I3 (I26567));
AN2X1 gate17326(.O (g20131), .I1 (g18486), .I2 (g3176));
AN2X1 gate17327(.O (g20132), .I1 (g18593), .I2 (g3182));
AN2X1 gate17328(.O (g20133), .I1 (g18170), .I2 (g9505));
AN2X1 gate17329(.O (g20134), .I1 (g18337), .I2 (g9506));
AN2X1 gate17330(.O (g20135), .I1 (g18486), .I2 (g9885));
AN2X1 gate17331(.O (g20136), .I1 (g17878), .I2 (g9423));
AN2X1 gate17332(.O (g20137), .I1 (g18070), .I2 (g9226));
AN2X1 gate17333(.O (g20138), .I1 (g18261), .I2 (g9756));
AN2X1 gate17334(.O (g20139), .I1 (g16836), .I2 (g3151));
AN3X1 gate17335(.O (g20144), .I1 (g16679), .I2 (g16884), .I3 (g16665));
AN4X1 gate17336(.O (g20145), .I1 (g14776), .I2 (g18670), .I3 (g16142), .I4 (g16189));
AN3X1 gate17337(.O (I26590), .I1 (g14811), .I2 (g18699), .I3 (g18758));
AN4X1 gate17338(.O (g20146), .I1 (g16201), .I2 (g13714), .I3 (g13756), .I4 (I26590));
AN3X1 gate17339(.O (I26593), .I1 (g14811), .I2 (g18758), .I3 (g13687));
AN3X1 gate17340(.O (g20147), .I1 (g16254), .I2 (g13756), .I3 (I26593));
AN3X1 gate17341(.O (I26596), .I1 (g18708), .I2 (g18735), .I3 (g18765));
AN4X1 gate17342(.O (g20148), .I1 (g13724), .I2 (g13764), .I3 (g13819), .I4 (I26596));
AN3X1 gate17343(.O (I26599), .I1 (g18708), .I2 (g14991), .I3 (g13724));
AN3X1 gate17344(.O (g20149), .I1 (g13764), .I2 (g13797), .I3 (I26599));
AN2X1 gate17345(.O (g20156), .I1 (g16809), .I2 (g3185));
AN2X1 gate17346(.O (g20157), .I1 (g18415), .I2 (g9287));
AN2X1 gate17347(.O (g20158), .I1 (g18543), .I2 (g9886));
AN2X1 gate17348(.O (g20159), .I1 (g16809), .I2 (g9288));
AN2X1 gate17349(.O (g20160), .I1 (g18170), .I2 (g9424));
AN2X1 gate17350(.O (g20161), .I1 (g18337), .I2 (g9426));
AN2X1 gate17351(.O (g20162), .I1 (g18486), .I2 (g9757));
AN3X1 gate17352(.O (I26615), .I1 (g14797), .I2 (g18692), .I3 (g13657));
AN3X1 gate17353(.O (g20177), .I1 (g13677), .I2 (g13750), .I3 (I26615));
AN3X1 gate17354(.O (g20182), .I1 (g16705), .I2 (g16913), .I3 (g16686));
AN4X1 gate17355(.O (g20183), .I1 (g14811), .I2 (g18699), .I3 (g16201), .I4 (g16254));
AN3X1 gate17356(.O (I26621), .I1 (g14863), .I2 (g18735), .I3 (g18789));
AN4X1 gate17357(.O (g20184), .I1 (g16266), .I2 (g13764), .I3 (g13797), .I4 (I26621));
AN3X1 gate17358(.O (I26624), .I1 (g14863), .I2 (g18789), .I3 (g13724));
AN3X1 gate17359(.O (g20185), .I1 (g16313), .I2 (g13797), .I3 (I26624));
AN3X1 gate17360(.O (I26627), .I1 (g18744), .I2 (g18772), .I3 (g18796));
AN4X1 gate17361(.O (g20186), .I1 (g13774), .I2 (g13805), .I3 (g13840), .I4 (I26627));
AN3X1 gate17362(.O (I26630), .I1 (g18744), .I2 (g15080), .I3 (g13774));
AN3X1 gate17363(.O (g20187), .I1 (g13805), .I2 (g13825), .I3 (I26630));
AN2X1 gate17364(.O (g20188), .I1 (g18593), .I2 (g9425));
AN2X1 gate17365(.O (g20189), .I1 (g16825), .I2 (g9289));
AN2X1 gate17366(.O (g20190), .I1 (g18415), .I2 (g9227));
AN2X1 gate17367(.O (g20191), .I1 (g18543), .I2 (g9758));
AN2X1 gate17368(.O (g20192), .I1 (g16809), .I2 (g9228));
AN3X1 gate17369(.O (I26639), .I1 (g18656), .I2 (g18670), .I3 (g16142));
AN3X1 gate17370(.O (g20197), .I1 (g13677), .I2 (g13706), .I3 (I26639));
AN3X1 gate17371(.O (I26645), .I1 (g14849), .I2 (g18728), .I3 (g13687));
AN3X1 gate17372(.O (g20211), .I1 (g13714), .I2 (g13791), .I3 (I26645));
AN3X1 gate17373(.O (g20216), .I1 (g16736), .I2 (g16943), .I3 (g16712));
AN4X1 gate17374(.O (g20217), .I1 (g14863), .I2 (g18735), .I3 (g16266), .I4 (g16313));
AN3X1 gate17375(.O (I26651), .I1 (g14936), .I2 (g18772), .I3 (g18815));
AN4X1 gate17376(.O (g20218), .I1 (g16325), .I2 (g13805), .I3 (g13825), .I4 (I26651));
AN3X1 gate17377(.O (I26654), .I1 (g14936), .I2 (g18815), .I3 (g13774));
AN3X1 gate17378(.O (g20219), .I1 (g16371), .I2 (g13825), .I3 (I26654));
AN2X1 gate17379(.O (g20220), .I1 (g18593), .I2 (g9355));
AN2X1 gate17380(.O (g20221), .I1 (g16825), .I2 (g10099));
AN4X1 gate17381(.O (g20222), .I1 (g18656), .I2 (g18720), .I3 (g13657), .I4 (g16293));
AN3X1 gate17382(.O (I26661), .I1 (g18679), .I2 (g18699), .I3 (g16201));
AN3X1 gate17383(.O (g20227), .I1 (g13714), .I2 (g13756), .I3 (I26661));
AN3X1 gate17384(.O (I26667), .I1 (g14922), .I2 (g18765), .I3 (g13724));
AN3X1 gate17385(.O (g20241), .I1 (g13764), .I2 (g13819), .I3 (I26667));
AN3X1 gate17386(.O (g20246), .I1 (g16778), .I2 (g16974), .I3 (g16743));
AN4X1 gate17387(.O (g20247), .I1 (g14936), .I2 (g18772), .I3 (g16325), .I4 (g16371));
AN3X1 gate17388(.O (g20248), .I1 (g18656), .I2 (g14837), .I3 (g16293));
AN4X1 gate17389(.O (g20249), .I1 (g18679), .I2 (g18758), .I3 (g13687), .I4 (g16351));
AN3X1 gate17390(.O (I26676), .I1 (g18708), .I2 (g18735), .I3 (g16266));
AN3X1 gate17391(.O (g20254), .I1 (g13764), .I2 (g13797), .I3 (I26676));
AN3X1 gate17392(.O (I26682), .I1 (g15003), .I2 (g18796), .I3 (g13774));
AN3X1 gate17393(.O (g20268), .I1 (g13805), .I2 (g13840), .I3 (I26682));
AN4X1 gate17394(.O (g20270), .I1 (g14797), .I2 (g18692), .I3 (g13657), .I4 (g16243));
AN3X1 gate17395(.O (g20271), .I1 (g18679), .I2 (g14910), .I3 (g16351));
AN4X1 gate17396(.O (g20272), .I1 (g18708), .I2 (g18789), .I3 (g13724), .I4 (g16395));
AN3X1 gate17397(.O (I26690), .I1 (g18744), .I2 (g18772), .I3 (g16325));
AN3X1 gate17398(.O (g20277), .I1 (g13805), .I2 (g13825), .I3 (I26690));
AN3X1 gate17399(.O (I26695), .I1 (g18670), .I2 (g18692), .I3 (g16142));
AN3X1 gate17400(.O (g20280), .I1 (g13677), .I2 (g16243), .I3 (I26695));
AN4X1 gate17401(.O (g20282), .I1 (g14849), .I2 (g18728), .I3 (g13687), .I4 (g16302));
AN3X1 gate17402(.O (g20283), .I1 (g18708), .I2 (g14991), .I3 (g16395));
AN4X1 gate17403(.O (g20284), .I1 (g18744), .I2 (g18815), .I3 (g13774), .I4 (g16433));
AN2X1 gate17404(.O (g20285), .I1 (g16846), .I2 (g8103));
AN3X1 gate17405(.O (I26708), .I1 (g18699), .I2 (g18728), .I3 (g16201));
AN3X1 gate17406(.O (g20291), .I1 (g13714), .I2 (g16302), .I3 (I26708));
AN4X1 gate17407(.O (g20293), .I1 (g14922), .I2 (g18765), .I3 (g13724), .I4 (g16360));
AN3X1 gate17408(.O (g20294), .I1 (g18744), .I2 (g15080), .I3 (g16433));
AN3X1 gate17409(.O (I26726), .I1 (g18735), .I2 (g18765), .I3 (g16266));
AN3X1 gate17410(.O (g20307), .I1 (g13764), .I2 (g16360), .I3 (I26726));
AN4X1 gate17411(.O (g20309), .I1 (g15003), .I2 (g18796), .I3 (g13774), .I4 (g16404));
AN3X1 gate17412(.O (I26745), .I1 (g18772), .I2 (g18796), .I3 (g16325));
AN3X1 gate17413(.O (g20326), .I1 (g13805), .I2 (g16404), .I3 (I26745));
AN2X1 gate17414(.O (g20460), .I1 (g17351), .I2 (g13644));
AN2X1 gate17415(.O (g20472), .I1 (g17314), .I2 (g13669));
AN2X1 gate17416(.O (g20480), .I1 (g17313), .I2 (g11827));
AN2X1 gate17417(.O (g20486), .I1 (g17281), .I2 (g11859));
AN2X1 gate17418(.O (g20492), .I1 (g17258), .I2 (g11894));
AN2X1 gate17419(.O (g20499), .I1 (g17648), .I2 (g11933));
AN2X1 gate17420(.O (g20502), .I1 (g17566), .I2 (g11973));
AN2X1 gate17421(.O (g20503), .I1 (g17507), .I2 (g13817));
AN2X1 gate17422(.O (g20506), .I1 (g17499), .I2 (g12025));
AN2X1 gate17423(.O (g20512), .I1 (g17445), .I2 (g13836));
AN2X1 gate17424(.O (g20525), .I1 (g17394), .I2 (g13849));
AN4X1 gate17425(.O (g20538), .I1 (g18656), .I2 (g14837), .I3 (g13657), .I4 (g16189));
AN2X1 gate17426(.O (g20640), .I1 (g4809), .I2 (g19064));
AN2X1 gate17427(.O (g20647), .I1 (g5888), .I2 (g19075));
AN2X1 gate17428(.O (g20665), .I1 (g4985), .I2 (g19081));
AN2X1 gate17429(.O (g20809), .I1 (g5712), .I2 (g19113));
AN2X1 gate17430(.O (g20826), .I1 (g5770), .I2 (g19118));
AN2X1 gate17431(.O (g20836), .I1 (g5829), .I2 (g19125));
AN2X1 gate17432(.O (g20840), .I1 (g5885), .I2 (g19132));
AN3X1 gate17433(.O (g21049), .I1 (g20016), .I2 (g14079), .I3 (g14165));
AN2X1 gate17434(.O (g21067), .I1 (g20193), .I2 (g12030));
AN3X1 gate17435(.O (g21068), .I1 (g20058), .I2 (g14194), .I3 (g14280));
AN2X1 gate17436(.O (g21077), .I1 (g20223), .I2 (g12094));
AN3X1 gate17437(.O (g21078), .I1 (g20099), .I2 (g14309), .I3 (g14402));
AN3X1 gate17438(.O (g21085), .I1 (g19484), .I2 (g14158), .I3 (g19001));
AN2X1 gate17439(.O (g21086), .I1 (g20193), .I2 (g12142));
AN2X1 gate17440(.O (g21091), .I1 (g20250), .I2 (g12166));
AN3X1 gate17441(.O (g21092), .I1 (g20124), .I2 (g14431), .I3 (g14514));
AN3X1 gate17442(.O (g21097), .I1 (g19505), .I2 (g14273), .I3 (g16507));
AN2X1 gate17443(.O (g21098), .I1 (g20223), .I2 (g12204));
AN2X1 gate17444(.O (g21103), .I1 (g20273), .I2 (g12228));
AN3X1 gate17445(.O (g21107), .I1 (g19444), .I2 (g17893), .I3 (g14079));
AN3X1 gate17446(.O (g21111), .I1 (g19524), .I2 (g14395), .I3 (g16529));
AN2X1 gate17447(.O (g21112), .I1 (g20250), .I2 (g12259));
AN2X1 gate17448(.O (g21121), .I1 (g20054), .I2 (g14244));
AN2X1 gate17449(.O (g21122), .I1 (g20140), .I2 (g12279));
AN2X1 gate17450(.O (g21123), .I1 (g19970), .I2 (g19982));
AN3X1 gate17451(.O (g21124), .I1 (g19471), .I2 (g18004), .I3 (g14194));
AN3X1 gate17452(.O (g21128), .I1 (g19534), .I2 (g14507), .I3 (g16560));
AN2X1 gate17453(.O (g21129), .I1 (g20273), .I2 (g12302));
AN3X1 gate17454(.O (I27695), .I1 (g19318), .I2 (g19300), .I3 (g19286));
AN3X1 gate17455(.O (g21136), .I1 (g19271), .I2 (g19261), .I3 (I27695));
AN2X1 gate17456(.O (g21137), .I1 (g5750), .I2 (g19272));
AN2X1 gate17457(.O (g21138), .I1 (g19484), .I2 (g14347));
AN2X1 gate17458(.O (g21140), .I1 (g20095), .I2 (g14366));
AN2X1 gate17459(.O (g21141), .I1 (g20178), .I2 (g12315));
AN2X1 gate17460(.O (g21142), .I1 (g20000), .I2 (g20020));
AN3X1 gate17461(.O (g21143), .I1 (g19494), .I2 (g18121), .I3 (g14309));
AN3X1 gate17462(.O (I27711), .I1 (g19262), .I2 (g19414), .I3 (g19386));
AN3X1 gate17463(.O (g21152), .I1 (g19357), .I2 (g19334), .I3 (I27711));
AN3X1 gate17464(.O (g21153), .I1 (g20054), .I2 (g16543), .I3 (g16501));
AN2X1 gate17465(.O (g21154), .I1 (g20193), .I2 (g12333));
AN2X1 gate17466(.O (g21155), .I1 (g20140), .I2 (g12336));
AN3X1 gate17467(.O (I27717), .I1 (g19345), .I2 (g19321), .I3 (g19304));
AN3X1 gate17468(.O (g21156), .I1 (g19290), .I2 (g19276), .I3 (I27717));
AN2X1 gate17469(.O (g21157), .I1 (g5809), .I2 (g19291));
AN2X1 gate17470(.O (g21158), .I1 (g19505), .I2 (g14459));
AN2X1 gate17471(.O (g21160), .I1 (g20120), .I2 (g14478));
AN2X1 gate17472(.O (g21161), .I1 (g20212), .I2 (g12343));
AN2X1 gate17473(.O (g21162), .I1 (g20038), .I2 (g20062));
AN3X1 gate17474(.O (g21163), .I1 (g19515), .I2 (g18237), .I3 (g14431));
AN3X1 gate17475(.O (I27733), .I1 (g19277), .I2 (g19451), .I3 (g19416));
AN3X1 gate17476(.O (g21172), .I1 (g19389), .I2 (g19368), .I3 (I27733));
AN3X1 gate17477(.O (g21173), .I1 (g20095), .I2 (g16575), .I3 (g16523));
AN2X1 gate17478(.O (g21174), .I1 (g20223), .I2 (g12363));
AN2X1 gate17479(.O (g21175), .I1 (g20178), .I2 (g12366));
AN3X1 gate17480(.O (I27739), .I1 (g19379), .I2 (g19348), .I3 (g19325));
AN3X1 gate17481(.O (g21176), .I1 (g19308), .I2 (g19295), .I3 (I27739));
AN2X1 gate17482(.O (g21177), .I1 (g5865), .I2 (g19309));
AN2X1 gate17483(.O (g21178), .I1 (g19524), .I2 (g14546));
AN2X1 gate17484(.O (g21180), .I1 (g20150), .I2 (g14565));
AN2X1 gate17485(.O (g21181), .I1 (g20242), .I2 (g12373));
AN2X1 gate17486(.O (g21182), .I1 (g20080), .I2 (g20103));
AN2X1 gate17487(.O (g21188), .I1 (g20140), .I2 (g12379));
AN3X1 gate17488(.O (I27755), .I1 (g19296), .I2 (g19478), .I3 (g19453));
AN3X1 gate17489(.O (g21192), .I1 (g19419), .I2 (g19400), .I3 (I27755));
AN3X1 gate17490(.O (g21193), .I1 (g20120), .I2 (g16599), .I3 (g16554));
AN2X1 gate17491(.O (g21194), .I1 (g20250), .I2 (g12382));
AN2X1 gate17492(.O (g21195), .I1 (g20212), .I2 (g12385));
AN3X1 gate17493(.O (I27761), .I1 (g19411), .I2 (g19382), .I3 (g19352));
AN3X1 gate17494(.O (g21196), .I1 (g19329), .I2 (g19313), .I3 (I27761));
AN2X1 gate17495(.O (g21197), .I1 (g5912), .I2 (g19330));
AN2X1 gate17496(.O (g21198), .I1 (g19534), .I2 (g14601));
AN2X1 gate17497(.O (g21203), .I1 (g20178), .I2 (g12409));
AN3X1 gate17498(.O (I27772), .I1 (g19314), .I2 (g19501), .I3 (g19480));
AN3X1 gate17499(.O (g21207), .I1 (g19456), .I2 (g19430), .I3 (I27772));
AN3X1 gate17500(.O (g21208), .I1 (g20150), .I2 (g16619), .I3 (g16586));
AN2X1 gate17501(.O (g21209), .I1 (g20273), .I2 (g12412));
AN2X1 gate17502(.O (g21210), .I1 (g20242), .I2 (g12415));
AN2X1 gate17503(.O (g21218), .I1 (g20212), .I2 (g12421));
AN2X1 gate17504(.O (g21226), .I1 (g20242), .I2 (g12426));
AN3X1 gate17505(.O (g21229), .I1 (g19578), .I2 (g14797), .I3 (g16665));
AN3X1 gate17506(.O (g21234), .I1 (g19608), .I2 (g14849), .I3 (g16686));
AN3X1 gate17507(.O (g21243), .I1 (g19641), .I2 (g14922), .I3 (g16712));
AN2X1 gate17508(.O (g21245), .I1 (g20299), .I2 (g14837));
AN3X1 gate17509(.O (g21251), .I1 (g19681), .I2 (g15003), .I3 (g16743));
AN2X1 gate17510(.O (g21252), .I1 (g19578), .I2 (g14895));
AN2X1 gate17511(.O (g21254), .I1 (g20318), .I2 (g14910));
AN3X1 gate17512(.O (g21259), .I1 (g20299), .I2 (g16722), .I3 (g16682));
AN2X1 gate17513(.O (g21260), .I1 (g19608), .I2 (g14976));
AN2X1 gate17514(.O (g21262), .I1 (g20337), .I2 (g14991));
AN3X1 gate17515(.O (g21267), .I1 (g20318), .I2 (g16764), .I3 (g16708));
AN2X1 gate17516(.O (g21268), .I1 (g19641), .I2 (g15065));
AN2X1 gate17517(.O (g21270), .I1 (g20357), .I2 (g15080));
AN3X1 gate17518(.O (g21276), .I1 (g20337), .I2 (g16791), .I3 (g16739));
AN2X1 gate17519(.O (g21277), .I1 (g19681), .I2 (g15161));
AN3X1 gate17520(.O (g21283), .I1 (g20357), .I2 (g16820), .I3 (g16781));
AN2X1 gate17521(.O (g21284), .I1 (g9356), .I2 (g20269));
AN2X1 gate17522(.O (g21290), .I1 (g9356), .I2 (g20278));
AN2X1 gate17523(.O (g21291), .I1 (g9293), .I2 (g20279));
AN2X1 gate17524(.O (g21292), .I1 (g9453), .I2 (g20281));
AN2X1 gate17525(.O (g21298), .I1 (g9356), .I2 (g20286));
AN2X1 gate17526(.O (g21299), .I1 (g9293), .I2 (g20287));
AN2X1 gate17527(.O (g21300), .I1 (g9232), .I2 (g20288));
AN2X1 gate17528(.O (g21301), .I1 (g9453), .I2 (g20289));
AN2X1 gate17529(.O (g21302), .I1 (g9374), .I2 (g20290));
AN2X1 gate17530(.O (g21303), .I1 (g9595), .I2 (g20292));
AN2X1 gate17531(.O (g21304), .I1 (g9293), .I2 (g20296));
AN2X1 gate17532(.O (g21305), .I1 (g9232), .I2 (g20297));
AN2X1 gate17533(.O (g21306), .I1 (g9187), .I2 (g20298));
AN2X1 gate17534(.O (g21307), .I1 (g9453), .I2 (g20302));
AN2X1 gate17535(.O (g21308), .I1 (g9374), .I2 (g20303));
AN2X1 gate17536(.O (g21309), .I1 (g9310), .I2 (g20304));
AN2X1 gate17537(.O (g21310), .I1 (g9595), .I2 (g20305));
AN2X1 gate17538(.O (g21311), .I1 (g9471), .I2 (g20306));
AN2X1 gate17539(.O (g21312), .I1 (g9737), .I2 (g20308));
AN2X1 gate17540(.O (g21313), .I1 (g9232), .I2 (g20311));
AN2X1 gate17541(.O (g21314), .I1 (g9187), .I2 (g20312));
AN2X1 gate17542(.O (g21315), .I1 (g9161), .I2 (g20313));
AN2X1 gate17543(.O (g21319), .I1 (g9374), .I2 (g20315));
AN2X1 gate17544(.O (g21320), .I1 (g9310), .I2 (g20316));
AN2X1 gate17545(.O (g21321), .I1 (g9248), .I2 (g20317));
AN2X1 gate17546(.O (g21322), .I1 (g9595), .I2 (g20321));
AN2X1 gate17547(.O (g21323), .I1 (g9471), .I2 (g20322));
AN2X1 gate17548(.O (g21324), .I1 (g9391), .I2 (g20323));
AN2X1 gate17549(.O (g21325), .I1 (g9737), .I2 (g20324));
AN2X1 gate17550(.O (g21326), .I1 (g9613), .I2 (g20325));
AN2X1 gate17551(.O (g21328), .I1 (g9187), .I2 (g20327));
AN2X1 gate17552(.O (g21329), .I1 (g9161), .I2 (g20328));
AN2X1 gate17553(.O (g21330), .I1 (g9150), .I2 (g20329));
AN2X1 gate17554(.O (g21334), .I1 (g9310), .I2 (g20330));
AN2X1 gate17555(.O (g21335), .I1 (g9248), .I2 (g20331));
AN2X1 gate17556(.O (g21336), .I1 (g9203), .I2 (g20332));
AN2X1 gate17557(.O (g21337), .I1 (g9471), .I2 (g20334));
AN2X1 gate17558(.O (g21338), .I1 (g9391), .I2 (g20335));
AN2X1 gate17559(.O (g21339), .I1 (g9326), .I2 (g20336));
AN2X1 gate17560(.O (g21340), .I1 (g9737), .I2 (g20340));
AN2X1 gate17561(.O (g21341), .I1 (g9613), .I2 (g20341));
AN2X1 gate17562(.O (g21342), .I1 (g9488), .I2 (g20342));
AN2X1 gate17563(.O (g21343), .I1 (g9161), .I2 (g20344));
AN2X1 gate17564(.O (g21344), .I1 (g9150), .I2 (g20345));
AN2X1 gate17565(.O (g21345), .I1 (g15096), .I2 (g20346));
AN2X1 gate17566(.O (g21349), .I1 (g9248), .I2 (g20347));
AN2X1 gate17567(.O (g21350), .I1 (g9203), .I2 (g20348));
AN2X1 gate17568(.O (g21351), .I1 (g9174), .I2 (g20349));
AN2X1 gate17569(.O (g21352), .I1 (g9391), .I2 (g20350));
AN2X1 gate17570(.O (g21353), .I1 (g9326), .I2 (g20351));
AN2X1 gate17571(.O (g21354), .I1 (g9264), .I2 (g20352));
AN2X1 gate17572(.O (g21355), .I1 (g9613), .I2 (g20354));
AN2X1 gate17573(.O (g21356), .I1 (g9488), .I2 (g20355));
AN2X1 gate17574(.O (g21357), .I1 (g9407), .I2 (g20356));
AN2X1 gate17575(.O (g21360), .I1 (g9507), .I2 (g20361));
AN2X1 gate17576(.O (g21361), .I1 (g9150), .I2 (g20362));
AN2X1 gate17577(.O (g21362), .I1 (g15096), .I2 (g20363));
AN2X1 gate17578(.O (g21363), .I1 (g15022), .I2 (g20364));
AN2X1 gate17579(.O (g21367), .I1 (g9203), .I2 (g20366));
AN2X1 gate17580(.O (g21368), .I1 (g9174), .I2 (g20367));
AN2X1 gate17581(.O (g21369), .I1 (g15188), .I2 (g20368));
AN2X1 gate17582(.O (g21370), .I1 (g9326), .I2 (g20369));
AN2X1 gate17583(.O (g21371), .I1 (g9264), .I2 (g20370));
AN2X1 gate17584(.O (g21372), .I1 (g9216), .I2 (g20371));
AN2X1 gate17585(.O (g21373), .I1 (g9488), .I2 (g20372));
AN2X1 gate17586(.O (g21374), .I1 (g9407), .I2 (g20373));
AN2X1 gate17587(.O (g21375), .I1 (g9342), .I2 (g20374));
AN2X1 gate17588(.O (g21378), .I1 (g9507), .I2 (g20378));
AN2X1 gate17589(.O (g21379), .I1 (g9427), .I2 (g20379));
AN2X1 gate17590(.O (g21380), .I1 (g15096), .I2 (g20380));
AN2X1 gate17591(.O (g21381), .I1 (g15022), .I2 (g20381));
AN2X1 gate17592(.O (g21388), .I1 (g6201), .I2 (g19657));
AN2X1 gate17593(.O (g21389), .I1 (g9649), .I2 (g20384));
AN2X1 gate17594(.O (g21390), .I1 (g9174), .I2 (g20385));
AN2X1 gate17595(.O (g21391), .I1 (g15188), .I2 (g20386));
AN2X1 gate17596(.O (g21392), .I1 (g15118), .I2 (g20387));
AN2X1 gate17597(.O (g21393), .I1 (g9264), .I2 (g20389));
AN2X1 gate17598(.O (g21394), .I1 (g9216), .I2 (g20390));
AN2X1 gate17599(.O (g21395), .I1 (g15274), .I2 (g20391));
AN2X1 gate17600(.O (g21396), .I1 (g9407), .I2 (g20392));
AN2X1 gate17601(.O (g21397), .I1 (g9342), .I2 (g20393));
AN2X1 gate17602(.O (g21398), .I1 (g9277), .I2 (g20394));
AN2X1 gate17603(.O (g21401), .I1 (g9507), .I2 (g20397));
AN2X1 gate17604(.O (g21402), .I1 (g9427), .I2 (g20398));
AN2X1 gate17605(.O (g21403), .I1 (g15022), .I2 (g20399));
AN2X1 gate17606(.O (g21410), .I1 (g6363), .I2 (g20402));
AN2X1 gate17607(.O (g21411), .I1 (g9649), .I2 (g20403));
AN2X1 gate17608(.O (g21412), .I1 (g9569), .I2 (g20404));
AN2X1 gate17609(.O (g21413), .I1 (g15188), .I2 (g20405));
AN2X1 gate17610(.O (g21414), .I1 (g15118), .I2 (g20406));
AN2X1 gate17611(.O (g21418), .I1 (g6290), .I2 (g19705));
AN2X1 gate17612(.O (g21419), .I1 (g9795), .I2 (g20409));
AN2X1 gate17613(.O (g21420), .I1 (g9216), .I2 (g20410));
AN2X1 gate17614(.O (g21421), .I1 (g15274), .I2 (g20411));
AN2X1 gate17615(.O (g21422), .I1 (g15210), .I2 (g20412));
AN2X1 gate17616(.O (g21423), .I1 (g9342), .I2 (g20414));
AN2X1 gate17617(.O (g21424), .I1 (g9277), .I2 (g20415));
AN2X1 gate17618(.O (g21425), .I1 (g15366), .I2 (g20416));
AN2X1 gate17619(.O (g21428), .I1 (g9427), .I2 (g20420));
AN2X1 gate17620(.O (g21438), .I1 (g9649), .I2 (g20422));
AN2X1 gate17621(.O (g21439), .I1 (g9569), .I2 (g20423));
AN2X1 gate17622(.O (g21440), .I1 (g15118), .I2 (g20424));
AN2X1 gate17623(.O (g21444), .I1 (g6568), .I2 (g20427));
AN2X1 gate17624(.O (g21445), .I1 (g9795), .I2 (g20428));
AN2X1 gate17625(.O (g21446), .I1 (g9711), .I2 (g20429));
AN2X1 gate17626(.O (g21447), .I1 (g15274), .I2 (g20430));
AN2X1 gate17627(.O (g21448), .I1 (g15210), .I2 (g20431));
AN2X1 gate17628(.O (g21452), .I1 (g6427), .I2 (g19749));
AN2X1 gate17629(.O (g21453), .I1 (g9941), .I2 (g20434));
AN2X1 gate17630(.O (g21454), .I1 (g9277), .I2 (g20435));
AN2X1 gate17631(.O (g21455), .I1 (g15366), .I2 (g20436));
AN2X1 gate17632(.O (g21456), .I1 (g15296), .I2 (g20437));
AN2X1 gate17633(.O (g21476), .I1 (g9569), .I2 (g20442));
AN2X1 gate17634(.O (g21480), .I1 (g9795), .I2 (g20444));
AN2X1 gate17635(.O (g21481), .I1 (g9711), .I2 (g20445));
AN2X1 gate17636(.O (g21482), .I1 (g15210), .I2 (g20446));
AN2X1 gate17637(.O (g21486), .I1 (g6832), .I2 (g20449));
AN2X1 gate17638(.O (g21487), .I1 (g9941), .I2 (g20450));
AN2X1 gate17639(.O (g21488), .I1 (g9857), .I2 (g20451));
AN2X1 gate17640(.O (g21489), .I1 (g15366), .I2 (g20452));
AN2X1 gate17641(.O (g21490), .I1 (g15296), .I2 (g20453));
AN2X1 gate17642(.O (g21494), .I1 (g6632), .I2 (g19792));
AN2X1 gate17643(.O (g21497), .I1 (g3006), .I2 (g20456));
AN2X1 gate17644(.O (g21517), .I1 (g9711), .I2 (g20461));
AN2X1 gate17645(.O (g21521), .I1 (g9941), .I2 (g20463));
AN2X1 gate17646(.O (g21522), .I1 (g9857), .I2 (g20464));
AN2X1 gate17647(.O (g21523), .I1 (g15296), .I2 (g20465));
AN2X1 gate17648(.O (g21527), .I1 (g7134), .I2 (g20468));
AN3X1 gate17649(.O (I28068), .I1 (g17802), .I2 (g18265), .I3 (g17882));
AN4X1 gate17650(.O (g21533), .I1 (g17724), .I2 (g18179), .I3 (g19799), .I4 (I28068));
AN2X1 gate17651(.O (g21553), .I1 (g9857), .I2 (g20476));
AN3X1 gate17652(.O (I28096), .I1 (g13907), .I2 (g14238), .I3 (g13946));
AN4X1 gate17653(.O (g21564), .I1 (g13886), .I2 (g14153), .I3 (g19799), .I4 (I28096));
AN3X1 gate17654(.O (I28103), .I1 (g17914), .I2 (g18358), .I3 (g17993));
AN4X1 gate17655(.O (g21569), .I1 (g17825), .I2 (g18286), .I3 (g19843), .I4 (I28103));
AN2X1 gate17656(.O (g21589), .I1 (g3002), .I2 (g19890));
AN3X1 gate17657(.O (g21593), .I1 (g16498), .I2 (g19484), .I3 (g14071));
AN3X1 gate17658(.O (I28126), .I1 (g13963), .I2 (g14360), .I3 (g14016));
AN4X1 gate17659(.O (g21597), .I1 (g13927), .I2 (g14268), .I3 (g19843), .I4 (I28126));
AN3X1 gate17660(.O (I28133), .I1 (g18025), .I2 (g18453), .I3 (g18110));
AN4X1 gate17661(.O (g21602), .I1 (g17937), .I2 (g18379), .I3 (g19876), .I4 (I28133));
AN2X1 gate17662(.O (g21610), .I1 (g7522), .I2 (g20490));
AN2X1 gate17663(.O (g21611), .I1 (g7471), .I2 (g19915));
AN3X1 gate17664(.O (g21622), .I1 (g16520), .I2 (g19505), .I3 (g14186));
AN3X1 gate17665(.O (I28155), .I1 (g14033), .I2 (g14472), .I3 (g14107));
AN4X1 gate17666(.O (g21626), .I1 (g13983), .I2 (g14390), .I3 (g19876), .I4 (I28155));
AN3X1 gate17667(.O (I28162), .I1 (g18142), .I2 (g18526), .I3 (g18226));
AN4X1 gate17668(.O (g21631), .I1 (g18048), .I2 (g18474), .I3 (g19907), .I4 (I28162));
AN2X1 gate17669(.O (g21635), .I1 (g7549), .I2 (g20496));
AN2X1 gate17670(.O (g21639), .I1 (g3398), .I2 (g20500));
AN3X1 gate17671(.O (g21650), .I1 (g16551), .I2 (g19524), .I3 (g14301));
AN3X1 gate17672(.O (I28181), .I1 (g14124), .I2 (g14559), .I3 (g14222));
AN4X1 gate17673(.O (g21654), .I1 (g14053), .I2 (g14502), .I3 (g19907), .I4 (I28181));
AN2X1 gate17674(.O (g21658), .I1 (g2896), .I2 (g20501));
AN2X1 gate17675(.O (g21666), .I1 (g3398), .I2 (g20504));
AN2X1 gate17676(.O (g21670), .I1 (g3554), .I2 (g20505));
AN3X1 gate17677(.O (g21681), .I1 (g16583), .I2 (g19534), .I3 (g14423));
AN2X1 gate17678(.O (g21687), .I1 (g3398), .I2 (g20516));
AN2X1 gate17679(.O (g21695), .I1 (g3554), .I2 (g20517));
AN2X1 gate17680(.O (g21699), .I1 (g3710), .I2 (g20518));
AN2X1 gate17681(.O (g21707), .I1 (g2892), .I2 (g19978));
AN2X1 gate17682(.O (g21723), .I1 (g3554), .I2 (g20534));
AN2X1 gate17683(.O (g21731), .I1 (g3710), .I2 (g20535));
AN2X1 gate17684(.O (g21735), .I1 (g3866), .I2 (g20536));
AN2X1 gate17685(.O (g21749), .I1 (g3710), .I2 (g20553));
AN2X1 gate17686(.O (g21757), .I1 (g3866), .I2 (g20554));
AN2X1 gate17687(.O (g21758), .I1 (g7607), .I2 (g20045));
AN2X1 gate17688(.O (g21773), .I1 (g3866), .I2 (g19078));
AN3X1 gate17689(.O (g21805), .I1 (g16679), .I2 (g19578), .I3 (g14776));
AN3X1 gate17690(.O (g21812), .I1 (g16705), .I2 (g19608), .I3 (g14811));
AN3X1 gate17691(.O (g21818), .I1 (g16736), .I2 (g19641), .I3 (g14863));
AN3X1 gate17692(.O (g21822), .I1 (g16778), .I2 (g19681), .I3 (g14936));
AN2X1 gate17693(.O (g21891), .I1 (g19302), .I2 (g11749));
AN2X1 gate17694(.O (g21892), .I1 (g19288), .I2 (g13011));
AN2X1 gate17695(.O (g21899), .I1 (g19323), .I2 (g11749));
AN2X1 gate17696(.O (g21900), .I1 (g19306), .I2 (g13011));
AN2X1 gate17697(.O (g21906), .I1 (g5715), .I2 (g20513));
AN2X1 gate17698(.O (g21911), .I1 (g19350), .I2 (g11749));
AN2X1 gate17699(.O (g21912), .I1 (g19327), .I2 (g13011));
AN2X1 gate17700(.O (g21913), .I1 (g4456), .I2 (g20519));
AN2X1 gate17701(.O (g21920), .I1 (g5773), .I2 (g20531));
AN2X1 gate17702(.O (g21925), .I1 (g19384), .I2 (g11749));
AN2X1 gate17703(.O (g21926), .I1 (g19354), .I2 (g13011));
AN2X1 gate17704(.O (g21931), .I1 (g4632), .I2 (g20539));
AN2X1 gate17705(.O (g21938), .I1 (g5832), .I2 (g20550));
AN2X1 gate17706(.O (g21990), .I1 (g291), .I2 (g21187));
AN2X1 gate17707(.O (g22004), .I1 (g978), .I2 (g21202));
AN2X1 gate17708(.O (g22015), .I1 (g1672), .I2 (g21217));
AN2X1 gate17709(.O (g22020), .I1 (g2366), .I2 (g21225));
AN3X1 gate17710(.O (I28582), .I1 (g19141), .I2 (g21133), .I3 (g21116));
AN4X1 gate17711(.O (g22036), .I1 (g21104), .I2 (g21095), .I3 (g21084), .I4 (I28582));
AN3X1 gate17712(.O (I28594), .I1 (g21167), .I2 (g21147), .I3 (g21134));
AN4X1 gate17713(.O (g22046), .I1 (g21117), .I2 (g21105), .I3 (g21096), .I4 (I28594));
AN3X1 gate17714(.O (I28609), .I1 (g21183), .I2 (g21168), .I3 (g21148));
AN4X1 gate17715(.O (g22062), .I1 (g21135), .I2 (g21118), .I3 (g21106), .I4 (I28609));
AN2X1 gate17716(.O (g22187), .I1 (g21564), .I2 (g20986));
AN2X1 gate17717(.O (g22196), .I1 (g21597), .I2 (g21012));
AN2X1 gate17718(.O (g22201), .I1 (g21271), .I2 (g16881));
AN2X1 gate17719(.O (g22202), .I1 (g21626), .I2 (g21036));
AN2X1 gate17720(.O (g22206), .I1 (g21895), .I2 (g11976));
AN2X1 gate17721(.O (g22207), .I1 (g21278), .I2 (g16910));
AN2X1 gate17722(.O (g22208), .I1 (g21654), .I2 (g21057));
AN2X1 gate17723(.O (g22211), .I1 (g21661), .I2 (g12027));
AN2X1 gate17724(.O (g22214), .I1 (g21907), .I2 (g12045));
AN2X1 gate17725(.O (g22215), .I1 (g21285), .I2 (g16940));
AN2X1 gate17726(.O (g22220), .I1 (g21690), .I2 (g12091));
AN2X1 gate17727(.O (g22223), .I1 (g21921), .I2 (g12109));
AN2X1 gate17728(.O (g22224), .I1 (g21293), .I2 (g16971));
AN2X1 gate17729(.O (g22228), .I1 (g21716), .I2 (g12136));
AN2X1 gate17730(.O (g22229), .I1 (g21661), .I2 (g12139));
AN2X1 gate17731(.O (g22235), .I1 (g21726), .I2 (g12163));
AN2X1 gate17732(.O (g22238), .I1 (g21939), .I2 (g12181));
AN2X1 gate17733(.O (g22244), .I1 (g21742), .I2 (g12198));
AN2X1 gate17734(.O (g22245), .I1 (g21690), .I2 (g12201));
AN2X1 gate17735(.O (g22250), .I1 (g21752), .I2 (g12225));
AN2X1 gate17736(.O (g22254), .I1 (g21716), .I2 (g12239));
AN2X1 gate17737(.O (g22255), .I1 (g21661), .I2 (g12242));
AN2X1 gate17738(.O (g22264), .I1 (g21766), .I2 (g12253));
AN2X1 gate17739(.O (g22265), .I1 (g21726), .I2 (g12256));
AN2X1 gate17740(.O (g22270), .I1 (g92), .I2 (g21529));
AN2X1 gate17741(.O (g22272), .I1 (g21742), .I2 (g12282));
AN2X1 gate17742(.O (g22273), .I1 (g21690), .I2 (g12285));
AN2X1 gate17743(.O (g22281), .I1 (g21782), .I2 (g12296));
AN2X1 gate17744(.O (g22282), .I1 (g21752), .I2 (g12299));
AN2X1 gate17745(.O (g22285), .I1 (g21716), .I2 (g12312));
AN2X1 gate17746(.O (g22289), .I1 (g780), .I2 (g21565));
AN2X1 gate17747(.O (g22291), .I1 (g21766), .I2 (g12318));
AN2X1 gate17748(.O (g22292), .I1 (g21726), .I2 (g12321));
AN2X1 gate17749(.O (g22305), .I1 (g21742), .I2 (g12340));
AN2X1 gate17750(.O (g22309), .I1 (g1466), .I2 (g21598));
AN2X1 gate17751(.O (g22311), .I1 (g21782), .I2 (g12346));
AN2X1 gate17752(.O (g22312), .I1 (g21752), .I2 (g12349));
AN2X1 gate17753(.O (g22333), .I1 (g21766), .I2 (g12370));
AN2X1 gate17754(.O (g22337), .I1 (g2160), .I2 (g21627));
AN2X1 gate17755(.O (g22340), .I1 (g88), .I2 (g21184));
AN2X1 gate17756(.O (g22358), .I1 (g21782), .I2 (g12389));
AN2X1 gate17757(.O (g22363), .I1 (g776), .I2 (g21199));
AN2X1 gate17758(.O (g22383), .I1 (g1462), .I2 (g21214));
AN2X1 gate17759(.O (g22398), .I1 (g2156), .I2 (g21222));
AN2X1 gate17760(.O (g22483), .I1 (g646), .I2 (g21861));
AN2X1 gate17761(.O (g22515), .I1 (g13873), .I2 (g21382));
AN2X1 gate17762(.O (g22516), .I1 (g20885), .I2 (g17442));
AN2X1 gate17763(.O (g22517), .I1 (g21895), .I2 (g12608));
AN2X1 gate17764(.O (g22526), .I1 (g1332), .I2 (g21867));
AN2X1 gate17765(.O (g22546), .I1 (g13886), .I2 (g21404));
AN2X1 gate17766(.O (g22555), .I1 (g13895), .I2 (g21415));
AN2X1 gate17767(.O (g22556), .I1 (g20904), .I2 (g17523));
AN2X1 gate17768(.O (g22557), .I1 (g21907), .I2 (g12654));
AN2X1 gate17769(.O (g22566), .I1 (g2026), .I2 (g21872));
AN2X1 gate17770(.O (g22577), .I1 (g13907), .I2 (g21429));
AN2X1 gate17771(.O (g22581), .I1 (g21895), .I2 (g12699));
AN2X1 gate17772(.O (g22587), .I1 (g13927), .I2 (g21441));
AN2X1 gate17773(.O (g22595), .I1 (g13936), .I2 (g21449));
AN2X1 gate17774(.O (g22596), .I1 (g20928), .I2 (g17613));
AN2X1 gate17775(.O (g22597), .I1 (g21921), .I2 (g12708));
AN2X1 gate17776(.O (g22606), .I1 (g2720), .I2 (g21876));
AN2X1 gate17777(.O (g22607), .I1 (g13946), .I2 (g21458));
AN2X1 gate17778(.O (g22610), .I1 (g660), .I2 (g21473));
AN2X1 gate17779(.O (g22614), .I1 (g13963), .I2 (g21477));
AN2X1 gate17780(.O (g22618), .I1 (g21907), .I2 (g12756));
AN2X1 gate17781(.O (g22624), .I1 (g13983), .I2 (g21483));
AN2X1 gate17782(.O (g22632), .I1 (g13992), .I2 (g21491));
AN2X1 gate17783(.O (g22633), .I1 (g20956), .I2 (g17710));
AN2X1 gate17784(.O (g22634), .I1 (g21939), .I2 (g12765));
AN2X1 gate17785(.O (g22637), .I1 (g20841), .I2 (g10927));
AN2X1 gate17786(.O (g22638), .I1 (g14001), .I2 (g21498));
AN2X1 gate17787(.O (g22643), .I1 (g14016), .I2 (g21505));
AN2X1 gate17788(.O (g22646), .I1 (g1346), .I2 (g21514));
AN2X1 gate17789(.O (g22650), .I1 (g14033), .I2 (g21518));
AN2X1 gate17790(.O (g22654), .I1 (g21921), .I2 (g12798));
AN2X1 gate17791(.O (g22660), .I1 (g14053), .I2 (g21524));
AN2X1 gate17792(.O (g22665), .I1 (g20920), .I2 (g6153));
AN2X1 gate17793(.O (g22666), .I1 (g21825), .I2 (g20014));
AN2X1 gate17794(.O (g22667), .I1 (g14062), .I2 (g21530));
AN2X1 gate17795(.O (g22674), .I1 (g14092), .I2 (g21537));
AN2X1 gate17796(.O (g22679), .I1 (g14107), .I2 (g21541));
AN2X1 gate17797(.O (g22682), .I1 (g2040), .I2 (g21550));
AN2X1 gate17798(.O (g22686), .I1 (g14124), .I2 (g21554));
AN2X1 gate17799(.O (g22690), .I1 (g21939), .I2 (g12837));
AN2X1 gate17800(.O (g22699), .I1 (g7338), .I2 (g21883));
AN2X1 gate17801(.O (g22700), .I1 (g7146), .I2 (g21558));
AN2X1 gate17802(.O (g22701), .I1 (g18174), .I2 (g21561));
AN2X1 gate17803(.O (g22707), .I1 (g14177), .I2 (g21566));
AN2X1 gate17804(.O (g22714), .I1 (g14207), .I2 (g21573));
AN2X1 gate17805(.O (g22719), .I1 (g14222), .I2 (g21577));
AN2X1 gate17806(.O (g22722), .I1 (g2734), .I2 (g21586));
AN2X1 gate17807(.O (g22726), .I1 (g3036), .I2 (g21886));
AN2X1 gate17808(.O (g22727), .I1 (g14238), .I2 (g21590));
AN2X1 gate17809(.O (g22732), .I1 (g18281), .I2 (g21594));
AN2X1 gate17810(.O (g22738), .I1 (g14292), .I2 (g21599));
AN2X1 gate17811(.O (g22745), .I1 (g14322), .I2 (g21606));
AN2X1 gate17812(.O (g22754), .I1 (g14342), .I2 (g21612));
AN2X1 gate17813(.O (g22759), .I1 (g14360), .I2 (g21619));
AN2X1 gate17814(.O (g22764), .I1 (g18374), .I2 (g21623));
AN2X1 gate17815(.O (g22770), .I1 (g14414), .I2 (g21628));
AN2X1 gate17816(.O (g22788), .I1 (g14454), .I2 (g21640));
AN2X1 gate17817(.O (g22793), .I1 (g14472), .I2 (g21647));
AN2X1 gate17818(.O (g22798), .I1 (g18469), .I2 (g21651));
AN2X1 gate17819(.O (g22804), .I1 (g2920), .I2 (g21655));
AN2X1 gate17820(.O (g22830), .I1 (g14541), .I2 (g21671));
AN2X1 gate17821(.O (g22835), .I1 (g14559), .I2 (g21678));
AN2X1 gate17822(.O (g22841), .I1 (g7583), .I2 (g21902));
AN2X1 gate17823(.O (g22842), .I1 (g3032), .I2 (g21682));
AN2X1 gate17824(.O (g22869), .I1 (g14596), .I2 (g21700));
AN2X1 gate17825(.O (g22874), .I1 (g7587), .I2 (g21708));
AN2X1 gate17826(.O (g22906), .I1 (g2924), .I2 (g21927));
AN2X1 gate17827(.O (g22984), .I1 (g16840), .I2 (g21400));
AN2X1 gate17828(.O (g23104), .I1 (g20842), .I2 (g15859));
AN2X1 gate17829(.O (g23106), .I1 (g5857), .I2 (g21050));
AN2X1 gate17830(.O (g23118), .I1 (g20850), .I2 (g15890));
AN2X1 gate17831(.O (g23119), .I1 (g5904), .I2 (g21069));
AN2X1 gate17832(.O (g23127), .I1 (g20858), .I2 (g15923));
AN2X1 gate17833(.O (g23128), .I1 (g5943), .I2 (g21079));
AN2X1 gate17834(.O (g23138), .I1 (g20866), .I2 (g15952));
AN2X1 gate17835(.O (g23139), .I1 (g5977), .I2 (g21093));
AN2X1 gate17836(.O (g23409), .I1 (g21533), .I2 (g22408));
AN2X1 gate17837(.O (g23414), .I1 (g21569), .I2 (g22421));
AN2X1 gate17838(.O (g23419), .I1 (g22755), .I2 (g19577));
AN2X1 gate17839(.O (g23423), .I1 (g21602), .I2 (g22443));
AN2X1 gate17840(.O (g23428), .I1 (g22789), .I2 (g19607));
AN2X1 gate17841(.O (g23432), .I1 (g21631), .I2 (g22476));
AN2X1 gate17842(.O (g23434), .I1 (g22831), .I2 (g19640));
AN2X1 gate17843(.O (g23440), .I1 (g22870), .I2 (g19680));
AN2X1 gate17844(.O (g23451), .I1 (g18552), .I2 (g22547));
AN2X1 gate17845(.O (g23458), .I1 (g18602), .I2 (g22588));
AN2X1 gate17846(.O (g23462), .I1 (g17988), .I2 (g22609));
AN2X1 gate17847(.O (g23467), .I1 (g18634), .I2 (g22625));
AN2X1 gate17848(.O (g23471), .I1 (g18105), .I2 (g22645));
AN2X1 gate17849(.O (g23476), .I1 (g18643), .I2 (g22661));
AN2X1 gate17850(.O (g23483), .I1 (g22945), .I2 (g8847));
AN2X1 gate17851(.O (g23484), .I1 (g18221), .I2 (g22681));
AN2X1 gate17852(.O (g23494), .I1 (g18328), .I2 (g22721));
AN2X1 gate17853(.O (g23496), .I1 (g5802), .I2 (g22300));
AN2X1 gate17854(.O (g23510), .I1 (g5890), .I2 (g22753));
AN2X1 gate17855(.O (g23512), .I1 (g5858), .I2 (g22328));
AN2X1 gate17856(.O (g23525), .I1 (g5929), .I2 (g22787));
AN2X1 gate17857(.O (g23527), .I1 (g5905), .I2 (g22353));
AN2X1 gate17858(.O (g23536), .I1 (g5963), .I2 (g22829));
AN2X1 gate17859(.O (g23538), .I1 (g5944), .I2 (g22376));
AN2X1 gate17860(.O (g23544), .I1 (g5992), .I2 (g22868));
AN2X1 gate17861(.O (g23547), .I1 (g8062), .I2 (g22405));
AN2X1 gate17862(.O (g23550), .I1 (g8132), .I2 (g22409));
AN2X1 gate17863(.O (g23551), .I1 (g8135), .I2 (g22412));
AN2X1 gate17864(.O (g23552), .I1 (g6136), .I2 (g22415));
AN2X1 gate17865(.O (g23554), .I1 (g8147), .I2 (g22418));
AN2X1 gate17866(.O (g23558), .I1 (g8200), .I2 (g22422));
AN2X1 gate17867(.O (g23559), .I1 (g8203), .I2 (g22425));
AN2X1 gate17868(.O (g23560), .I1 (g8206), .I2 (g22428));
AN2X1 gate17869(.O (g23563), .I1 (g8218), .I2 (g22431));
AN2X1 gate17870(.O (g23564), .I1 (g8221), .I2 (g22434));
AN2X1 gate17871(.O (g23565), .I1 (g6146), .I2 (g22437));
AN2X1 gate17872(.O (g23567), .I1 (g8233), .I2 (g22440));
AN2X1 gate17873(.O (g23571), .I1 (g3931), .I2 (g22445));
AN2X1 gate17874(.O (g23572), .I1 (g3934), .I2 (g22448));
AN2X1 gate17875(.O (g23573), .I1 (g3937), .I2 (g22451));
AN2X1 gate17876(.O (g23577), .I1 (g3957), .I2 (g22455));
AN2X1 gate17877(.O (g23578), .I1 (g3960), .I2 (g22458));
AN2X1 gate17878(.O (g23579), .I1 (g3963), .I2 (g22461));
AN2X1 gate17879(.O (g23582), .I1 (g3975), .I2 (g22464));
AN2X1 gate17880(.O (g23583), .I1 (g3978), .I2 (g22467));
AN2X1 gate17881(.O (g23584), .I1 (g6167), .I2 (g22470));
AN2X1 gate17882(.O (g23586), .I1 (g3990), .I2 (g22473));
AN2X1 gate17883(.O (g23590), .I1 (g4009), .I2 (g22477));
AN2X1 gate17884(.O (g23591), .I1 (g4012), .I2 (g22480));
AN2X1 gate17885(.O (g23592), .I1 (g17640), .I2 (g22986));
AN2X1 gate17886(.O (g23593), .I1 (g22845), .I2 (g20365));
AN2X1 gate17887(.O (g23598), .I1 (g4038), .I2 (g22484));
AN2X1 gate17888(.O (g23599), .I1 (g4041), .I2 (g22487));
AN2X1 gate17889(.O (g23600), .I1 (g4044), .I2 (g22490));
AN2X1 gate17890(.O (g23604), .I1 (g4064), .I2 (g22494));
AN2X1 gate17891(.O (g23605), .I1 (g4067), .I2 (g22497));
AN2X1 gate17892(.O (g23606), .I1 (g4070), .I2 (g22500));
AN2X1 gate17893(.O (g23609), .I1 (g4082), .I2 (g22503));
AN2X1 gate17894(.O (g23610), .I1 (g4085), .I2 (g22506));
AN2X1 gate17895(.O (g23611), .I1 (g6194), .I2 (g22509));
AN2X1 gate17896(.O (g23615), .I1 (g4107), .I2 (g22512));
AN2X1 gate17897(.O (g23616), .I1 (g17724), .I2 (g22988));
AN2X1 gate17898(.O (g23617), .I1 (g22810), .I2 (g20382));
AN2X1 gate17899(.O (g23618), .I1 (g22608), .I2 (g20383));
AN2X1 gate17900(.O (g23622), .I1 (g4136), .I2 (g22520));
AN2X1 gate17901(.O (g23623), .I1 (g4139), .I2 (g22523));
AN2X1 gate17902(.O (g23624), .I1 (g17741), .I2 (g22989));
AN2X1 gate17903(.O (g23625), .I1 (g22880), .I2 (g20388));
AN2X1 gate17904(.O (g23630), .I1 (g4165), .I2 (g22527));
AN2X1 gate17905(.O (g23631), .I1 (g4168), .I2 (g22530));
AN2X1 gate17906(.O (g23632), .I1 (g4171), .I2 (g22533));
AN2X1 gate17907(.O (g23636), .I1 (g4191), .I2 (g22537));
AN2X1 gate17908(.O (g23637), .I1 (g4194), .I2 (g22540));
AN2X1 gate17909(.O (g23638), .I1 (g4197), .I2 (g22543));
AN2X1 gate17910(.O (g23639), .I1 (g21825), .I2 (g22805));
AN2X1 gate17911(.O (g23643), .I1 (g17802), .I2 (g22991));
AN2X1 gate17912(.O (g23659), .I1 (g22784), .I2 (g17500));
AN2X1 gate17913(.O (g23664), .I1 (g4246), .I2 (g22552));
AN2X1 gate17914(.O (g23665), .I1 (g17825), .I2 (g22995));
AN2X1 gate17915(.O (g23666), .I1 (g22851), .I2 (g20407));
AN2X1 gate17916(.O (g23667), .I1 (g22644), .I2 (g20408));
AN2X1 gate17917(.O (g23671), .I1 (g4275), .I2 (g22560));
AN2X1 gate17918(.O (g23672), .I1 (g4278), .I2 (g22563));
AN2X1 gate17919(.O (g23673), .I1 (g17842), .I2 (g22996));
AN2X1 gate17920(.O (g23674), .I1 (g22915), .I2 (g20413));
AN2X1 gate17921(.O (g23679), .I1 (g4304), .I2 (g22567));
AN2X1 gate17922(.O (g23680), .I1 (g4307), .I2 (g22570));
AN2X1 gate17923(.O (g23681), .I1 (g4310), .I2 (g22573));
AN2X1 gate17924(.O (g23686), .I1 (g17882), .I2 (g22998));
AN2X1 gate17925(.O (g23687), .I1 (g22668), .I2 (g17570));
AN2X1 gate17926(.O (g23689), .I1 (g6513), .I2 (g23001));
AN2X1 gate17927(.O (g23693), .I1 (g17914), .I2 (g23002));
AN2X1 gate17928(.O (g23709), .I1 (g22826), .I2 (g17591));
AN2X1 gate17929(.O (g23714), .I1 (g4401), .I2 (g22592));
AN2X1 gate17930(.O (g23715), .I1 (g17937), .I2 (g23006));
AN2X1 gate17931(.O (g23716), .I1 (g22886), .I2 (g20432));
AN2X1 gate17932(.O (g23717), .I1 (g22680), .I2 (g20433));
AN2X1 gate17933(.O (g23721), .I1 (g4430), .I2 (g22600));
AN2X1 gate17934(.O (g23722), .I1 (g4433), .I2 (g22603));
AN2X1 gate17935(.O (g23723), .I1 (g17954), .I2 (g23007));
AN2X1 gate17936(.O (g23724), .I1 (g22940), .I2 (g20438));
AN2X1 gate17937(.O (g23726), .I1 (g21825), .I2 (g22843));
AN2X1 gate17938(.O (g23734), .I1 (g17974), .I2 (g23008));
AN2X1 gate17939(.O (g23735), .I1 (g22949), .I2 (g9450));
AN2X1 gate17940(.O (g23740), .I1 (g17993), .I2 (g23012));
AN2X1 gate17941(.O (g23741), .I1 (g22708), .I2 (g17667));
AN2X1 gate17942(.O (g23743), .I1 (g6777), .I2 (g23015));
AN2X1 gate17943(.O (g23747), .I1 (g18025), .I2 (g23016));
AN2X1 gate17944(.O (g23763), .I1 (g22865), .I2 (g17688));
AN2X1 gate17945(.O (g23768), .I1 (g4570), .I2 (g22629));
AN2X1 gate17946(.O (g23769), .I1 (g18048), .I2 (g23020));
AN2X1 gate17947(.O (g23770), .I1 (g22921), .I2 (g20454));
AN2X1 gate17948(.O (g23771), .I1 (g22720), .I2 (g20455));
AN2X1 gate17949(.O (g23772), .I1 (g21825), .I2 (g22875));
AN2X1 gate17950(.O (g23776), .I1 (g18074), .I2 (g23021));
AN2X1 gate17951(.O (g23777), .I1 (g22949), .I2 (g9528));
AN2X1 gate17952(.O (g23778), .I1 (g22954), .I2 (g9531));
AN2X1 gate17953(.O (g23789), .I1 (g18091), .I2 (g23024));
AN2X1 gate17954(.O (g23790), .I1 (g22958), .I2 (g9592));
AN2X1 gate17955(.O (g23795), .I1 (g18110), .I2 (g23028));
AN2X1 gate17956(.O (g23796), .I1 (g22739), .I2 (g17767));
AN2X1 gate17957(.O (g23798), .I1 (g7079), .I2 (g23031));
AN2X1 gate17958(.O (g23802), .I1 (g18142), .I2 (g23032));
AN2X1 gate17959(.O (g23818), .I1 (g22900), .I2 (g17788));
AN2X1 gate17960(.O (g23820), .I1 (g3013), .I2 (g23036));
AN2X1 gate17961(.O (g23822), .I1 (g14148), .I2 (g23037));
AN2X1 gate17962(.O (g23824), .I1 (g22949), .I2 (g9641));
AN2X1 gate17963(.O (g23825), .I1 (g22954), .I2 (g9644));
AN2X1 gate17964(.O (g23829), .I1 (g18190), .I2 (g23038));
AN2X1 gate17965(.O (g23830), .I1 (g22958), .I2 (g9670));
AN2X1 gate17966(.O (g23831), .I1 (g22962), .I2 (g9673));
AN2X1 gate17967(.O (g23842), .I1 (g18207), .I2 (g23041));
AN2X1 gate17968(.O (g23843), .I1 (g22966), .I2 (g9734));
AN2X1 gate17969(.O (g23848), .I1 (g18226), .I2 (g23045));
AN2X1 gate17970(.O (g23849), .I1 (g22771), .I2 (g17868));
AN2X1 gate17971(.O (g23851), .I1 (g7329), .I2 (g23048));
AN2X1 gate17972(.O (g23852), .I1 (g19179), .I2 (g22696));
AN2X1 gate17973(.O (g23854), .I1 (g18265), .I2 (g23049));
AN2X1 gate17974(.O (g23855), .I1 (g22954), .I2 (g9767));
AN2X1 gate17975(.O (g23857), .I1 (g14263), .I2 (g23056));
AN2X1 gate17976(.O (g23859), .I1 (g22958), .I2 (g9787));
AN2X1 gate17977(.O (g23860), .I1 (g22962), .I2 (g9790));
AN2X1 gate17978(.O (g23864), .I1 (g18297), .I2 (g23057));
AN2X1 gate17979(.O (g23865), .I1 (g22966), .I2 (g9816));
AN2X1 gate17980(.O (g23866), .I1 (g22971), .I2 (g9819));
AN2X1 gate17981(.O (g23877), .I1 (g18314), .I2 (g23060));
AN2X1 gate17982(.O (g23878), .I1 (g22975), .I2 (g9880));
AN2X1 gate17983(.O (g23886), .I1 (g18341), .I2 (g23064));
AN2X1 gate17984(.O (g23888), .I1 (g18358), .I2 (g23069));
AN2X1 gate17985(.O (g23889), .I1 (g22962), .I2 (g9913));
AN2X1 gate17986(.O (g23891), .I1 (g14385), .I2 (g23074));
AN2X1 gate17987(.O (g23893), .I1 (g22966), .I2 (g9933));
AN2X1 gate17988(.O (g23894), .I1 (g22971), .I2 (g9936));
AN2X1 gate17989(.O (g23898), .I1 (g18390), .I2 (g23075));
AN2X1 gate17990(.O (g23899), .I1 (g22975), .I2 (g9962));
AN2X1 gate17991(.O (g23900), .I1 (g22980), .I2 (g9965));
AN2X1 gate17992(.O (g23904), .I1 (g3010), .I2 (g22750));
AN2X1 gate17993(.O (g23907), .I1 (g18436), .I2 (g23079));
AN2X1 gate17994(.O (g23909), .I1 (g18453), .I2 (g23082));
AN2X1 gate17995(.O (g23910), .I1 (g22971), .I2 (g10067));
AN2X1 gate17996(.O (g23912), .I1 (g14497), .I2 (g23087));
AN2X1 gate17997(.O (g23914), .I1 (g22975), .I2 (g10087));
AN2X1 gate17998(.O (g23915), .I1 (g22980), .I2 (g10090));
AN2X1 gate17999(.O (g23917), .I1 (g7545), .I2 (g23088));
AN2X1 gate18000(.O (g23939), .I1 (g18509), .I2 (g23095));
AN2X1 gate18001(.O (g23941), .I1 (g18526), .I2 (g23098));
AN2X1 gate18002(.O (g23942), .I1 (g22980), .I2 (g10176));
AN2X1 gate18003(.O (g23944), .I1 (g7570), .I2 (g23103));
AN2X1 gate18004(.O (g23971), .I1 (g18573), .I2 (g23112));
AN2X1 gate18005(.O (g23972), .I1 (g2903), .I2 (g23115));
AN2X1 gate18006(.O (g24029), .I1 (g2900), .I2 (g22903));
AN2X1 gate18007(.O (g24211), .I1 (g22014), .I2 (g10969));
AN2X1 gate18008(.O (g24217), .I1 (g22825), .I2 (g10999));
AN2X1 gate18009(.O (g24221), .I1 (g22979), .I2 (g11042));
AN2X1 gate18010(.O (g24224), .I1 (g22219), .I2 (g11045));
AN2X1 gate18011(.O (g24229), .I1 (g22232), .I2 (g11105));
AN2X1 gate18012(.O (g24236), .I1 (g22243), .I2 (g11157));
AN2X1 gate18013(.O (g24241), .I1 (g22259), .I2 (g11228));
AN2X1 gate18014(.O (g24246), .I1 (g21982), .I2 (g11291));
AN2X1 gate18015(.O (g24247), .I1 (g22551), .I2 (g11297));
AN2X1 gate18016(.O (g24253), .I1 (g21995), .I2 (g11370));
AN2X1 gate18017(.O (g24256), .I1 (g22003), .I2 (g11438));
AN3X1 gate18018(.O (g24427), .I1 (g17086), .I2 (g24134), .I3 (g13626));
AN2X1 gate18019(.O (g24429), .I1 (g24115), .I2 (g13614));
AN3X1 gate18020(.O (g24431), .I1 (g17124), .I2 (g24153), .I3 (g13637));
AN3X1 gate18021(.O (g24432), .I1 (g14642), .I2 (g15904), .I3 (g24115));
AN2X1 gate18022(.O (g24433), .I1 (g24134), .I2 (g13626));
AN3X1 gate18023(.O (g24435), .I1 (g17151), .I2 (g24168), .I3 (g13649));
AN3X1 gate18024(.O (g24436), .I1 (g14669), .I2 (g15933), .I3 (g24134));
AN2X1 gate18025(.O (g24437), .I1 (g24153), .I2 (g13637));
AN3X1 gate18026(.O (g24439), .I1 (g14703), .I2 (g15962), .I3 (g24153));
AN2X1 gate18027(.O (g24440), .I1 (g24168), .I2 (g13649));
AN3X1 gate18028(.O (g24441), .I1 (g14737), .I2 (g15981), .I3 (g24168));
AN3X1 gate18029(.O (g24478), .I1 (g23545), .I2 (g21119), .I3 (g21227));
AN3X1 gate18030(.O (g24529), .I1 (g19933), .I2 (g17896), .I3 (g23403));
AN3X1 gate18031(.O (g24540), .I1 (g18548), .I2 (g23089), .I3 (g23403));
AN3X1 gate18032(.O (g24541), .I1 (g23420), .I2 (g17896), .I3 (g23052));
AN3X1 gate18033(.O (g24542), .I1 (g19950), .I2 (g18007), .I3 (g23410));
AN3X1 gate18034(.O (g24550), .I1 (g18548), .I2 (g23420), .I3 (g19948));
AN3X1 gate18035(.O (g24552), .I1 (g18598), .I2 (g23107), .I3 (g23410));
AN3X1 gate18036(.O (g24553), .I1 (g23429), .I2 (g18007), .I3 (g23071));
AN3X1 gate18037(.O (g24554), .I1 (g19977), .I2 (g18124), .I3 (g23415));
AN2X1 gate18038(.O (g24559), .I1 (g79), .I2 (g23448));
AN3X1 gate18039(.O (g24561), .I1 (g18598), .I2 (g23429), .I3 (g19975));
AN3X1 gate18040(.O (g24563), .I1 (g18630), .I2 (g23120), .I3 (g23415));
AN3X1 gate18041(.O (g24564), .I1 (g23435), .I2 (g18124), .I3 (g23084));
AN3X1 gate18042(.O (g24565), .I1 (g20007), .I2 (g18240), .I3 (g23424));
AN2X1 gate18043(.O (g24569), .I1 (g767), .I2 (g23455));
AN3X1 gate18044(.O (g24571), .I1 (g18630), .I2 (g23435), .I3 (g20005));
AN3X1 gate18045(.O (g24573), .I1 (g18639), .I2 (g23129), .I3 (g23424));
AN3X1 gate18046(.O (g24574), .I1 (g23441), .I2 (g18240), .I3 (g23100));
AN2X1 gate18047(.O (g24578), .I1 (g1453), .I2 (g23464));
AN3X1 gate18048(.O (g24580), .I1 (g18639), .I2 (g23441), .I3 (g20043));
AN2X1 gate18049(.O (g24585), .I1 (g2147), .I2 (g23473));
AN2X1 gate18050(.O (g24590), .I1 (g23486), .I2 (g23478));
AN2X1 gate18051(.O (g24591), .I1 (g83), .I2 (g23853));
AN2X1 gate18052(.O (g24595), .I1 (g23502), .I2 (g23489));
AN2X1 gate18053(.O (g24596), .I1 (g771), .I2 (g23887));
AN2X1 gate18054(.O (g24603), .I1 (g23518), .I2 (g23505));
AN2X1 gate18055(.O (g24604), .I1 (g1457), .I2 (g23908));
AN2X1 gate18056(.O (g24610), .I1 (g23533), .I2 (g23521));
AN2X1 gate18057(.O (g24611), .I1 (g2151), .I2 (g23940));
AN2X1 gate18058(.O (g24644), .I1 (g17203), .I2 (g24115));
AN2X1 gate18059(.O (g24664), .I1 (g17208), .I2 (g24134));
AN2X1 gate18060(.O (g24676), .I1 (g13568), .I2 (g24115));
AN2X1 gate18061(.O (g24683), .I1 (g17214), .I2 (g24153));
AN2X1 gate18062(.O (g24695), .I1 (g13576), .I2 (g24134));
AN2X1 gate18063(.O (g24700), .I1 (g17217), .I2 (g24168));
AN2X1 gate18064(.O (g24712), .I1 (g13585), .I2 (g24153));
AN2X1 gate18065(.O (g24723), .I1 (g13605), .I2 (g24168));
AN2X1 gate18066(.O (g24745), .I1 (g15454), .I2 (g24096));
AN2X1 gate18067(.O (g24746), .I1 (g15454), .I2 (g24098));
AN2X1 gate18068(.O (g24747), .I1 (g9427), .I2 (g24099));
AN2X1 gate18069(.O (g24748), .I1 (g672), .I2 (g24101));
AN2X1 gate18070(.O (g24749), .I1 (g15540), .I2 (g24102));
AN2X1 gate18071(.O (g24750), .I1 (g15454), .I2 (g24104));
AN2X1 gate18072(.O (g24751), .I1 (g9427), .I2 (g24105));
AN2X1 gate18073(.O (g24752), .I1 (g9507), .I2 (g24106));
AN2X1 gate18074(.O (g24754), .I1 (g15540), .I2 (g24107));
AN2X1 gate18075(.O (g24755), .I1 (g9569), .I2 (g24108));
AN2X1 gate18076(.O (g24757), .I1 (g1358), .I2 (g24110));
AN2X1 gate18077(.O (g24758), .I1 (g15618), .I2 (g24111));
AN2X1 gate18078(.O (g24759), .I1 (g21825), .I2 (g23885));
AN2X1 gate18079(.O (g24760), .I1 (g9427), .I2 (g24112));
AN2X1 gate18080(.O (g24761), .I1 (g9507), .I2 (g24113));
AN2X1 gate18081(.O (g24762), .I1 (g12876), .I2 (g24114));
AN2X1 gate18082(.O (g24767), .I1 (g15540), .I2 (g24121));
AN2X1 gate18083(.O (g24768), .I1 (g9569), .I2 (g24122));
AN2X1 gate18084(.O (g24769), .I1 (g9649), .I2 (g24123));
AN2X1 gate18085(.O (g24772), .I1 (g15618), .I2 (g24124));
AN2X1 gate18086(.O (g24773), .I1 (g9711), .I2 (g24125));
AN2X1 gate18087(.O (g24774), .I1 (g2052), .I2 (g24127));
AN2X1 gate18088(.O (g24775), .I1 (g15694), .I2 (g24128));
AN2X1 gate18089(.O (g24776), .I1 (g9507), .I2 (g24129));
AN2X1 gate18090(.O (g24777), .I1 (g12876), .I2 (g24130));
AN2X1 gate18091(.O (g24779), .I1 (g9569), .I2 (g24131));
AN2X1 gate18092(.O (g24780), .I1 (g9649), .I2 (g24132));
AN2X1 gate18093(.O (g24781), .I1 (g12916), .I2 (g24133));
AN2X1 gate18094(.O (g24788), .I1 (g15618), .I2 (g24140));
AN2X1 gate18095(.O (g24789), .I1 (g9711), .I2 (g24141));
AN2X1 gate18096(.O (g24790), .I1 (g9795), .I2 (g24142));
AN2X1 gate18097(.O (g24792), .I1 (g15694), .I2 (g24143));
AN2X1 gate18098(.O (g24793), .I1 (g9857), .I2 (g24144));
AN2X1 gate18099(.O (g24794), .I1 (g2746), .I2 (g24146));
AN2X1 gate18100(.O (g24795), .I1 (g12017), .I2 (g24232));
AN2X1 gate18101(.O (g24796), .I1 (g12876), .I2 (g24147));
AN2X1 gate18102(.O (g24798), .I1 (g9649), .I2 (g24148));
AN2X1 gate18103(.O (g24799), .I1 (g12916), .I2 (g24149));
AN2X1 gate18104(.O (g24802), .I1 (g9711), .I2 (g24150));
AN2X1 gate18105(.O (g24803), .I1 (g9795), .I2 (g24151));
AN2X1 gate18106(.O (g24804), .I1 (g12945), .I2 (g24152));
AN2X1 gate18107(.O (g24809), .I1 (g15694), .I2 (g24159));
AN2X1 gate18108(.O (g24810), .I1 (g9857), .I2 (g24160));
AN2X1 gate18109(.O (g24811), .I1 (g9941), .I2 (g24161));
AN2X1 gate18110(.O (g24813), .I1 (g21825), .I2 (g23905));
AN2X1 gate18111(.O (g24818), .I1 (g12916), .I2 (g24162));
AN2X1 gate18112(.O (g24821), .I1 (g9795), .I2 (g24163));
AN2X1 gate18113(.O (g24822), .I1 (g12945), .I2 (g24164));
AN2X1 gate18114(.O (g24824), .I1 (g9857), .I2 (g24165));
AN2X1 gate18115(.O (g24825), .I1 (g9941), .I2 (g24166));
AN2X1 gate18116(.O (g24826), .I1 (g12974), .I2 (g24167));
AN2X1 gate18117(.O (g24831), .I1 (g24100), .I2 (g20401));
AN2X1 gate18118(.O (g24838), .I1 (g12945), .I2 (g24175));
AN2X1 gate18119(.O (g24840), .I1 (g9941), .I2 (g24176));
AN2X1 gate18120(.O (g24841), .I1 (g12974), .I2 (g24177));
AN2X1 gate18121(.O (g24843), .I1 (g21825), .I2 (g23918));
AN2X1 gate18122(.O (g24846), .I1 (g24109), .I2 (g20426));
AN2X1 gate18123(.O (g24853), .I1 (g12974), .I2 (g24180));
AN2X1 gate18124(.O (g24855), .I1 (g18174), .I2 (g23731));
AN2X1 gate18125(.O (g24858), .I1 (g24047), .I2 (g18873));
AN2X1 gate18126(.O (g24861), .I1 (g24126), .I2 (g20448));
AN2X1 gate18127(.O (g24867), .I1 (g666), .I2 (g23779));
AN2X1 gate18128(.O (g24869), .I1 (g24047), .I2 (g18894));
AN2X1 gate18129(.O (g24870), .I1 (g18281), .I2 (g23786));
AN2X1 gate18130(.O (g24874), .I1 (g24060), .I2 (g18899));
AN2X1 gate18131(.O (g24876), .I1 (g24145), .I2 (g20467));
AN2X1 gate18132(.O (g24878), .I1 (g19830), .I2 (g24210));
AN2X1 gate18133(.O (g24881), .I1 (g24047), .I2 (g18912));
AN2X1 gate18134(.O (g24882), .I1 (g1352), .I2 (g23832));
AN2X1 gate18135(.O (g24884), .I1 (g24060), .I2 (g18917));
AN2X1 gate18136(.O (g24885), .I1 (g18374), .I2 (g23839));
AN2X1 gate18137(.O (g24888), .I1 (g24073), .I2 (g18922));
AN2X1 gate18138(.O (g24898), .I1 (g24060), .I2 (g18931));
AN2X1 gate18139(.O (g24899), .I1 (g2046), .I2 (g23867));
AN2X1 gate18140(.O (g24901), .I1 (g24073), .I2 (g18936));
AN2X1 gate18141(.O (g24902), .I1 (g18469), .I2 (g23874));
AN2X1 gate18142(.O (g24905), .I1 (g24084), .I2 (g18941));
AN2X1 gate18143(.O (g24906), .I1 (g18886), .I2 (g23879));
AN2X1 gate18144(.O (g24907), .I1 (g7466), .I2 (g24220));
AN2X1 gate18145(.O (g24908), .I1 (g7342), .I2 (g23882));
AN2X1 gate18146(.O (g24921), .I1 (g24073), .I2 (g18951));
AN2X1 gate18147(.O (g24922), .I1 (g2740), .I2 (g23901));
AN2X1 gate18148(.O (g24924), .I1 (g24084), .I2 (g18956));
AN2X1 gate18149(.O (g24938), .I1 (g24084), .I2 (g18967));
AN2X1 gate18150(.O (g24964), .I1 (g7595), .I2 (g24251));
AN2X1 gate18151(.O (g24974), .I1 (g7600), .I2 (g24030));
AN2X1 gate18152(.O (g25086), .I1 (g23444), .I2 (g10880));
AN2X1 gate18153(.O (g25102), .I1 (g23444), .I2 (g10915));
AN2X1 gate18154(.O (g25117), .I1 (g23444), .I2 (g10974));
AN3X1 gate18155(.O (g25128), .I1 (g17051), .I2 (g24115), .I3 (g13614));
AN2X1 gate18156(.O (g25178), .I1 (g24623), .I2 (g20634));
AN2X1 gate18157(.O (g25181), .I1 (g24636), .I2 (g20673));
AN2X1 gate18158(.O (g25182), .I1 (g24681), .I2 (g20676));
AN2X1 gate18159(.O (g25184), .I1 (g24694), .I2 (g20735));
AN2X1 gate18160(.O (g25187), .I1 (g24633), .I2 (g16608));
AN2X1 gate18161(.O (g25188), .I1 (g24652), .I2 (g20763));
AN2X1 gate18162(.O (g25192), .I1 (g24711), .I2 (g20790));
AN2X1 gate18163(.O (g25193), .I1 (g24653), .I2 (g16626));
AN2X1 gate18164(.O (g25196), .I1 (g24672), .I2 (g16640));
AN2X1 gate18165(.O (g25198), .I1 (g24691), .I2 (g16651));
AN2X1 gate18166(.O (g25269), .I1 (g24648), .I2 (g8700));
AN2X1 gate18167(.O (g25277), .I1 (g24648), .I2 (g8714));
AN2X1 gate18168(.O (g25278), .I1 (g24668), .I2 (g8719));
AN2X1 gate18169(.O (g25281), .I1 (g5606), .I2 (g24815));
AN2X1 gate18170(.O (g25282), .I1 (g24648), .I2 (g8748));
AN2X1 gate18171(.O (g25286), .I1 (g24668), .I2 (g8752));
AN2X1 gate18172(.O (g25287), .I1 (g24687), .I2 (g8757));
AN2X1 gate18173(.O (g25289), .I1 (g5631), .I2 (g24834));
AN2X1 gate18174(.O (g25290), .I1 (g24668), .I2 (g8771));
AN2X1 gate18175(.O (g25294), .I1 (g24687), .I2 (g8775));
AN2X1 gate18176(.O (g25295), .I1 (g24704), .I2 (g8780));
AN2X1 gate18177(.O (g25299), .I1 (g5659), .I2 (g24850));
AN2X1 gate18178(.O (g25300), .I1 (g24687), .I2 (g8794));
AN2X1 gate18179(.O (g25304), .I1 (g24704), .I2 (g8798));
AN2X1 gate18180(.O (g25309), .I1 (g5697), .I2 (g24864));
AN2X1 gate18181(.O (g25310), .I1 (g24704), .I2 (g8813));
AN3X1 gate18182(.O (g25318), .I1 (g24682), .I2 (g19358), .I3 (g19335));
AN2X1 gate18183(.O (g25321), .I1 (g25075), .I2 (g9669));
AN2X1 gate18184(.O (g25328), .I1 (g24644), .I2 (g17892));
AN2X1 gate18185(.O (g25334), .I1 (g24644), .I2 (g17984));
AN2X1 gate18186(.O (g25337), .I1 (g24664), .I2 (g18003));
AN2X1 gate18187(.O (g25342), .I1 (g5851), .I2 (g24600));
AN2X1 gate18188(.O (g25346), .I1 (g24644), .I2 (g18084));
AN2X1 gate18189(.O (g25348), .I1 (g24664), .I2 (g18101));
AN2X1 gate18190(.O (g25351), .I1 (g24683), .I2 (g18120));
AN2X1 gate18191(.O (g25356), .I1 (g5898), .I2 (g24607));
AN2X1 gate18192(.O (g25360), .I1 (g24664), .I2 (g18200));
AN2X1 gate18193(.O (g25362), .I1 (g24683), .I2 (g18217));
AN2X1 gate18194(.O (g25365), .I1 (g24700), .I2 (g18236));
AN2X1 gate18195(.O (g25371), .I1 (g5937), .I2 (g24619));
AN2X1 gate18196(.O (g25375), .I1 (g24683), .I2 (g18307));
AN2X1 gate18197(.O (g25377), .I1 (g24700), .I2 (g18324));
AN2X1 gate18198(.O (g25388), .I1 (g5971), .I2 (g24630));
AN2X1 gate18199(.O (g25392), .I1 (g24700), .I2 (g18400));
AN2X1 gate18200(.O (g25453), .I1 (g6142), .I2 (g24763));
AN2X1 gate18201(.O (g25457), .I1 (g6163), .I2 (g24784));
AN2X1 gate18202(.O (g25461), .I1 (g6190), .I2 (g24805));
AN2X1 gate18203(.O (g25466), .I1 (g6222), .I2 (g24827));
AN2X1 gate18204(.O (g25470), .I1 (g24479), .I2 (g20400));
AN2X1 gate18205(.O (g25475), .I1 (g14148), .I2 (g25087));
AN2X1 gate18206(.O (g25482), .I1 (g24480), .I2 (g17567));
AN2X1 gate18207(.O (g25483), .I1 (g24481), .I2 (g20421));
AN2X1 gate18208(.O (g25487), .I1 (g24485), .I2 (g20425));
AN2X1 gate18209(.O (g25505), .I1 (g6707), .I2 (g25094));
AN2X1 gate18210(.O (g25506), .I1 (g14263), .I2 (g25095));
AN2X1 gate18211(.O (g25513), .I1 (g24487), .I2 (g17664));
AN2X1 gate18212(.O (g25514), .I1 (g24488), .I2 (g20443));
AN2X1 gate18213(.O (g25518), .I1 (g24489), .I2 (g20447));
AN2X1 gate18214(.O (g25552), .I1 (g7009), .I2 (g25104));
AN2X1 gate18215(.O (g25553), .I1 (g14385), .I2 (g25105));
AN2X1 gate18216(.O (g25560), .I1 (g24494), .I2 (g17764));
AN2X1 gate18217(.O (g25561), .I1 (g24495), .I2 (g20462));
AN2X1 gate18218(.O (g25565), .I1 (g24496), .I2 (g20466));
AN2X1 gate18219(.O (g25618), .I1 (g7259), .I2 (g25110));
AN2X1 gate18220(.O (g25619), .I1 (g14497), .I2 (g25111));
AN2X1 gate18221(.O (g25626), .I1 (g24504), .I2 (g17865));
AN2X1 gate18222(.O (g25627), .I1 (g24505), .I2 (g20477));
AN2X1 gate18223(.O (g25628), .I1 (g21008), .I2 (g25115));
AN2X1 gate18224(.O (g25629), .I1 (g3024), .I2 (g25116));
AN2X1 gate18225(.O (g25697), .I1 (g7455), .I2 (g25120));
AN2X1 gate18226(.O (g25881), .I1 (g2908), .I2 (g25126));
AN2X1 gate18227(.O (g25951), .I1 (g24800), .I2 (g13670));
AN2X1 gate18228(.O (g25953), .I1 (g24783), .I2 (g13699));
AN2X1 gate18229(.O (g25957), .I1 (g24782), .I2 (g11869));
AN2X1 gate18230(.O (g25961), .I1 (g24770), .I2 (g11901));
AN2X1 gate18231(.O (g25963), .I1 (g24756), .I2 (g11944));
AN2X1 gate18232(.O (g25968), .I1 (g24871), .I2 (g11986));
AN2X1 gate18233(.O (g25972), .I1 (g24859), .I2 (g12042));
AN2X1 gate18234(.O (g25973), .I1 (g24847), .I2 (g13838));
AN2X1 gate18235(.O (g25975), .I1 (g24606), .I2 (g21917));
AN2X1 gate18236(.O (g25977), .I1 (g24845), .I2 (g12089));
AN2X1 gate18237(.O (g25978), .I1 (g24836), .I2 (g13850));
AN2X1 gate18238(.O (g25980), .I1 (g24663), .I2 (g21928));
AN2X1 gate18239(.O (g25981), .I1 (g24819), .I2 (g13858));
AN2X1 gate18240(.O (g26023), .I1 (g25422), .I2 (g24912));
AN2X1 gate18241(.O (g26024), .I1 (g25301), .I2 (g21102));
AN2X1 gate18242(.O (g26026), .I1 (g25431), .I2 (g24929));
AN2X1 gate18243(.O (g26027), .I1 (g25418), .I2 (g22271));
AN2X1 gate18244(.O (g26028), .I1 (g25438), .I2 (g24941));
AN2X1 gate18245(.O (g26029), .I1 (g25445), .I2 (g24952));
AN2X1 gate18246(.O (g26030), .I1 (g25429), .I2 (g22304));
AN2X1 gate18247(.O (g26032), .I1 (g25379), .I2 (g19415));
AN2X1 gate18248(.O (g26033), .I1 (g25395), .I2 (g19452));
AN2X1 gate18249(.O (g26034), .I1 (g25405), .I2 (g19479));
AN2X1 gate18250(.O (g26035), .I1 (g25523), .I2 (g19483));
AN2X1 gate18251(.O (g26036), .I1 (g25413), .I2 (g19502));
AN2X1 gate18252(.O (g26038), .I1 (g25589), .I2 (g19504));
AN2X1 gate18253(.O (g26039), .I1 (g25668), .I2 (g19523));
AN2X1 gate18254(.O (g26040), .I1 (g25745), .I2 (g19533));
AN2X1 gate18255(.O (g26051), .I1 (g70), .I2 (g25296));
AN2X1 gate18256(.O (g26052), .I1 (g25941), .I2 (g21087));
AN2X1 gate18257(.O (g26053), .I1 (g758), .I2 (g25306));
AN2X1 gate18258(.O (g26054), .I1 (g25944), .I2 (g21099));
AN2X1 gate18259(.O (g26060), .I1 (g25943), .I2 (g21108));
AN2X1 gate18260(.O (g26061), .I1 (g1444), .I2 (g25315));
AN2X1 gate18261(.O (g26062), .I1 (g25947), .I2 (g21113));
AN2X1 gate18262(.O (g26067), .I1 (g25946), .I2 (g21125));
AN2X1 gate18263(.O (g26068), .I1 (g2138), .I2 (g25324));
AN2X1 gate18264(.O (g26069), .I1 (g25949), .I2 (g21130));
AN2X1 gate18265(.O (g26074), .I1 (g25948), .I2 (g21144));
AN2X1 gate18266(.O (g26075), .I1 (g74), .I2 (g25698));
AN2X1 gate18267(.O (g26080), .I1 (g25950), .I2 (g21164));
AN2X1 gate18268(.O (g26082), .I1 (g762), .I2 (g25771));
AN2X1 gate18269(.O (g26085), .I1 (g1448), .I2 (g25825));
AN2X1 gate18270(.O (g26091), .I1 (g2142), .I2 (g25860));
AN2X1 gate18271(.O (g26157), .I1 (g21825), .I2 (g25630));
AN2X1 gate18272(.O (g26158), .I1 (g679), .I2 (g25937));
AN2X1 gate18273(.O (g26163), .I1 (g1365), .I2 (g25939));
AN2X1 gate18274(.O (g26166), .I1 (g686), .I2 (g25454));
AN2X1 gate18275(.O (g26171), .I1 (g2059), .I2 (g25942));
AN2X1 gate18276(.O (g26186), .I1 (g1372), .I2 (g25458));
AN2X1 gate18277(.O (g26188), .I1 (g2753), .I2 (g25945));
AN2X1 gate18278(.O (g26207), .I1 (g2066), .I2 (g25463));
AN2X1 gate18279(.O (g26212), .I1 (g4217), .I2 (g25467));
AN2X1 gate18280(.O (g26213), .I1 (g25895), .I2 (g9306));
AN2X1 gate18281(.O (g26231), .I1 (g2760), .I2 (g25472));
AN2X1 gate18282(.O (g26233), .I1 (g4340), .I2 (g25476));
AN2X1 gate18283(.O (g26234), .I1 (g4343), .I2 (g25479));
AN2X1 gate18284(.O (g26235), .I1 (g25895), .I2 (g9368));
AN2X1 gate18285(.O (g26236), .I1 (g25899), .I2 (g9371));
AN2X1 gate18286(.O (g26243), .I1 (g4372), .I2 (g25484));
AN2X1 gate18287(.O (g26244), .I1 (g25903), .I2 (g9387));
AN2X1 gate18288(.O (g26257), .I1 (g4465), .I2 (g25493));
AN2X1 gate18289(.O (g26258), .I1 (g4468), .I2 (g25496));
AN2X1 gate18290(.O (g26259), .I1 (g4471), .I2 (g25499));
AN2X1 gate18291(.O (g26260), .I1 (g25254), .I2 (g17649));
AN2X1 gate18292(.O (g26261), .I1 (g25895), .I2 (g9443));
AN2X1 gate18293(.O (g26262), .I1 (g25899), .I2 (g9446));
AN2X1 gate18294(.O (g26263), .I1 (g4476), .I2 (g25502));
AN2X1 gate18295(.O (g26268), .I1 (g4509), .I2 (g25507));
AN2X1 gate18296(.O (g26269), .I1 (g4512), .I2 (g25510));
AN2X1 gate18297(.O (g26270), .I1 (g25903), .I2 (g9465));
AN2X1 gate18298(.O (g26271), .I1 (g25907), .I2 (g9468));
AN2X1 gate18299(.O (g26278), .I1 (g4541), .I2 (g25515));
AN2X1 gate18300(.O (g26279), .I1 (g25911), .I2 (g9484));
AN2X1 gate18301(.O (g26288), .I1 (g4592), .I2 (g25524));
AN2X1 gate18302(.O (g26289), .I1 (g4595), .I2 (g25527));
AN2X1 gate18303(.O (g26290), .I1 (g4598), .I2 (g25530));
AN2X1 gate18304(.O (g26291), .I1 (g25899), .I2 (g9524));
AN2X1 gate18305(.O (g26292), .I1 (g4603), .I2 (g25533));
AN2X1 gate18306(.O (g26293), .I1 (g4606), .I2 (g25536));
AN2X1 gate18307(.O (g26298), .I1 (g4641), .I2 (g25540));
AN2X1 gate18308(.O (g26299), .I1 (g4644), .I2 (g25543));
AN2X1 gate18309(.O (g26300), .I1 (g4647), .I2 (g25546));
AN2X1 gate18310(.O (g26301), .I1 (g25258), .I2 (g17749));
AN2X1 gate18311(.O (g26302), .I1 (g25903), .I2 (g9585));
AN2X1 gate18312(.O (g26303), .I1 (g25907), .I2 (g9588));
AN2X1 gate18313(.O (g26307), .I1 (g4652), .I2 (g25549));
AN2X1 gate18314(.O (g26309), .I1 (g4685), .I2 (g25554));
AN2X1 gate18315(.O (g26310), .I1 (g4688), .I2 (g25557));
AN2X1 gate18316(.O (g26311), .I1 (g25911), .I2 (g9607));
AN2X1 gate18317(.O (g26312), .I1 (g25915), .I2 (g9610));
AN2X1 gate18318(.O (g26316), .I1 (g4717), .I2 (g25562));
AN2X1 gate18319(.O (g26317), .I1 (g25919), .I2 (g9626));
AN2X1 gate18320(.O (g26318), .I1 (g4737), .I2 (g25573));
AN2X1 gate18321(.O (g26319), .I1 (g4740), .I2 (g25576));
AN2X1 gate18322(.O (g26324), .I1 (g4743), .I2 (g25579));
AN2X1 gate18323(.O (g26325), .I1 (g4746), .I2 (g25582));
AN2X1 gate18324(.O (g26326), .I1 (g4749), .I2 (g25585));
AN2X1 gate18325(.O (g26332), .I1 (g4769), .I2 (g25590));
AN2X1 gate18326(.O (g26333), .I1 (g4772), .I2 (g25593));
AN2X1 gate18327(.O (g26334), .I1 (g4775), .I2 (g25596));
AN2X1 gate18328(.O (g26335), .I1 (g25907), .I2 (g9666));
AN2X1 gate18329(.O (g26339), .I1 (g4780), .I2 (g25599));
AN2X1 gate18330(.O (g26340), .I1 (g4783), .I2 (g25602));
AN2X1 gate18331(.O (g26342), .I1 (g4818), .I2 (g25606));
AN2X1 gate18332(.O (g26343), .I1 (g4821), .I2 (g25609));
AN2X1 gate18333(.O (g26344), .I1 (g4824), .I2 (g25612));
AN2X1 gate18334(.O (g26345), .I1 (g25261), .I2 (g17850));
AN2X1 gate18335(.O (g26346), .I1 (g25911), .I2 (g9727));
AN2X1 gate18336(.O (g26347), .I1 (g25915), .I2 (g9730));
AN2X1 gate18337(.O (g26348), .I1 (g4829), .I2 (g25615));
AN2X1 gate18338(.O (g26350), .I1 (g4862), .I2 (g25620));
AN2X1 gate18339(.O (g26351), .I1 (g4865), .I2 (g25623));
AN2X1 gate18340(.O (g26352), .I1 (g25919), .I2 (g9749));
AN2X1 gate18341(.O (g26353), .I1 (g25923), .I2 (g9752));
AN2X1 gate18342(.O (g26357), .I1 (g4882), .I2 (g25634));
AN2X1 gate18343(.O (g26361), .I1 (g4888), .I2 (g25637));
AN2X1 gate18344(.O (g26362), .I1 (g4891), .I2 (g25640));
AN2X1 gate18345(.O (g26363), .I1 (g4894), .I2 (g25643));
AN2X1 gate18346(.O (g26365), .I1 (g4913), .I2 (g25652));
AN2X1 gate18347(.O (g26366), .I1 (g4916), .I2 (g25655));
AN2X1 gate18348(.O (g26371), .I1 (g4919), .I2 (g25658));
AN2X1 gate18349(.O (g26372), .I1 (g4922), .I2 (g25661));
AN2X1 gate18350(.O (g26373), .I1 (g4925), .I2 (g25664));
AN2X1 gate18351(.O (g26379), .I1 (g4945), .I2 (g25669));
AN2X1 gate18352(.O (g26380), .I1 (g4948), .I2 (g25672));
AN2X1 gate18353(.O (g26381), .I1 (g4951), .I2 (g25675));
AN2X1 gate18354(.O (g26382), .I1 (g25915), .I2 (g9812));
AN2X1 gate18355(.O (g26383), .I1 (g4956), .I2 (g25678));
AN2X1 gate18356(.O (g26384), .I1 (g4959), .I2 (g25681));
AN2X1 gate18357(.O (g26386), .I1 (g4994), .I2 (g25685));
AN2X1 gate18358(.O (g26387), .I1 (g4997), .I2 (g25688));
AN2X1 gate18359(.O (g26388), .I1 (g5000), .I2 (g25691));
AN2X1 gate18360(.O (g26389), .I1 (g25264), .I2 (g17962));
AN2X1 gate18361(.O (g26390), .I1 (g25919), .I2 (g9873));
AN2X1 gate18362(.O (g26391), .I1 (g25923), .I2 (g9876));
AN2X1 gate18363(.O (g26392), .I1 (g5005), .I2 (g25694));
AN2X1 gate18364(.O (g26396), .I1 (g5027), .I2 (g25700));
AN2X1 gate18365(.O (g26397), .I1 (g5030), .I2 (g25703));
AN2X1 gate18366(.O (g26400), .I1 (g5041), .I2 (g25711));
AN2X1 gate18367(.O (g26404), .I1 (g5047), .I2 (g25714));
AN2X1 gate18368(.O (g26405), .I1 (g5050), .I2 (g25717));
AN2X1 gate18369(.O (g26406), .I1 (g5053), .I2 (g25720));
AN2X1 gate18370(.O (g26408), .I1 (g5072), .I2 (g25729));
AN2X1 gate18371(.O (g26409), .I1 (g5075), .I2 (g25732));
AN2X1 gate18372(.O (g26414), .I1 (g5078), .I2 (g25735));
AN2X1 gate18373(.O (g26415), .I1 (g5081), .I2 (g25738));
AN2X1 gate18374(.O (g26416), .I1 (g5084), .I2 (g25741));
AN2X1 gate18375(.O (g26422), .I1 (g5104), .I2 (g25746));
AN2X1 gate18376(.O (g26423), .I1 (g5107), .I2 (g25749));
AN2X1 gate18377(.O (g26424), .I1 (g5110), .I2 (g25752));
AN2X1 gate18378(.O (g26425), .I1 (g25923), .I2 (g9958));
AN2X1 gate18379(.O (g26426), .I1 (g5115), .I2 (g25755));
AN2X1 gate18380(.O (g26427), .I1 (g5118), .I2 (g25758));
AN2X1 gate18381(.O (g26432), .I1 (g5145), .I2 (g25767));
AN2X1 gate18382(.O (g26437), .I1 (g5156), .I2 (g25773));
AN2X1 gate18383(.O (g26438), .I1 (g5159), .I2 (g25776));
AN2X1 gate18384(.O (g26441), .I1 (g5170), .I2 (g25784));
AN2X1 gate18385(.O (g26445), .I1 (g5176), .I2 (g25787));
AN2X1 gate18386(.O (g26446), .I1 (g5179), .I2 (g25790));
AN2X1 gate18387(.O (g26447), .I1 (g5182), .I2 (g25793));
AN2X1 gate18388(.O (g26449), .I1 (g5201), .I2 (g25802));
AN2X1 gate18389(.O (g26450), .I1 (g5204), .I2 (g25805));
AN2X1 gate18390(.O (g26455), .I1 (g5207), .I2 (g25808));
AN2X1 gate18391(.O (g26456), .I1 (g5210), .I2 (g25811));
AN2X1 gate18392(.O (g26457), .I1 (g5213), .I2 (g25814));
AN2X1 gate18393(.O (g26464), .I1 (g5238), .I2 (g25821));
AN2X1 gate18394(.O (g26469), .I1 (g5249), .I2 (g25827));
AN2X1 gate18395(.O (g26470), .I1 (g5252), .I2 (g25830));
AN2X1 gate18396(.O (g26473), .I1 (g5263), .I2 (g25838));
AN2X1 gate18397(.O (g26477), .I1 (g5269), .I2 (g25841));
AN2X1 gate18398(.O (g26478), .I1 (g5272), .I2 (g25844));
AN2X1 gate18399(.O (g26479), .I1 (g5275), .I2 (g25847));
AN2X1 gate18400(.O (g26488), .I1 (g5301), .I2 (g25856));
AN2X1 gate18401(.O (g26493), .I1 (g5312), .I2 (g25862));
AN2X1 gate18402(.O (g26494), .I1 (g5315), .I2 (g25865));
AN2X1 gate18403(.O (g26504), .I1 (g5338), .I2 (g25877));
AN2X1 gate18404(.O (g26663), .I1 (g25274), .I2 (g21066));
AN2X1 gate18405(.O (g26668), .I1 (g25283), .I2 (g21076));
AN2X1 gate18406(.O (g26673), .I1 (g12431), .I2 (g25318));
AN2X1 gate18407(.O (g26674), .I1 (g25291), .I2 (g21090));
AN2X1 gate18408(.O (g26754), .I1 (g14657), .I2 (g26508));
AN2X1 gate18409(.O (g26755), .I1 (g26083), .I2 (g22239));
AN2X1 gate18410(.O (g26756), .I1 (g26113), .I2 (g22240));
AN3X1 gate18411(.O (g26758), .I1 (g16614), .I2 (g26521), .I3 (g13637));
AN2X1 gate18412(.O (g26759), .I1 (g26356), .I2 (g19251));
AN2X1 gate18413(.O (g26760), .I1 (g26137), .I2 (g22256));
AN2X1 gate18414(.O (g26761), .I1 (g26154), .I2 (g22257));
AN2X1 gate18415(.O (g26763), .I1 (g14691), .I2 (g26516));
AN3X1 gate18416(.O (g26764), .I1 (g16632), .I2 (g26525), .I3 (g13649));
AN2X1 gate18417(.O (g26765), .I1 (g26399), .I2 (g19265));
AN2X1 gate18418(.O (g26766), .I1 (g14725), .I2 (g26521));
AN2X1 gate18419(.O (g26767), .I1 (g26087), .I2 (g22287));
AN2X1 gate18420(.O (g26768), .I1 (g26440), .I2 (g19280));
AN2X1 gate18421(.O (g26769), .I1 (g14753), .I2 (g26525));
AN2X1 gate18422(.O (g26770), .I1 (g26059), .I2 (g19287));
AN3X1 gate18423(.O (g26771), .I1 (g24912), .I2 (g26508), .I3 (g13614));
AN2X1 gate18424(.O (g26773), .I1 (g26145), .I2 (g22303));
AN2X1 gate18425(.O (g26774), .I1 (g26472), .I2 (g19299));
AN2X1 gate18426(.O (g26775), .I1 (g26099), .I2 (g22318));
AN2X1 gate18427(.O (g26777), .I1 (g26066), .I2 (g19305));
AN3X1 gate18428(.O (g26778), .I1 (g24929), .I2 (g26516), .I3 (g13626));
AN2X1 gate18429(.O (g26780), .I1 (g26119), .I2 (g16622));
AN2X1 gate18430(.O (g26783), .I1 (g26073), .I2 (g19326));
AN3X1 gate18431(.O (g26784), .I1 (g24941), .I2 (g26521), .I3 (g13637));
AN2X1 gate18432(.O (g26787), .I1 (g26129), .I2 (g16636));
AN2X1 gate18433(.O (g26790), .I1 (g26079), .I2 (g19353));
AN3X1 gate18434(.O (g26791), .I1 (g24952), .I2 (g26525), .I3 (g13649));
AN2X1 gate18435(.O (g26794), .I1 (g26143), .I2 (g16647));
AN2X1 gate18436(.O (g26797), .I1 (g26148), .I2 (g16659));
AN2X1 gate18437(.O (g26829), .I1 (g5623), .I2 (g26209));
AN2X1 gate18438(.O (g26833), .I1 (g5651), .I2 (g26237));
AN2X1 gate18439(.O (g26842), .I1 (g5689), .I2 (g26275));
AN2X1 gate18440(.O (g26845), .I1 (g5664), .I2 (g26056));
AN2X1 gate18441(.O (g26851), .I1 (g5741), .I2 (g26313));
AN2X1 gate18442(.O (g26853), .I1 (g5716), .I2 (g26063));
AN2X1 gate18443(.O (g26860), .I1 (g5774), .I2 (g26070));
AN2X1 gate18444(.O (g26866), .I1 (g5833), .I2 (g26076));
AN2X1 gate18445(.O (g26955), .I1 (g6157), .I2 (g26533));
AN2X1 gate18446(.O (g26958), .I1 (g6184), .I2 (g26538));
AN2X1 gate18447(.O (g26961), .I1 (g13907), .I2 (g26175));
AN2X1 gate18448(.O (g26962), .I1 (g6180), .I2 (g26178));
AN2X1 gate18449(.O (g26963), .I1 (g6216), .I2 (g26539));
AN2X1 gate18450(.O (g26965), .I1 (g23320), .I2 (g26540));
AN2X1 gate18451(.O (g26966), .I1 (g13963), .I2 (g26196));
AN2X1 gate18452(.O (g26967), .I1 (g6212), .I2 (g26202));
AN2X1 gate18453(.O (g26968), .I1 (g6305), .I2 (g26542));
AN2X1 gate18454(.O (g26969), .I1 (g23320), .I2 (g26543));
AN2X1 gate18455(.O (g26970), .I1 (g21976), .I2 (g26544));
AN2X1 gate18456(.O (g26971), .I1 (g23325), .I2 (g26546));
AN2X1 gate18457(.O (g26972), .I1 (g14033), .I2 (g26223));
AN2X1 gate18458(.O (g26973), .I1 (g6301), .I2 (g26226));
AN2X1 gate18459(.O (g26977), .I1 (g23320), .I2 (g26550));
AN2X1 gate18460(.O (g26978), .I1 (g21976), .I2 (g26551));
AN2X1 gate18461(.O (g26979), .I1 (g23331), .I2 (g26552));
AN2X1 gate18462(.O (g26980), .I1 (g23360), .I2 (g26554));
AN2X1 gate18463(.O (g26981), .I1 (g23325), .I2 (g26555));
AN2X1 gate18464(.O (g26982), .I1 (g21983), .I2 (g26556));
AN2X1 gate18465(.O (g26984), .I1 (g23335), .I2 (g26558));
AN2X1 gate18466(.O (g26985), .I1 (g14124), .I2 (g26251));
AN2X1 gate18467(.O (g26986), .I1 (g6438), .I2 (g26254));
AN2X1 gate18468(.O (g26993), .I1 (g21976), .I2 (g26561));
AN2X1 gate18469(.O (g26994), .I1 (g23331), .I2 (g26562));
AN2X1 gate18470(.O (g26995), .I1 (g21991), .I2 (g26563));
AN2X1 gate18471(.O (g26996), .I1 (g23360), .I2 (g26564));
AN2X1 gate18472(.O (g26997), .I1 (g22050), .I2 (g26565));
AN2X1 gate18473(.O (g26998), .I1 (g23325), .I2 (g26566));
AN2X1 gate18474(.O (g26999), .I1 (g21983), .I2 (g26567));
AN2X1 gate18475(.O (g27000), .I1 (g23340), .I2 (g26568));
AN2X1 gate18476(.O (g27001), .I1 (g23364), .I2 (g26570));
AN2X1 gate18477(.O (g27002), .I1 (g23335), .I2 (g26571));
AN2X1 gate18478(.O (g27003), .I1 (g21996), .I2 (g26572));
AN2X1 gate18479(.O (g27004), .I1 (g23344), .I2 (g26574));
AN2X1 gate18480(.O (g27005), .I1 (g23331), .I2 (g26578));
AN2X1 gate18481(.O (g27006), .I1 (g21991), .I2 (g26579));
AN2X1 gate18482(.O (g27007), .I1 (g23360), .I2 (g26580));
AN2X1 gate18483(.O (g27008), .I1 (g22050), .I2 (g26581));
AN2X1 gate18484(.O (g27009), .I1 (g23368), .I2 (g26582));
AN2X1 gate18485(.O (g27016), .I1 (g21983), .I2 (g26584));
AN2X1 gate18486(.O (g27017), .I1 (g23340), .I2 (g26585));
AN2X1 gate18487(.O (g27018), .I1 (g22005), .I2 (g26586));
AN2X1 gate18488(.O (g27019), .I1 (g23364), .I2 (g26587));
AN2X1 gate18489(.O (g27020), .I1 (g22069), .I2 (g26588));
AN2X1 gate18490(.O (g27021), .I1 (g23335), .I2 (g26589));
AN2X1 gate18491(.O (g27022), .I1 (g21996), .I2 (g26590));
AN2X1 gate18492(.O (g27023), .I1 (g23349), .I2 (g26591));
AN2X1 gate18493(.O (g27024), .I1 (g23372), .I2 (g26593));
AN2X1 gate18494(.O (g27025), .I1 (g23344), .I2 (g26594));
AN2X1 gate18495(.O (g27026), .I1 (g22009), .I2 (g26595));
AN2X1 gate18496(.O (g27027), .I1 (g21991), .I2 (g26598));
AN2X1 gate18497(.O (g27028), .I1 (g22050), .I2 (g26599));
AN2X1 gate18498(.O (g27029), .I1 (g23368), .I2 (g26600));
AN2X1 gate18499(.O (g27030), .I1 (g22083), .I2 (g26601));
AN2X1 gate18500(.O (g27031), .I1 (g23340), .I2 (g26602));
AN2X1 gate18501(.O (g27032), .I1 (g22005), .I2 (g26603));
AN2X1 gate18502(.O (g27033), .I1 (g23364), .I2 (g26604));
AN2X1 gate18503(.O (g27034), .I1 (g22069), .I2 (g26605));
AN2X1 gate18504(.O (g27035), .I1 (g23377), .I2 (g26606));
AN2X1 gate18505(.O (g27042), .I1 (g21996), .I2 (g26608));
AN2X1 gate18506(.O (g27043), .I1 (g23349), .I2 (g26609));
AN2X1 gate18507(.O (g27044), .I1 (g22016), .I2 (g26610));
AN2X1 gate18508(.O (g27045), .I1 (g23372), .I2 (g26611));
AN2X1 gate18509(.O (g27046), .I1 (g22093), .I2 (g26612));
AN2X1 gate18510(.O (g27047), .I1 (g23344), .I2 (g26613));
AN2X1 gate18511(.O (g27048), .I1 (g22009), .I2 (g26614));
AN2X1 gate18512(.O (g27049), .I1 (g23353), .I2 (g26615));
AN2X1 gate18513(.O (g27050), .I1 (g23381), .I2 (g26617));
AN2X1 gate18514(.O (g27052), .I1 (g4885), .I2 (g26358));
AN2X1 gate18515(.O (g27053), .I1 (g23368), .I2 (g26619));
AN2X1 gate18516(.O (g27054), .I1 (g22083), .I2 (g26620));
AN2X1 gate18517(.O (g27055), .I1 (g22005), .I2 (g26621));
AN2X1 gate18518(.O (g27056), .I1 (g22069), .I2 (g26622));
AN2X1 gate18519(.O (g27057), .I1 (g23377), .I2 (g26623));
AN2X1 gate18520(.O (g27058), .I1 (g22108), .I2 (g26624));
AN2X1 gate18521(.O (g27059), .I1 (g23349), .I2 (g26625));
AN2X1 gate18522(.O (g27060), .I1 (g22016), .I2 (g26626));
AN2X1 gate18523(.O (g27061), .I1 (g23372), .I2 (g26627));
AN2X1 gate18524(.O (g27062), .I1 (g22093), .I2 (g26628));
AN2X1 gate18525(.O (g27063), .I1 (g23388), .I2 (g26629));
AN2X1 gate18526(.O (g27070), .I1 (g22009), .I2 (g26631));
AN2X1 gate18527(.O (g27071), .I1 (g23353), .I2 (g26632));
AN2X1 gate18528(.O (g27072), .I1 (g22021), .I2 (g26633));
AN2X1 gate18529(.O (g27073), .I1 (g23381), .I2 (g26634));
AN2X1 gate18530(.O (g27074), .I1 (g22118), .I2 (g26635));
AN2X1 gate18531(.O (g27076), .I1 (g5024), .I2 (g26393));
AN2X1 gate18532(.O (g27077), .I1 (g22083), .I2 (g26636));
AN2X1 gate18533(.O (g27079), .I1 (g5044), .I2 (g26401));
AN2X1 gate18534(.O (g27080), .I1 (g23377), .I2 (g26637));
AN2X1 gate18535(.O (g27081), .I1 (g22108), .I2 (g26638));
AN2X1 gate18536(.O (g27082), .I1 (g22016), .I2 (g26639));
AN2X1 gate18537(.O (g27083), .I1 (g22093), .I2 (g26640));
AN2X1 gate18538(.O (g27084), .I1 (g23388), .I2 (g26641));
AN2X1 gate18539(.O (g27085), .I1 (g22134), .I2 (g26642));
AN2X1 gate18540(.O (g27086), .I1 (g23353), .I2 (g26643));
AN2X1 gate18541(.O (g27087), .I1 (g22021), .I2 (g26644));
AN2X1 gate18542(.O (g27088), .I1 (g23381), .I2 (g26645));
AN2X1 gate18543(.O (g27089), .I1 (g22118), .I2 (g26646));
AN2X1 gate18544(.O (g27090), .I1 (g23395), .I2 (g26647));
AN2X1 gate18545(.O (g27091), .I1 (g5142), .I2 (g26429));
AN2X1 gate18546(.O (g27092), .I1 (g5153), .I2 (g26434));
AN2X1 gate18547(.O (g27093), .I1 (g22108), .I2 (g26648));
AN2X1 gate18548(.O (g27095), .I1 (g5173), .I2 (g26442));
AN2X1 gate18549(.O (g27096), .I1 (g23388), .I2 (g26649));
AN2X1 gate18550(.O (g27097), .I1 (g22134), .I2 (g26650));
AN2X1 gate18551(.O (g27098), .I1 (g22021), .I2 (g26651));
AN2X1 gate18552(.O (g27099), .I1 (g22118), .I2 (g26652));
AN2X1 gate18553(.O (g27100), .I1 (g23395), .I2 (g26653));
AN2X1 gate18554(.O (g27101), .I1 (g22157), .I2 (g26654));
AN2X1 gate18555(.O (g27103), .I1 (g5235), .I2 (g26461));
AN2X1 gate18556(.O (g27104), .I1 (g5246), .I2 (g26466));
AN2X1 gate18557(.O (g27105), .I1 (g22134), .I2 (g26656));
AN2X1 gate18558(.O (g27107), .I1 (g5266), .I2 (g26474));
AN2X1 gate18559(.O (g27108), .I1 (g23395), .I2 (g26657));
AN2X1 gate18560(.O (g27109), .I1 (g22157), .I2 (g26658));
AN2X1 gate18561(.O (g27110), .I1 (g5298), .I2 (g26485));
AN2X1 gate18562(.O (g27111), .I1 (g5309), .I2 (g26490));
AN2X1 gate18563(.O (g27112), .I1 (g22157), .I2 (g26662));
AN2X1 gate18564(.O (g27115), .I1 (g5335), .I2 (g26501));
AN2X1 gate18565(.O (g27178), .I1 (g26110), .I2 (g22213));
AN3X1 gate18566(.O (g27181), .I1 (g16570), .I2 (g26508), .I3 (g13614));
AN2X1 gate18567(.O (g27182), .I1 (g26151), .I2 (g22217));
AN2X1 gate18568(.O (g27185), .I1 (g26126), .I2 (g22230));
AN3X1 gate18569(.O (g27187), .I1 (g16594), .I2 (g26516), .I3 (g13626));
AN2X1 gate18570(.O (g27240), .I1 (g26905), .I2 (g22241));
AN2X1 gate18571(.O (g27241), .I1 (g10730), .I2 (g26934));
AN2X1 gate18572(.O (g27242), .I1 (g26793), .I2 (g8357));
AN2X1 gate18573(.O (g27244), .I1 (g26914), .I2 (g22258));
AN2X1 gate18574(.O (g27245), .I1 (g26877), .I2 (g22286));
AN2X1 gate18575(.O (g27246), .I1 (g26988), .I2 (g16676));
AN2X1 gate18576(.O (g27247), .I1 (g27011), .I2 (g16702));
AN2X1 gate18577(.O (g27248), .I1 (g27037), .I2 (g16733));
AN2X1 gate18578(.O (g27249), .I1 (g27065), .I2 (g16775));
AN2X1 gate18579(.O (g27355), .I1 (g61), .I2 (g26837));
AN2X1 gate18580(.O (g27356), .I1 (g65), .I2 (g26987));
AN2X1 gate18581(.O (g27358), .I1 (g749), .I2 (g26846));
AN2X1 gate18582(.O (g27359), .I1 (g753), .I2 (g27010));
AN2X1 gate18583(.O (g27364), .I1 (g1435), .I2 (g26855));
AN2X1 gate18584(.O (g27365), .I1 (g1439), .I2 (g27036));
AN2X1 gate18585(.O (g27370), .I1 (g27126), .I2 (g8874));
AN2X1 gate18586(.O (g27371), .I1 (g2129), .I2 (g26861));
AN2X1 gate18587(.O (g27372), .I1 (g2133), .I2 (g27064));
AN2X1 gate18588(.O (g27394), .I1 (g17802), .I2 (g27134));
AN2X1 gate18589(.O (g27396), .I1 (g692), .I2 (g27135));
AN2X1 gate18590(.O (g27407), .I1 (g17914), .I2 (g27136));
AN2X1 gate18591(.O (g27409), .I1 (g1378), .I2 (g27137));
AN2X1 gate18592(.O (g27425), .I1 (g18025), .I2 (g27138));
AN2X1 gate18593(.O (g27427), .I1 (g2072), .I2 (g27139));
AN2X1 gate18594(.O (g27446), .I1 (g18142), .I2 (g27141));
AN2X1 gate18595(.O (g27448), .I1 (g2766), .I2 (g27142));
AN2X1 gate18596(.O (g27495), .I1 (g23945), .I2 (g27146));
AN2X1 gate18597(.O (g27509), .I1 (g23945), .I2 (g27148));
AN2X1 gate18598(.O (g27516), .I1 (g23974), .I2 (g27151));
AN2X1 gate18599(.O (g27530), .I1 (g23945), .I2 (g27153));
AN2X1 gate18600(.O (g27534), .I1 (g23974), .I2 (g27155));
AN2X1 gate18601(.O (g27541), .I1 (g24004), .I2 (g27159));
AN2X1 gate18602(.O (g27552), .I1 (g23974), .I2 (g27162));
AN2X1 gate18603(.O (g27554), .I1 (g24004), .I2 (g27164));
AN2X1 gate18604(.O (g27561), .I1 (g24038), .I2 (g27167));
AN2X1 gate18605(.O (g27568), .I1 (g24004), .I2 (g27172));
AN2X1 gate18606(.O (g27570), .I1 (g24038), .I2 (g27173));
AN2X1 gate18607(.O (g27578), .I1 (g24038), .I2 (g27177));
AN2X1 gate18608(.O (g27656), .I1 (g26796), .I2 (g11004));
AN2X1 gate18609(.O (g27657), .I1 (g27114), .I2 (g11051));
AN2X1 gate18610(.O (g27659), .I1 (g27132), .I2 (g11114));
AN2X1 gate18611(.O (g27660), .I1 (g26835), .I2 (g11117));
AN2X1 gate18612(.O (g27661), .I1 (g26841), .I2 (g11173));
AN2X1 gate18613(.O (g27666), .I1 (g26849), .I2 (g11243));
AN2X1 gate18614(.O (g27671), .I1 (g26885), .I2 (g22212));
AN2X1 gate18615(.O (g27673), .I1 (g26854), .I2 (g11312));
AN2X1 gate18616(.O (g27679), .I1 (g26782), .I2 (g11386));
AN2X1 gate18617(.O (g27680), .I1 (g26983), .I2 (g11392));
AN2X1 gate18618(.O (g27681), .I1 (g26788), .I2 (g11456));
AN2X1 gate18619(.O (g27719), .I1 (g27496), .I2 (g20649));
AN2X1 gate18620(.O (g27720), .I1 (g27481), .I2 (g20652));
AN2X1 gate18621(.O (g27721), .I1 (g27579), .I2 (g20655));
AN2X1 gate18622(.O (g27723), .I1 (g27464), .I2 (g20679));
AN2X1 gate18623(.O (g27725), .I1 (g27532), .I2 (g20704));
AN2X1 gate18624(.O (g27726), .I1 (g27531), .I2 (g20732));
AN2X1 gate18625(.O (g27727), .I1 (g27414), .I2 (g19301));
AN2X1 gate18626(.O (g27728), .I1 (g27564), .I2 (g20766));
AN2X1 gate18627(.O (g27729), .I1 (g27435), .I2 (g19322));
AN2X1 gate18628(.O (g27730), .I1 (g27454), .I2 (g19349));
AN2X1 gate18629(.O (g27731), .I1 (g27470), .I2 (g19383));
AN2X1 gate18630(.O (g27732), .I1 (g27492), .I2 (g16758));
AN2X1 gate18631(.O (g27733), .I1 (g27513), .I2 (g16785));
AN2X1 gate18632(.O (g27734), .I1 (g27538), .I2 (g16814));
AN2X1 gate18633(.O (g27737), .I1 (g27558), .I2 (g16832));
AN2X1 gate18634(.O (g27770), .I1 (g5642), .I2 (g27449));
AN2X1 gate18635(.O (g27772), .I1 (g5680), .I2 (g27465));
AN2X1 gate18636(.O (g27773), .I1 (g5732), .I2 (g27484));
AN2X1 gate18637(.O (g27774), .I1 (g5702), .I2 (g27361));
AN2X1 gate18638(.O (g27775), .I1 (g5790), .I2 (g27506));
AN2X1 gate18639(.O (g27779), .I1 (g5760), .I2 (g27367));
AN2X1 gate18640(.O (g27783), .I1 (g5819), .I2 (g27373));
AN2X1 gate18641(.O (g27790), .I1 (g5875), .I2 (g27376));
AN2X1 gate18642(.O (g27904), .I1 (g13873), .I2 (g27387));
AN2X1 gate18643(.O (g27908), .I1 (g13886), .I2 (g27391));
AN2X1 gate18644(.O (g27909), .I1 (g13895), .I2 (g27397));
AN2X1 gate18645(.O (g27913), .I1 (g4017), .I2 (g27401));
AN2X1 gate18646(.O (g27914), .I1 (g13927), .I2 (g27404));
AN2X1 gate18647(.O (g27915), .I1 (g13936), .I2 (g27410));
AN2X1 gate18648(.O (g27922), .I1 (g4112), .I2 (g27416));
AN2X1 gate18649(.O (g27923), .I1 (g4144), .I2 (g27419));
AN2X1 gate18650(.O (g27924), .I1 (g13983), .I2 (g27422));
AN2X1 gate18651(.O (g27926), .I1 (g13992), .I2 (g27428));
AN2X1 gate18652(.O (g27931), .I1 (g4221), .I2 (g27432));
AN2X1 gate18653(.O (g27935), .I1 (g4251), .I2 (g27437));
AN2X1 gate18654(.O (g27936), .I1 (g4283), .I2 (g27440));
AN2X1 gate18655(.O (g27938), .I1 (g14053), .I2 (g27443));
AN2X1 gate18656(.O (g27945), .I1 (g4376), .I2 (g27451));
AN2X1 gate18657(.O (g27949), .I1 (g4406), .I2 (g27456));
AN2X1 gate18658(.O (g27951), .I1 (g4438), .I2 (g27459));
AN2X1 gate18659(.O (g27963), .I1 (g4545), .I2 (g27467));
AN2X1 gate18660(.O (g27968), .I1 (g4575), .I2 (g27472));
AN2X1 gate18661(.O (g27970), .I1 (g14238), .I2 (g27475));
AN2X1 gate18662(.O (g27984), .I1 (g4721), .I2 (g27486));
AN2X1 gate18663(.O (g27985), .I1 (g14342), .I2 (g27489));
AN2X1 gate18664(.O (g27991), .I1 (g14360), .I2 (g27498));
AN2X1 gate18665(.O (g28008), .I1 (g27590), .I2 (g9770));
AN2X1 gate18666(.O (g28009), .I1 (g14454), .I2 (g27510));
AN2X1 gate18667(.O (g28015), .I1 (g14472), .I2 (g27518));
AN2X1 gate18668(.O (g28027), .I1 (g27590), .I2 (g9895));
AN2X1 gate18669(.O (g28028), .I1 (g27595), .I2 (g9898));
AN2X1 gate18670(.O (g28035), .I1 (g27599), .I2 (g9916));
AN2X1 gate18671(.O (g28036), .I1 (g14541), .I2 (g27535));
AN2X1 gate18672(.O (g28042), .I1 (g14559), .I2 (g27543));
AN2X1 gate18673(.O (g28050), .I1 (g27590), .I2 (g10018));
AN2X1 gate18674(.O (g28051), .I1 (g27595), .I2 (g10021));
AN2X1 gate18675(.O (g28057), .I1 (g27599), .I2 (g10049));
AN2X1 gate18676(.O (g28058), .I1 (g27604), .I2 (g10052));
AN2X1 gate18677(.O (g28065), .I1 (g27608), .I2 (g10070));
AN2X1 gate18678(.O (g28066), .I1 (g14596), .I2 (g27555));
AN2X1 gate18679(.O (g28073), .I1 (g27595), .I2 (g10109));
AN2X1 gate18680(.O (g28079), .I1 (g27599), .I2 (g10127));
AN2X1 gate18681(.O (g28080), .I1 (g27604), .I2 (g10130));
AN2X1 gate18682(.O (g28086), .I1 (g27608), .I2 (g10158));
AN2X1 gate18683(.O (g28087), .I1 (g27613), .I2 (g10161));
AN2X1 gate18684(.O (g28094), .I1 (g27617), .I2 (g10179));
AN2X1 gate18685(.O (g28098), .I1 (g27604), .I2 (g10214));
AN2X1 gate18686(.O (g28104), .I1 (g27608), .I2 (g10232));
AN2X1 gate18687(.O (g28105), .I1 (g27613), .I2 (g10235));
AN2X1 gate18688(.O (g28111), .I1 (g27617), .I2 (g10263));
AN2X1 gate18689(.O (g28112), .I1 (g27622), .I2 (g10266));
AN2X1 gate18690(.O (g28116), .I1 (g27613), .I2 (g10316));
AN2X1 gate18691(.O (g28122), .I1 (g27617), .I2 (g10334));
AN2X1 gate18692(.O (g28123), .I1 (g27622), .I2 (g10337));
AN2X1 gate18693(.O (g28127), .I1 (g27622), .I2 (g10409));
AN2X1 gate18694(.O (g28171), .I1 (g27349), .I2 (g10898));
AN2X1 gate18695(.O (g28176), .I1 (g27349), .I2 (g10940));
AN2X1 gate18696(.O (g28188), .I1 (g27349), .I2 (g11008));
AN2X1 gate18697(.O (g28193), .I1 (g27573), .I2 (g21914));
AN2X1 gate18698(.O (g28319), .I1 (g27855), .I2 (g22246));
AN2X1 gate18699(.O (g28320), .I1 (g27854), .I2 (g20637));
AN2X1 gate18700(.O (g28322), .I1 (g27937), .I2 (g13868));
AN2X1 gate18701(.O (g28323), .I1 (g8580), .I2 (g27838));
AN2X1 gate18702(.O (g28324), .I1 (g27810), .I2 (g20659));
AN2X1 gate18703(.O (g28326), .I1 (g27865), .I2 (g22274));
AN2X1 gate18704(.O (g28327), .I1 (g27900), .I2 (g22275));
AN2X1 gate18705(.O (g28329), .I1 (g27823), .I2 (g20708));
AN2X1 gate18706(.O (g28330), .I1 (g27864), .I2 (g20711));
AN2X1 gate18707(.O (g28331), .I1 (g27802), .I2 (g22307));
AN2X1 gate18708(.O (g28332), .I1 (g27883), .I2 (g22331));
AN2X1 gate18709(.O (g28333), .I1 (g27882), .I2 (g20772));
AN2X1 gate18710(.O (g28334), .I1 (g27842), .I2 (g20793));
AN2X1 gate18711(.O (g28335), .I1 (g27814), .I2 (g22343));
AN2X1 gate18712(.O (g28336), .I1 (g27896), .I2 (g20810));
AN2X1 gate18713(.O (g28337), .I1 (g28002), .I2 (g19448));
AN2X1 gate18714(.O (g28338), .I1 (g28029), .I2 (g19475));
AN2X1 gate18715(.O (g28339), .I1 (g28059), .I2 (g19498));
AN2X1 gate18716(.O (g28340), .I1 (g28088), .I2 (g19519));
AN2X1 gate18717(.O (g28373), .I1 (g56), .I2 (g27969));
AN2X1 gate18718(.O (g28376), .I1 (g744), .I2 (g27990));
AN2X1 gate18719(.O (g28378), .I1 (g52), .I2 (g27776));
AN3X1 gate18720(.O (g28379), .I1 (g27868), .I2 (g19390), .I3 (g19369));
AN2X1 gate18721(.O (g28380), .I1 (g1430), .I2 (g28014));
AN2X1 gate18722(.O (g28381), .I1 (g28157), .I2 (g9815));
AN2X1 gate18723(.O (g28383), .I1 (g740), .I2 (g27780));
AN2X1 gate18724(.O (g28385), .I1 (g2124), .I2 (g28041));
AN2X1 gate18725(.O (g28387), .I1 (g1426), .I2 (g27787));
AN2X1 gate18726(.O (g28389), .I1 (g2120), .I2 (g27794));
AN2X1 gate18727(.O (g28396), .I1 (g7754), .I2 (g27806));
AN2X1 gate18728(.O (g28398), .I1 (g7769), .I2 (g27817));
AN2X1 gate18729(.O (g28399), .I1 (g7776), .I2 (g27820));
AN2X1 gate18730(.O (g28401), .I1 (g7782), .I2 (g27831));
AN2X1 gate18731(.O (g28402), .I1 (g7785), .I2 (g27839));
AN2X1 gate18732(.O (g28404), .I1 (g7792), .I2 (g27843));
AN2X1 gate18733(.O (g28405), .I1 (g7796), .I2 (g27847));
AN2X1 gate18734(.O (g28407), .I1 (g7799), .I2 (g27858));
AN2X1 gate18735(.O (g28408), .I1 (g7806), .I2 (g27861));
AN2X1 gate18736(.O (g28411), .I1 (g7809), .I2 (g27872));
AN2X1 gate18737(.O (g28412), .I1 (g7812), .I2 (g27879));
AN2X1 gate18738(.O (g28416), .I1 (g7823), .I2 (g27889));
AN2X1 gate18739(.O (g28422), .I1 (g17640), .I2 (g28150));
AN2X1 gate18740(.O (g28423), .I1 (g17724), .I2 (g28152));
AN2X1 gate18741(.O (g28424), .I1 (g17741), .I2 (g28153));
AN2X1 gate18742(.O (g28426), .I1 (g28128), .I2 (g9170));
AN2X1 gate18743(.O (g28427), .I1 (g26092), .I2 (g28154));
AN2X1 gate18744(.O (g28428), .I1 (g17825), .I2 (g28155));
AN2X1 gate18745(.O (g28429), .I1 (g17842), .I2 (g28156));
AN2X1 gate18746(.O (g28430), .I1 (g28128), .I2 (g9196));
AN2X1 gate18747(.O (g28431), .I1 (g26092), .I2 (g28158));
AN2X1 gate18748(.O (g28433), .I1 (g28133), .I2 (g9212));
AN2X1 gate18749(.O (g28434), .I1 (g26114), .I2 (g28159));
AN2X1 gate18750(.O (g28435), .I1 (g17937), .I2 (g28160));
AN2X1 gate18751(.O (g28436), .I1 (g17954), .I2 (g28161));
AN2X1 gate18752(.O (g28438), .I1 (g17882), .I2 (g27919));
AN2X1 gate18753(.O (g28439), .I1 (g28128), .I2 (g9242));
AN2X1 gate18754(.O (g28440), .I1 (g26092), .I2 (g28162));
AN2X1 gate18755(.O (g28441), .I1 (g28133), .I2 (g9257));
AN2X1 gate18756(.O (g28442), .I1 (g26114), .I2 (g28163));
AN2X1 gate18757(.O (g28444), .I1 (g28137), .I2 (g9273));
AN2X1 gate18758(.O (g28445), .I1 (g26121), .I2 (g28164));
AN2X1 gate18759(.O (g28446), .I1 (g18048), .I2 (g28165));
AN2X1 gate18760(.O (g28448), .I1 (g17974), .I2 (g27928));
AN2X1 gate18761(.O (g28450), .I1 (g17993), .I2 (g27932));
AN2X1 gate18762(.O (g28451), .I1 (g28133), .I2 (g9320));
AN2X1 gate18763(.O (g28452), .I1 (g26114), .I2 (g28166));
AN2X1 gate18764(.O (g28453), .I1 (g28137), .I2 (g9335));
AN2X1 gate18765(.O (g28454), .I1 (g26121), .I2 (g28167));
AN2X1 gate18766(.O (g28456), .I1 (g28141), .I2 (g9351));
AN2X1 gate18767(.O (g28457), .I1 (g26131), .I2 (g28168));
AN2X1 gate18768(.O (g28459), .I1 (g18074), .I2 (g27939));
AN2X1 gate18769(.O (g28460), .I1 (g18091), .I2 (g27942));
AN2X1 gate18770(.O (g28462), .I1 (g18110), .I2 (g27946));
AN2X1 gate18771(.O (g28463), .I1 (g28137), .I2 (g9401));
AN2X1 gate18772(.O (g28464), .I1 (g26121), .I2 (g28169));
AN2X1 gate18773(.O (g28465), .I1 (g28141), .I2 (g9416));
AN2X1 gate18774(.O (g28466), .I1 (g26131), .I2 (g28170));
AN2X1 gate18775(.O (g28468), .I1 (g18265), .I2 (g28172));
AN2X1 gate18776(.O (g28469), .I1 (g18179), .I2 (g27952));
AN2X1 gate18777(.O (g28471), .I1 (g18190), .I2 (g27956));
AN2X1 gate18778(.O (g28472), .I1 (g18207), .I2 (g27959));
AN2X1 gate18779(.O (g28474), .I1 (g18226), .I2 (g27965));
AN2X1 gate18780(.O (g28475), .I1 (g28141), .I2 (g9498));
AN2X1 gate18781(.O (g28476), .I1 (g26131), .I2 (g28173));
AN2X1 gate18782(.O (g28477), .I1 (g18341), .I2 (g28174));
AN2X1 gate18783(.O (g28478), .I1 (g18358), .I2 (g28175));
AN2X1 gate18784(.O (g28479), .I1 (g18286), .I2 (g27973));
AN2X1 gate18785(.O (g28480), .I1 (g18297), .I2 (g27977));
AN2X1 gate18786(.O (g28481), .I1 (g18314), .I2 (g27981));
AN2X1 gate18787(.O (g28484), .I1 (g18436), .I2 (g28177));
AN2X1 gate18788(.O (g28485), .I1 (g18453), .I2 (g28178));
AN2X1 gate18789(.O (g28486), .I1 (g18379), .I2 (g27994));
AN2X1 gate18790(.O (g28487), .I1 (g18390), .I2 (g27999));
AN2X1 gate18791(.O (g28492), .I1 (g18509), .I2 (g28186));
AN2X1 gate18792(.O (g28493), .I1 (g18526), .I2 (g28187));
AN2X1 gate18793(.O (g28494), .I1 (g18474), .I2 (g28018));
AN2X1 gate18794(.O (g28497), .I1 (g18573), .I2 (g28190));
AN2X1 gate18795(.O (g28657), .I1 (g27925), .I2 (g13700));
AN2X1 gate18796(.O (g28659), .I1 (g27917), .I2 (g13736));
AN2X1 gate18797(.O (g28660), .I1 (g27916), .I2 (g11911));
AN2X1 gate18798(.O (g28662), .I1 (g27911), .I2 (g11951));
AN2X1 gate18799(.O (g28663), .I1 (g27906), .I2 (g11997));
AN2X1 gate18800(.O (g28664), .I1 (g27997), .I2 (g12055));
AN2X1 gate18801(.O (g28665), .I1 (g27827), .I2 (g22222));
AN2X1 gate18802(.O (g28666), .I1 (g27980), .I2 (g12106));
AN2X1 gate18803(.O (g28667), .I1 (g27964), .I2 (g13852));
AN2X1 gate18804(.O (g28669), .I1 (g27897), .I2 (g22233));
AN2X1 gate18805(.O (g28670), .I1 (g27798), .I2 (g21935));
AN2X1 gate18806(.O (g28671), .I1 (g27962), .I2 (g12161));
AN2X1 gate18807(.O (g28672), .I1 (g27950), .I2 (g13859));
AN2X1 gate18808(.O (g28707), .I1 (g12436), .I2 (g28379));
AN2X1 gate18809(.O (g28708), .I1 (g28392), .I2 (g22260));
AN2X1 gate18810(.O (g28709), .I1 (g28400), .I2 (g22261));
AN2X1 gate18811(.O (g28710), .I1 (g28403), .I2 (g22262));
AN2X1 gate18812(.O (g28711), .I1 (g10749), .I2 (g28415));
AN2X1 gate18813(.O (g28712), .I1 (g28406), .I2 (g22276));
AN2X1 gate18814(.O (g28713), .I1 (g28410), .I2 (g22290));
AN2X1 gate18815(.O (g28714), .I1 (g28394), .I2 (g22306));
AN2X1 gate18816(.O (g28715), .I1 (g28414), .I2 (g22332));
AN2X1 gate18817(.O (g28716), .I1 (g28449), .I2 (g19319));
AN2X1 gate18818(.O (g28717), .I1 (g28461), .I2 (g19346));
AN2X1 gate18819(.O (g28718), .I1 (g28473), .I2 (g19380));
AN2X1 gate18820(.O (g28719), .I1 (g28482), .I2 (g19412));
AN2X1 gate18821(.O (g28722), .I1 (g28523), .I2 (g16694));
AN2X1 gate18822(.O (g28724), .I1 (g28551), .I2 (g16725));
AN2X1 gate18823(.O (g28726), .I1 (g28578), .I2 (g16767));
AN2X1 gate18824(.O (g28729), .I1 (g28606), .I2 (g16794));
AN2X1 gate18825(.O (g28834), .I1 (g5751), .I2 (g28483));
AN2X1 gate18826(.O (g28836), .I1 (g5810), .I2 (g28491));
AN2X1 gate18827(.O (g28838), .I1 (g5866), .I2 (g28496));
AN2X1 gate18828(.O (g28840), .I1 (g5913), .I2 (g28500));
AN2X1 gate18829(.O (g28841), .I1 (g27834), .I2 (g28554));
AN2X1 gate18830(.O (g28843), .I1 (g27834), .I2 (g28581));
AN2X1 gate18831(.O (g28844), .I1 (g27850), .I2 (g28582));
AN2X1 gate18832(.O (g28846), .I1 (g27834), .I2 (g28608));
AN2X1 gate18833(.O (g28847), .I1 (g27850), .I2 (g28609));
AN2X1 gate18834(.O (g28848), .I1 (g27875), .I2 (g28610));
AN2X1 gate18835(.O (g28849), .I1 (g27850), .I2 (g28616));
AN2X1 gate18836(.O (g28850), .I1 (g27875), .I2 (g28617));
AN2X1 gate18837(.O (g28851), .I1 (g27892), .I2 (g28618));
AN2X1 gate18838(.O (g28852), .I1 (g27875), .I2 (g28623));
AN2X1 gate18839(.O (g28853), .I1 (g27892), .I2 (g28624));
AN2X1 gate18840(.O (g28854), .I1 (g27892), .I2 (g28629));
AN2X1 gate18841(.O (g28880), .I1 (g13946), .I2 (g28639));
AN2X1 gate18842(.O (g28881), .I1 (g28612), .I2 (g9199));
AN2X1 gate18843(.O (g28892), .I1 (g14001), .I2 (g28640));
AN2X1 gate18844(.O (g28893), .I1 (g28612), .I2 (g9245));
AN2X1 gate18845(.O (g28897), .I1 (g14016), .I2 (g28641));
AN2X1 gate18846(.O (g28898), .I1 (g28619), .I2 (g9260));
AN2X1 gate18847(.O (g28909), .I1 (g14062), .I2 (g28642));
AN2X1 gate18848(.O (g28910), .I1 (g28612), .I2 (g9303));
AN2X1 gate18849(.O (g28914), .I1 (g14092), .I2 (g28643));
AN2X1 gate18850(.O (g28915), .I1 (g28619), .I2 (g9323));
AN2X1 gate18851(.O (g28919), .I1 (g14107), .I2 (g28644));
AN2X1 gate18852(.O (g28923), .I1 (g28625), .I2 (g9338));
AN2X1 gate18853(.O (g28931), .I1 (g14153), .I2 (g28645));
AN2X1 gate18854(.O (g28935), .I1 (g14177), .I2 (g28646));
AN2X1 gate18855(.O (g28936), .I1 (g28619), .I2 (g9384));
AN2X1 gate18856(.O (g28940), .I1 (g14207), .I2 (g28647));
AN2X1 gate18857(.O (g28944), .I1 (g28625), .I2 (g9404));
AN2X1 gate18858(.O (g28948), .I1 (g14222), .I2 (g28648));
AN2X1 gate18859(.O (g28949), .I1 (g28630), .I2 (g9419));
AN2X1 gate18860(.O (g28958), .I1 (g14268), .I2 (g28649));
AN2X1 gate18861(.O (g28962), .I1 (g14292), .I2 (g28650));
AN2X1 gate18862(.O (g28966), .I1 (g28625), .I2 (g9481));
AN2X1 gate18863(.O (g28970), .I1 (g14322), .I2 (g28651));
AN2X1 gate18864(.O (g28971), .I1 (g28630), .I2 (g9501));
AN2X1 gate18865(.O (g28986), .I1 (g14390), .I2 (g28652));
AN2X1 gate18866(.O (g28996), .I1 (g14414), .I2 (g28653));
AN2X1 gate18867(.O (g28997), .I1 (g28630), .I2 (g9623));
AN2X1 gate18868(.O (g29022), .I1 (g14502), .I2 (g28655));
AN2X1 gate18869(.O (g29130), .I1 (g28397), .I2 (g22221));
AN2X1 gate18870(.O (g29174), .I1 (g29031), .I2 (g20684));
AN2X1 gate18871(.O (g29175), .I1 (g29009), .I2 (g20687));
AN2X1 gate18872(.O (g29176), .I1 (g29097), .I2 (g20690));
AN2X1 gate18873(.O (g29180), .I1 (g28982), .I2 (g20714));
AN2X1 gate18874(.O (g29183), .I1 (g29064), .I2 (g20739));
AN2X1 gate18875(.O (g29186), .I1 (g29063), .I2 (g20769));
AN2X1 gate18876(.O (g29188), .I1 (g29083), .I2 (g20796));
AN2X1 gate18877(.O (g29196), .I1 (g15022), .I2 (g28741));
AN2X1 gate18878(.O (g29200), .I1 (g15096), .I2 (g28751));
AN2X1 gate18879(.O (g29203), .I1 (g15118), .I2 (g28755));
AN2X1 gate18880(.O (g29208), .I1 (g15188), .I2 (g28764));
AN2X1 gate18881(.O (g29211), .I1 (g15210), .I2 (g28768));
AN2X1 gate18882(.O (g29217), .I1 (g15274), .I2 (g28775));
AN2X1 gate18883(.O (g29220), .I1 (g15296), .I2 (g28779));
AN2X1 gate18884(.O (g29225), .I1 (g15366), .I2 (g28785));
AN2X1 gate18885(.O (g29229), .I1 (g9293), .I2 (g28791));
AN2X1 gate18886(.O (g29232), .I1 (g9356), .I2 (g28796));
AN2X1 gate18887(.O (g29233), .I1 (g9374), .I2 (g28799));
AN2X1 gate18888(.O (g29234), .I1 (g9427), .I2 (g28804));
AN2X1 gate18889(.O (g29235), .I1 (g9453), .I2 (g28807));
AN2X1 gate18890(.O (g29236), .I1 (g9471), .I2 (g28810));
AN2X1 gate18891(.O (g29238), .I1 (g9569), .I2 (g28814));
AN2X1 gate18892(.O (g29239), .I1 (g9595), .I2 (g28817));
AN2X1 gate18893(.O (g29240), .I1 (g9613), .I2 (g28820));
AN2X1 gate18894(.O (g29241), .I1 (g9711), .I2 (g28823));
AN2X1 gate18895(.O (g29242), .I1 (g9737), .I2 (g28826));
AN2X1 gate18896(.O (g29243), .I1 (g9857), .I2 (g28829));
AN2X1 gate18897(.O (g29248), .I1 (g28855), .I2 (g8836));
AN2X1 gate18898(.O (g29251), .I1 (g28855), .I2 (g8856));
AN2X1 gate18899(.O (g29252), .I1 (g28859), .I2 (g8863));
AN2X1 gate18900(.O (g29255), .I1 (g28855), .I2 (g8885));
AN2X1 gate18901(.O (g29256), .I1 (g28859), .I2 (g8894));
AN2X1 gate18902(.O (g29257), .I1 (g28863), .I2 (g8901));
AN2X1 gate18903(.O (g29259), .I1 (g28859), .I2 (g8925));
AN2X1 gate18904(.O (g29260), .I1 (g28863), .I2 (g8934));
AN2X1 gate18905(.O (g29261), .I1 (g28867), .I2 (g8941));
AN2X1 gate18906(.O (g29262), .I1 (g28863), .I2 (g8965));
AN2X1 gate18907(.O (g29263), .I1 (g28867), .I2 (g8974));
AN2X1 gate18908(.O (g29264), .I1 (g28867), .I2 (g8997));
AN2X1 gate18909(.O (g29284), .I1 (g29001), .I2 (g28871));
AN2X1 gate18910(.O (g29289), .I1 (g29030), .I2 (g28883));
AN2X1 gate18911(.O (g29294), .I1 (g29053), .I2 (g28900));
AN2X1 gate18912(.O (g29300), .I1 (g29072), .I2 (g28925));
AN2X1 gate18913(.O (g29302), .I1 (g29026), .I2 (g28928));
AN2X1 gate18914(.O (g29310), .I1 (g28978), .I2 (g28951));
AN2X1 gate18915(.O (g29312), .I1 (g29049), .I2 (g28955));
AN2X1 gate18916(.O (g29320), .I1 (g29088), .I2 (g28972));
AN2X1 gate18917(.O (g29321), .I1 (g29008), .I2 (g28979));
AN2X1 gate18918(.O (g29323), .I1 (g29068), .I2 (g28983));
AN2X1 gate18919(.O (g29329), .I1 (g29096), .I2 (g29002));
AN2X1 gate18920(.O (g29330), .I1 (g29038), .I2 (g29010));
AN2X1 gate18921(.O (g29332), .I1 (g29080), .I2 (g29019));
AN2X1 gate18922(.O (g29336), .I1 (g29045), .I2 (g29023));
AN2X1 gate18923(.O (g29337), .I1 (g29103), .I2 (g29032));
AN2X1 gate18924(.O (g29338), .I1 (g29060), .I2 (g29042));
AN2X1 gate18925(.O (g29341), .I1 (g29062), .I2 (g29046));
AN2X1 gate18926(.O (g29342), .I1 (g29107), .I2 (g29054));
AN2X1 gate18927(.O (g29344), .I1 (g29076), .I2 (g29065));
AN2X1 gate18928(.O (g29346), .I1 (g29087), .I2 (g29077));
AN2X1 gate18929(.O (g29411), .I1 (g29090), .I2 (g21932));
AN2X1 gate18930(.O (g29464), .I1 (g29190), .I2 (g8375));
AN2X1 gate18931(.O (g29465), .I1 (g29191), .I2 (g8424));
AN2X1 gate18932(.O (g29466), .I1 (g8587), .I2 (g29265));
AN2X1 gate18933(.O (g29467), .I1 (g29340), .I2 (g19467));
AN2X1 gate18934(.O (g29468), .I1 (g29343), .I2 (g19490));
AN2X1 gate18935(.O (g29469), .I1 (g29345), .I2 (g19511));
AN2X1 gate18936(.O (g29470), .I1 (g29347), .I2 (g19530));
AN2X1 gate18937(.O (g29471), .I1 (g21461), .I2 (g29266));
AN2X1 gate18938(.O (g29472), .I1 (g21461), .I2 (g29268));
AN2X1 gate18939(.O (g29473), .I1 (g21508), .I2 (g29269));
AN2X1 gate18940(.O (g29474), .I1 (g21508), .I2 (g29271));
AN2X1 gate18941(.O (g29475), .I1 (g21544), .I2 (g29272));
AN2X1 gate18942(.O (g29476), .I1 (g21544), .I2 (g29274));
AN2X1 gate18943(.O (g29477), .I1 (g21580), .I2 (g29275));
AN2X1 gate18944(.O (g29478), .I1 (g21580), .I2 (g29277));
AN2X1 gate18945(.O (g29479), .I1 (g21461), .I2 (g29280));
AN2X1 gate18946(.O (g29480), .I1 (g21461), .I2 (g29282));
AN2X1 gate18947(.O (g29481), .I1 (g21508), .I2 (g29283));
AN2X1 gate18948(.O (g29482), .I1 (g21461), .I2 (g29285));
AN2X1 gate18949(.O (g29483), .I1 (g21508), .I2 (g29286));
AN2X1 gate18950(.O (g29484), .I1 (g21544), .I2 (g29287));
AN2X1 gate18951(.O (g29485), .I1 (g21508), .I2 (g29290));
AN2X1 gate18952(.O (g29486), .I1 (g21544), .I2 (g29291));
AN2X1 gate18953(.O (g29487), .I1 (g21580), .I2 (g29292));
AN2X1 gate18954(.O (g29488), .I1 (g21544), .I2 (g29295));
AN2X1 gate18955(.O (g29489), .I1 (g21580), .I2 (g29296));
AN2X1 gate18956(.O (g29490), .I1 (g21580), .I2 (g29301));
AN2X1 gate18957(.O (g29502), .I1 (g29350), .I2 (g8912));
AN2X1 gate18958(.O (g29518), .I1 (g28728), .I2 (g29360));
AN2X1 gate18959(.O (g29520), .I1 (g28731), .I2 (g29361));
AN2X1 gate18960(.O (g29521), .I1 (g28733), .I2 (g29362));
AN2X1 gate18961(.O (g29522), .I1 (g27735), .I2 (g29363));
AN2X1 gate18962(.O (g29523), .I1 (g28737), .I2 (g29364));
AN2X1 gate18963(.O (g29524), .I1 (g28739), .I2 (g29365));
AN2X1 gate18964(.O (g29525), .I1 (g29195), .I2 (g29366));
AN2X1 gate18965(.O (g29526), .I1 (g27741), .I2 (g29367));
AN2X1 gate18966(.O (g29527), .I1 (g28748), .I2 (g29368));
AN2X1 gate18967(.O (g29528), .I1 (g28750), .I2 (g29369));
AN2X1 gate18968(.O (g29529), .I1 (g29199), .I2 (g29370));
AN2X1 gate18969(.O (g29531), .I1 (g29202), .I2 (g29371));
AN2X1 gate18970(.O (g29532), .I1 (g27746), .I2 (g29372));
AN2X1 gate18971(.O (g29533), .I1 (g28762), .I2 (g29373));
AN2X1 gate18972(.O (g29534), .I1 (g29206), .I2 (g29374));
AN2X1 gate18973(.O (g29536), .I1 (g29207), .I2 (g29375));
AN2X1 gate18974(.O (g29538), .I1 (g29210), .I2 (g29376));
AN2X1 gate18975(.O (g29539), .I1 (g27754), .I2 (g29377));
AN2X1 gate18976(.O (g29540), .I1 (g26041), .I2 (g29378));
AN2X1 gate18977(.O (g29541), .I1 (g29214), .I2 (g29379));
AN2X1 gate18978(.O (g29543), .I1 (g29215), .I2 (g29380));
AN2X1 gate18979(.O (g29545), .I1 (g29216), .I2 (g29381));
AN2X1 gate18980(.O (g29547), .I1 (g29219), .I2 (g29382));
AN2X1 gate18981(.O (g29548), .I1 (g28784), .I2 (g29383));
AN2X1 gate18982(.O (g29549), .I1 (g26043), .I2 (g29384));
AN2X1 gate18983(.O (g29550), .I1 (g29222), .I2 (g29385));
AN2X1 gate18984(.O (g29553), .I1 (g29223), .I2 (g29386));
AN2X1 gate18985(.O (g29555), .I1 (g29224), .I2 (g29387));
AN2X1 gate18986(.O (g29557), .I1 (g28789), .I2 (g29388));
AN2X1 gate18987(.O (g29558), .I1 (g28790), .I2 (g29389));
AN2X1 gate18988(.O (g29559), .I1 (g26045), .I2 (g29390));
AN2X1 gate18989(.O (g29560), .I1 (g29227), .I2 (g29391));
AN2X1 gate18990(.O (g29562), .I1 (g29228), .I2 (g29392));
AN2X1 gate18991(.O (g29564), .I1 (g28794), .I2 (g29393));
AN2X1 gate18992(.O (g29565), .I1 (g28795), .I2 (g29394));
AN2X1 gate18993(.O (g29566), .I1 (g26047), .I2 (g29395));
AN2X1 gate18994(.O (g29567), .I1 (g29231), .I2 (g29396));
AN2X1 gate18995(.O (g29572), .I1 (g28802), .I2 (g29397));
AN2X1 gate18996(.O (g29573), .I1 (g28803), .I2 (g29398));
AN2X1 gate18997(.O (g29575), .I1 (g28813), .I2 (g29402));
AN2X1 gate18998(.O (g29607), .I1 (g29193), .I2 (g11056));
AN2X1 gate18999(.O (g29610), .I1 (g29349), .I2 (g11123));
AN2X1 gate19000(.O (g29614), .I1 (g29359), .I2 (g11182));
AN2X1 gate19001(.O (g29615), .I1 (g29245), .I2 (g11185));
AN2X1 gate19002(.O (g29619), .I1 (g29247), .I2 (g11259));
AN2X1 gate19003(.O (g29622), .I1 (g29250), .I2 (g11327));
AN2X1 gate19004(.O (g29624), .I1 (g29254), .I2 (g11407));
AN2X1 gate19005(.O (g29625), .I1 (g29189), .I2 (g11472));
AN2X1 gate19006(.O (g29626), .I1 (g29318), .I2 (g11478));
AN2X1 gate19007(.O (g29790), .I1 (g29491), .I2 (g10918));
AN2X1 gate19008(.O (g29792), .I1 (g29491), .I2 (g10977));
AN2X1 gate19009(.O (g29793), .I1 (g29491), .I2 (g11063));
AN2X1 gate19010(.O (g29810), .I1 (g29748), .I2 (g22248));
AN2X1 gate19011(.O (g29811), .I1 (g29703), .I2 (g20644));
AN2X1 gate19012(.O (g29812), .I1 (g29762), .I2 (g12223));
AN2X1 gate19013(.O (g29813), .I1 (g29760), .I2 (g13869));
AN2X1 gate19014(.O (g29814), .I1 (g29728), .I2 (g22266));
AN2X1 gate19015(.O (g29815), .I1 (g29727), .I2 (g20662));
AN2X1 gate19016(.O (g29816), .I1 (g29759), .I2 (g13883));
AN2X1 gate19017(.O (g29817), .I1 (g29709), .I2 (g20694));
AN2X1 gate19018(.O (g29818), .I1 (g29732), .I2 (g22293));
AN2X1 gate19019(.O (g29819), .I1 (g29751), .I2 (g22294));
AN2X1 gate19020(.O (g29820), .I1 (g29717), .I2 (g20743));
AN2X1 gate19021(.O (g29821), .I1 (g29731), .I2 (g20746));
AN2X1 gate19022(.O (g29822), .I1 (g29705), .I2 (g22335));
AN2X1 gate19023(.O (g29827), .I1 (g29741), .I2 (g22356));
AN2X1 gate19024(.O (g29828), .I1 (g29740), .I2 (g20802));
AN2X1 gate19025(.O (g29833), .I1 (g29725), .I2 (g20813));
AN2X1 gate19026(.O (g29834), .I1 (g29713), .I2 (g22366));
AN2X1 gate19027(.O (g29839), .I1 (g29747), .I2 (g20827));
AN3X1 gate19028(.O (g29909), .I1 (g29735), .I2 (g19420), .I3 (g19401));
AN2X1 gate19029(.O (g29910), .I1 (g29779), .I2 (g9961));
AN2X1 gate19030(.O (g29942), .I1 (g29771), .I2 (g28877));
AN2X1 gate19031(.O (g29944), .I1 (g29782), .I2 (g28889));
AN2X1 gate19032(.O (g29945), .I1 (g29773), .I2 (g28894));
AN2X1 gate19033(.O (g29946), .I1 (g29778), .I2 (g28906));
AN2X1 gate19034(.O (g29947), .I1 (g29785), .I2 (g28911));
AN2X1 gate19035(.O (g29948), .I1 (g29775), .I2 (g28916));
AN2X1 gate19036(.O (g29949), .I1 (g29781), .I2 (g28932));
AN2X1 gate19037(.O (g29950), .I1 (g29788), .I2 (g28937));
AN2X1 gate19038(.O (g29951), .I1 (g29777), .I2 (g28945));
AN2X1 gate19039(.O (g29952), .I1 (g29784), .I2 (g28959));
AN2X1 gate19040(.O (g29953), .I1 (g29791), .I2 (g28967));
AN2X1 gate19041(.O (g29954), .I1 (g29770), .I2 (g28975));
AN2X1 gate19042(.O (g29955), .I1 (g29787), .I2 (g28993));
AN2X1 gate19043(.O (g29956), .I1 (g29780), .I2 (g28998));
AN2X1 gate19044(.O (g29957), .I1 (g29772), .I2 (g29005));
AN2X1 gate19045(.O (g29958), .I1 (g29783), .I2 (g29027));
AN2X1 gate19046(.O (g29959), .I1 (g29774), .I2 (g29035));
AN2X1 gate19047(.O (g29960), .I1 (g29786), .I2 (g29050));
AN2X1 gate19048(.O (g29961), .I1 (g29776), .I2 (g29057));
AN2X1 gate19049(.O (g29962), .I1 (g29789), .I2 (g29069));
AN2X1 gate19050(.O (g29963), .I1 (g29758), .I2 (g13737));
AN2X1 gate19051(.O (g29964), .I1 (g29757), .I2 (g13786));
AN2X1 gate19052(.O (g29965), .I1 (g29756), .I2 (g11961));
AN2X1 gate19053(.O (g29966), .I1 (g29755), .I2 (g12004));
AN2X1 gate19054(.O (g29967), .I1 (g29754), .I2 (g12066));
AN2X1 gate19055(.O (g29968), .I1 (g29765), .I2 (g12119));
AN2X1 gate19056(.O (g29969), .I1 (g29721), .I2 (g22237));
AN2X1 gate19057(.O (g29970), .I1 (g29764), .I2 (g12178));
AN2X1 gate19058(.O (g29971), .I1 (g29763), .I2 (g13861));
AN2X1 gate19059(.O (g29980), .I1 (g29881), .I2 (g8324));
AN2X1 gate19060(.O (g29981), .I1 (g29869), .I2 (g8330));
AN2X1 gate19061(.O (g29982), .I1 (g29893), .I2 (g8336));
AN2X1 gate19062(.O (g29983), .I1 (g29885), .I2 (g8344));
AN2X1 gate19063(.O (g29984), .I1 (g29873), .I2 (g8351));
AN2X1 gate19064(.O (g29985), .I1 (g29897), .I2 (g8363));
AN2X1 gate19065(.O (g29986), .I1 (g29877), .I2 (g8366));
AN2X1 gate19066(.O (g29987), .I1 (g29889), .I2 (g8369));
AN2X1 gate19067(.O (g29988), .I1 (g29881), .I2 (g8382));
AN2X1 gate19068(.O (g29989), .I1 (g29893), .I2 (g8391));
AN2X1 gate19069(.O (g29990), .I1 (g29885), .I2 (g8397));
AN2X1 gate19070(.O (g29991), .I1 (g29901), .I2 (g8403));
AN2X1 gate19071(.O (g29992), .I1 (g12441), .I2 (g29909));
AN2X1 gate19072(.O (g29993), .I1 (g29897), .I2 (g8411));
AN2X1 gate19073(.O (g29994), .I1 (g29889), .I2 (g8418));
AN2X1 gate19074(.O (g29995), .I1 (g29893), .I2 (g8434));
AN2X1 gate19075(.O (g29996), .I1 (g29901), .I2 (g8443));
AN2X1 gate19076(.O (g29997), .I1 (g29918), .I2 (g22277));
AN2X1 gate19077(.O (g29998), .I1 (g29922), .I2 (g22278));
AN2X1 gate19078(.O (g29999), .I1 (g29924), .I2 (g22279));
AN2X1 gate19079(.O (g30000), .I1 (g10767), .I2 (g29930));
AN2X1 gate19080(.O (g30001), .I1 (g29897), .I2 (g8449));
AN2X1 gate19081(.O (g30002), .I1 (g29905), .I2 (g8455));
AN2X1 gate19082(.O (g30003), .I1 (g29901), .I2 (g8469));
AN2X1 gate19083(.O (g30004), .I1 (g29926), .I2 (g22295));
AN2X1 gate19084(.O (g30005), .I1 (g29905), .I2 (g8478));
AN2X1 gate19085(.O (g30006), .I1 (g29928), .I2 (g22310));
AN2X1 gate19086(.O (g30007), .I1 (g29905), .I2 (g8494));
AN2X1 gate19087(.O (g30008), .I1 (g29919), .I2 (g22334));
AN2X1 gate19088(.O (g30009), .I1 (g29929), .I2 (g22357));
AN2X1 gate19089(.O (g30077), .I1 (g29823), .I2 (g10963));
AN2X1 gate19090(.O (g30079), .I1 (g29823), .I2 (g10988));
AN2X1 gate19091(.O (g30080), .I1 (g29829), .I2 (g10996));
AN2X1 gate19092(.O (g30081), .I1 (g29823), .I2 (g11022));
AN2X1 gate19093(.O (g30082), .I1 (g29829), .I2 (g11036));
AN2X1 gate19094(.O (g30083), .I1 (g29835), .I2 (g11048));
AN2X1 gate19095(.O (g30085), .I1 (g29829), .I2 (g11092));
AN2X1 gate19096(.O (g30086), .I1 (g29835), .I2 (g11108));
AN2X1 gate19097(.O (g30087), .I1 (g29840), .I2 (g11120));
AN2X1 gate19098(.O (g30088), .I1 (g29844), .I2 (g11138));
AN2X1 gate19099(.O (g30089), .I1 (g29835), .I2 (g11160));
AN2X1 gate19100(.O (g30090), .I1 (g29840), .I2 (g11176));
AN2X1 gate19101(.O (g30091), .I1 (g29844), .I2 (g11202));
AN2X1 gate19102(.O (g30092), .I1 (g29849), .I2 (g11205));
AN2X1 gate19103(.O (g30093), .I1 (g29853), .I2 (g11222));
AN2X1 gate19104(.O (g30094), .I1 (g29840), .I2 (g11246));
AN2X1 gate19105(.O (g30095), .I1 (g29857), .I2 (g11265));
AN2X1 gate19106(.O (g30096), .I1 (g29844), .I2 (g11268));
AN2X1 gate19107(.O (g30097), .I1 (g29849), .I2 (g11271));
AN2X1 gate19108(.O (g30098), .I1 (g29853), .I2 (g11284));
AN2X1 gate19109(.O (g30099), .I1 (g29861), .I2 (g11287));
AN2X1 gate19110(.O (g30100), .I1 (g29865), .I2 (g11306));
AN2X1 gate19111(.O (g30101), .I1 (g29857), .I2 (g11341));
AN2X1 gate19112(.O (g30102), .I1 (g29849), .I2 (g11348));
AN2X1 gate19113(.O (g30103), .I1 (g29869), .I2 (g11358));
AN2X1 gate19114(.O (g30104), .I1 (g29853), .I2 (g11361));
AN2X1 gate19115(.O (g30105), .I1 (g29861), .I2 (g11364));
AN2X1 gate19116(.O (g30106), .I1 (g29865), .I2 (g11379));
AN2X1 gate19117(.O (g30107), .I1 (g29873), .I2 (g11382));
AN2X1 gate19118(.O (g30108), .I1 (g29877), .I2 (g11401));
AN2X1 gate19119(.O (g30109), .I1 (g29857), .I2 (g11411));
AN2X1 gate19120(.O (g30110), .I1 (g29881), .I2 (g11417));
AN2X1 gate19121(.O (g30111), .I1 (g29869), .I2 (g11425));
AN2X1 gate19122(.O (g30112), .I1 (g29861), .I2 (g11432));
AN2X1 gate19123(.O (g30113), .I1 (g29885), .I2 (g11444));
AN2X1 gate19124(.O (g30114), .I1 (g29865), .I2 (g11447));
AN2X1 gate19125(.O (g30115), .I1 (g29873), .I2 (g11450));
AN2X1 gate19126(.O (g30116), .I1 (g29921), .I2 (g22236));
AN2X1 gate19127(.O (g30117), .I1 (g29877), .I2 (g11465));
AN2X1 gate19128(.O (g30118), .I1 (g29889), .I2 (g11468));
AN2X1 gate19129(.O (g30123), .I1 (g30070), .I2 (g20641));
AN2X1 gate19130(.O (g30127), .I1 (g30065), .I2 (g20719));
AN2X1 gate19131(.O (g30128), .I1 (g30062), .I2 (g20722));
AN2X1 gate19132(.O (g30129), .I1 (g30071), .I2 (g20725));
AN2X1 gate19133(.O (g30131), .I1 (g30059), .I2 (g20749));
AN2X1 gate19134(.O (g30132), .I1 (g30068), .I2 (g20776));
AN2X1 gate19135(.O (g30133), .I1 (g30067), .I2 (g20799));
AN2X1 gate19136(.O (g30138), .I1 (g30069), .I2 (g20816));
AN2X1 gate19137(.O (g30216), .I1 (g30036), .I2 (g8921));
AN2X1 gate19138(.O (g30217), .I1 (g30036), .I2 (g8955));
AN2X1 gate19139(.O (g30218), .I1 (g30040), .I2 (g8961));
AN2X1 gate19140(.O (g30219), .I1 (g30036), .I2 (g8980));
AN2X1 gate19141(.O (g30220), .I1 (g30040), .I2 (g8987));
AN2X1 gate19142(.O (g30221), .I1 (g30044), .I2 (g8993));
AN2X1 gate19143(.O (g30222), .I1 (g30040), .I2 (g9010));
AN2X1 gate19144(.O (g30223), .I1 (g30044), .I2 (g9016));
AN2X1 gate19145(.O (g30224), .I1 (g30048), .I2 (g9022));
AN2X1 gate19146(.O (g30225), .I1 (g30044), .I2 (g9035));
AN2X1 gate19147(.O (g30226), .I1 (g30048), .I2 (g9041));
AN2X1 gate19148(.O (g30227), .I1 (g30048), .I2 (g9058));
AN2X1 gate19149(.O (g30327), .I1 (g30187), .I2 (g8321));
AN2X1 gate19150(.O (g30330), .I1 (g30195), .I2 (g8333));
AN2X1 gate19151(.O (g30333), .I1 (g30191), .I2 (g8341));
AN2X1 gate19152(.O (g30334), .I1 (g30203), .I2 (g8347));
AN2X1 gate19153(.O (g30337), .I1 (g30199), .I2 (g8354));
AN2X1 gate19154(.O (g30340), .I1 (g30207), .I2 (g8372));
AN2X1 gate19155(.O (g30345), .I1 (g30195), .I2 (g8388));
AN2X1 gate19156(.O (g30348), .I1 (g30203), .I2 (g8400));
AN2X1 gate19157(.O (g30351), .I1 (g30199), .I2 (g8408));
AN2X1 gate19158(.O (g30352), .I1 (g30211), .I2 (g8414));
AN2X1 gate19159(.O (g30355), .I1 (g30207), .I2 (g8421));
AN2X1 gate19160(.O (g30361), .I1 (g30203), .I2 (g8440));
AN2X1 gate19161(.O (g30364), .I1 (g30211), .I2 (g8452));
AN2X1 gate19162(.O (g30367), .I1 (g30207), .I2 (g8460));
AN2X1 gate19163(.O (g30372), .I1 (g8594), .I2 (g30228));
AN2X1 gate19164(.O (g30374), .I1 (g30211), .I2 (g8475));
AN2X1 gate19165(.O (g30387), .I1 (g30229), .I2 (g8888));
AN2X1 gate19166(.O (g30388), .I1 (g30229), .I2 (g8918));
AN2X1 gate19167(.O (g30389), .I1 (g30233), .I2 (g8928));
AN2X1 gate19168(.O (g30390), .I1 (g30229), .I2 (g8952));
AN2X1 gate19169(.O (g30391), .I1 (g30233), .I2 (g8958));
AN2X1 gate19170(.O (g30392), .I1 (g30237), .I2 (g8968));
AN2X1 gate19171(.O (g30393), .I1 (g30233), .I2 (g8984));
AN2X1 gate19172(.O (g30394), .I1 (g30237), .I2 (g8990));
AN2X1 gate19173(.O (g30395), .I1 (g30241), .I2 (g9000));
AN2X1 gate19174(.O (g30396), .I1 (g30237), .I2 (g9013));
AN2X1 gate19175(.O (g30397), .I1 (g30241), .I2 (g9019));
AN2X1 gate19176(.O (g30398), .I1 (g30241), .I2 (g9038));
AN2X1 gate19177(.O (g30407), .I1 (g30134), .I2 (g10991));
AN2X1 gate19178(.O (g30409), .I1 (g30134), .I2 (g11025));
AN2X1 gate19179(.O (g30410), .I1 (g30139), .I2 (g11028));
AN2X1 gate19180(.O (g30411), .I1 (g30143), .I2 (g11039));
AN2X1 gate19181(.O (g30436), .I1 (g30134), .I2 (g11079));
AN2X1 gate19182(.O (g30437), .I1 (g30139), .I2 (g11082));
AN2X1 gate19183(.O (g30438), .I1 (g30147), .I2 (g11085));
AN2X1 gate19184(.O (g30440), .I1 (g30143), .I2 (g11095));
AN2X1 gate19185(.O (g30441), .I1 (g30151), .I2 (g11098));
AN2X1 gate19186(.O (g30442), .I1 (g30155), .I2 (g11111));
AN2X1 gate19187(.O (g30444), .I1 (g30139), .I2 (g11132));
AN2X1 gate19188(.O (g30445), .I1 (g30147), .I2 (g11135));
AN2X1 gate19189(.O (g30447), .I1 (g30143), .I2 (g11145));
AN2X1 gate19190(.O (g30448), .I1 (g30151), .I2 (g11148));
AN2X1 gate19191(.O (g30449), .I1 (g30159), .I2 (g11151));
AN2X1 gate19192(.O (g30451), .I1 (g30155), .I2 (g11163));
AN2X1 gate19193(.O (g30452), .I1 (g30163), .I2 (g11166));
AN2X1 gate19194(.O (g30453), .I1 (g30167), .I2 (g11179));
AN2X1 gate19195(.O (g30454), .I1 (g30147), .I2 (g11199));
AN2X1 gate19196(.O (g30457), .I1 (g30151), .I2 (g11216));
AN2X1 gate19197(.O (g30458), .I1 (g30159), .I2 (g11219));
AN2X1 gate19198(.O (g30460), .I1 (g30155), .I2 (g11231));
AN2X1 gate19199(.O (g30461), .I1 (g30163), .I2 (g11234));
AN2X1 gate19200(.O (g30462), .I1 (g30171), .I2 (g11237));
AN2X1 gate19201(.O (g30464), .I1 (g30167), .I2 (g11249));
AN2X1 gate19202(.O (g30465), .I1 (g30175), .I2 (g11252));
AN2X1 gate19203(.O (g30467), .I1 (g30179), .I2 (g11274));
AN2X1 gate19204(.O (g30469), .I1 (g30159), .I2 (g11281));
AN2X1 gate19205(.O (g30472), .I1 (g30163), .I2 (g11300));
AN2X1 gate19206(.O (g30473), .I1 (g30171), .I2 (g11303));
AN2X1 gate19207(.O (g30475), .I1 (g30167), .I2 (g11315));
AN2X1 gate19208(.O (g30476), .I1 (g30175), .I2 (g11318));
AN2X1 gate19209(.O (g30477), .I1 (g30183), .I2 (g11321));
AN2X1 gate19210(.O (g30478), .I1 (g30187), .I2 (g11344));
AN2X1 gate19211(.O (g30481), .I1 (g30179), .I2 (g11351));
AN2X1 gate19212(.O (g30484), .I1 (g30191), .I2 (g11367));
AN2X1 gate19213(.O (g30486), .I1 (g30171), .I2 (g11376));
AN2X1 gate19214(.O (g30489), .I1 (g30175), .I2 (g11395));
AN2X1 gate19215(.O (g30490), .I1 (g30183), .I2 (g11398));
AN2X1 gate19216(.O (g30492), .I1 (g30187), .I2 (g11414));
AN2X1 gate19217(.O (g30495), .I1 (g30179), .I2 (g11422));
AN2X1 gate19218(.O (g30496), .I1 (g30195), .I2 (g11428));
AN2X1 gate19219(.O (g30499), .I1 (g30191), .I2 (g11435));
AN2X1 gate19220(.O (g30502), .I1 (g30199), .I2 (g11453));
AN2X1 gate19221(.O (g30504), .I1 (g30183), .I2 (g11462));
AN2X1 gate19222(.O (g30696), .I1 (g30383), .I2 (g10943));
AN2X1 gate19223(.O (g30697), .I1 (g30383), .I2 (g11011));
AN2X1 gate19224(.O (g30698), .I1 (g30383), .I2 (g11126));
AN2X1 gate19225(.O (g30728), .I1 (g30605), .I2 (g22252));
AN2X1 gate19226(.O (g30735), .I1 (g30629), .I2 (g22268));
AN2X1 gate19227(.O (g30736), .I1 (g30584), .I2 (g20669));
AN2X1 gate19228(.O (g30743), .I1 (g30610), .I2 (g22283));
AN2X1 gate19229(.O (g30744), .I1 (g30609), .I2 (g20697));
AN2X1 gate19230(.O (g30750), .I1 (g30593), .I2 (g20729));
AN2X1 gate19231(.O (g30754), .I1 (g30614), .I2 (g22313));
AN2X1 gate19232(.O (g30755), .I1 (g30632), .I2 (g22314));
AN2X1 gate19233(.O (g30757), .I1 (g30601), .I2 (g20780));
AN2X1 gate19234(.O (g30758), .I1 (g30613), .I2 (g20783));
AN2X1 gate19235(.O (g30759), .I1 (g30588), .I2 (g22360));
AN2X1 gate19236(.O (g30760), .I1 (g30622), .I2 (g22379));
AN2X1 gate19237(.O (g30761), .I1 (g30621), .I2 (g20822));
AN2X1 gate19238(.O (g30762), .I1 (g30608), .I2 (g20830));
AN2X1 gate19239(.O (g30763), .I1 (g30597), .I2 (g22386));
AN2X1 gate19240(.O (g30764), .I1 (g30628), .I2 (g20837));
AN3X1 gate19241(.O (g30766), .I1 (g30617), .I2 (g19457), .I3 (g19431));
AN2X1 gate19242(.O (g30916), .I1 (g30785), .I2 (g22251));
AN2X1 gate19243(.O (g30917), .I1 (g12446), .I2 (g30766));
AN2X1 gate19244(.O (g30918), .I1 (g30780), .I2 (g22296));
AN2X1 gate19245(.O (g30919), .I1 (g30786), .I2 (g22297));
AN2X1 gate19246(.O (g30920), .I1 (g30787), .I2 (g22298));
AN2X1 gate19247(.O (g30921), .I1 (g10773), .I2 (g30791));
AN2X1 gate19248(.O (g30922), .I1 (g30788), .I2 (g22315));
AN2X1 gate19249(.O (g30923), .I1 (g30789), .I2 (g22338));
AN2X1 gate19250(.O (g30924), .I1 (g30783), .I2 (g22359));
AN2X1 gate19251(.O (g30925), .I1 (g30790), .I2 (g22380));
AN2X1 gate19252(.O (g30944), .I1 (g30935), .I2 (g20666));
AN2X1 gate19253(.O (g30945), .I1 (g30931), .I2 (g20754));
AN2X1 gate19254(.O (g30946), .I1 (g30930), .I2 (g20757));
AN2X1 gate19255(.O (g30947), .I1 (g30936), .I2 (g20760));
AN2X1 gate19256(.O (g30948), .I1 (g30929), .I2 (g20786));
AN2X1 gate19257(.O (g30949), .I1 (g30933), .I2 (g20806));
AN2X1 gate19258(.O (g30950), .I1 (g30932), .I2 (g20819));
AN2X1 gate19259(.O (g30951), .I1 (g30934), .I2 (g20833));
AN2X1 gate19260(.O (g30953), .I1 (g8605), .I2 (g30952));
OR2X1 gate19261(.O (g9144), .I1 (g2986), .I2 (g5389));
OR2X1 gate19262(.O (g10778), .I1 (g2929), .I2 (g8022));
OR2X1 gate19263(.O (g12377), .I1 (g7553), .I2 (g11059));
OR2X1 gate19264(.O (g12407), .I1 (g7573), .I2 (g10779));
OR2X1 gate19265(.O (g12886), .I1 (g9534), .I2 (g3398));
OR2X1 gate19266(.O (g12926), .I1 (g9676), .I2 (g3554));
OR2X1 gate19267(.O (g12955), .I1 (g9822), .I2 (g3710));
OR2X1 gate19268(.O (g12984), .I1 (g9968), .I2 (g3866));
OR2X1 gate19269(.O (g16539), .I1 (g15880), .I2 (g14657));
OR2X1 gate19270(.O (g16571), .I1 (g15913), .I2 (g14691));
OR2X1 gate19271(.O (g16595), .I1 (g15942), .I2 (g14725));
OR2X1 gate19272(.O (g16615), .I1 (g15971), .I2 (g14753));
OR2X1 gate19273(.O (g17973), .I1 (g11623), .I2 (g15659));
OR2X1 gate19274(.O (g19181), .I1 (g17729), .I2 (g17979));
OR2X1 gate19275(.O (g19186), .I1 (g18419), .I2 (g17887));
OR2X1 gate19276(.O (g19187), .I1 (g18419), .I2 (g17729));
OR2X1 gate19277(.O (g19188), .I1 (g17830), .I2 (g18096));
OR2X1 gate19278(.O (g19191), .I1 (g17807), .I2 (g17887));
OR2X1 gate19279(.O (g19192), .I1 (g18183), .I2 (g18270));
OR2X1 gate19280(.O (g19193), .I1 (g18492), .I2 (g17998));
OR2X1 gate19281(.O (g19194), .I1 (g18492), .I2 (g17830));
OR2X1 gate19282(.O (g19195), .I1 (g17942), .I2 (g18212));
OR2X1 gate19283(.O (g19200), .I1 (g18346), .I2 (g18424));
OR2X1 gate19284(.O (g19201), .I1 (g18183), .I2 (g18424));
OR2X1 gate19285(.O (g19202), .I1 (g17919), .I2 (g17998));
OR2X1 gate19286(.O (g19203), .I1 (g18290), .I2 (g18363));
OR2X1 gate19287(.O (g19204), .I1 (g18556), .I2 (g18115));
OR2X1 gate19288(.O (g19205), .I1 (g18556), .I2 (g17942));
OR2X1 gate19289(.O (g19206), .I1 (g18053), .I2 (g18319));
OR2X1 gate19290(.O (g19209), .I1 (g18079), .I2 (g18346));
OR2X1 gate19291(.O (g19210), .I1 (g18079), .I2 (g18183));
OR2X1 gate19292(.O (g19211), .I1 (g18441), .I2 (g18497));
OR2X1 gate19293(.O (g19212), .I1 (g18290), .I2 (g18497));
OR2X1 gate19294(.O (g19213), .I1 (g18030), .I2 (g18115));
OR2X1 gate19295(.O (g19214), .I1 (g18383), .I2 (g18458));
OR2X1 gate19296(.O (g19215), .I1 (g18606), .I2 (g18231));
OR2X1 gate19297(.O (g19216), .I1 (g18606), .I2 (g18053));
OR2X1 gate19298(.O (g19221), .I1 (g18270), .I2 (g18346));
OR2X1 gate19299(.O (g19222), .I1 (g18195), .I2 (g18441));
OR2X1 gate19300(.O (g19223), .I1 (g18195), .I2 (g18290));
OR2X1 gate19301(.O (g19224), .I1 (g18514), .I2 (g18561));
OR2X1 gate19302(.O (g19225), .I1 (g18383), .I2 (g18561));
OR2X1 gate19303(.O (g19226), .I1 (g18147), .I2 (g18231));
OR2X1 gate19304(.O (g19227), .I1 (g18478), .I2 (g18531));
OR3X1 gate19305(.O (I25477), .I1 (g17024), .I2 (g17000), .I3 (g16992));
OR3X1 gate19306(.O (g19230), .I1 (g16985), .I2 (g16965), .I3 (I25477));
OR2X1 gate19307(.O (g19231), .I1 (g18363), .I2 (g18441));
OR2X1 gate19308(.O (g19232), .I1 (g18302), .I2 (g18514));
OR2X1 gate19309(.O (g19233), .I1 (g18302), .I2 (g18383));
OR2X1 gate19310(.O (g19234), .I1 (g18578), .I2 (g18611));
OR2X1 gate19311(.O (g19235), .I1 (g18478), .I2 (g18611));
OR3X1 gate19312(.O (I25495), .I1 (g17158), .I2 (g17137), .I3 (g17115));
OR3X1 gate19313(.O (g19240), .I1 (g17083), .I2 (g17050), .I3 (I25495));
OR2X1 gate19314(.O (g19242), .I1 (g14244), .I2 (g16501));
OR3X1 gate19315(.O (I25500), .I1 (g17058), .I2 (g17030), .I3 (g17016));
OR3X1 gate19316(.O (g19243), .I1 (g16995), .I2 (g16986), .I3 (I25500));
OR2X1 gate19317(.O (g19244), .I1 (g18458), .I2 (g18514));
OR2X1 gate19318(.O (g19245), .I1 (g18395), .I2 (g18578));
OR2X1 gate19319(.O (g19246), .I1 (g18395), .I2 (g18478));
OR2X1 gate19320(.O (g19250), .I1 (g17729), .I2 (g17807));
OR3X1 gate19321(.O (I25516), .I1 (g17173), .I2 (g17160), .I3 (g17142));
OR3X1 gate19322(.O (g19253), .I1 (g17121), .I2 (g17085), .I3 (I25516));
OR2X1 gate19323(.O (g19255), .I1 (g14366), .I2 (g16523));
OR3X1 gate19324(.O (I25521), .I1 (g17093), .I2 (g17064), .I3 (g17046));
OR3X1 gate19325(.O (g19256), .I1 (g17019), .I2 (g16996), .I3 (I25521));
OR2X1 gate19326(.O (g19257), .I1 (g18531), .I2 (g18578));
OR2X1 gate19327(.O (g19263), .I1 (g17887), .I2 (g17979));
OR2X1 gate19328(.O (g19264), .I1 (g17830), .I2 (g17919));
OR3X1 gate19329(.O (I25549), .I1 (g17190), .I2 (g17175), .I3 (g17165));
OR3X1 gate19330(.O (g19266), .I1 (g17148), .I2 (g17123), .I3 (I25549));
OR2X1 gate19331(.O (g19268), .I1 (g14478), .I2 (g16554));
OR3X1 gate19332(.O (I25554), .I1 (g17131), .I2 (g17099), .I3 (g17080));
OR3X1 gate19333(.O (g19269), .I1 (g17049), .I2 (g17020), .I3 (I25554));
OR3X1 gate19334(.O (g19275), .I1 (g16867), .I2 (g16515), .I3 (g19001));
OR2X1 gate19335(.O (g19278), .I1 (g17998), .I2 (g18096));
OR2X1 gate19336(.O (g19279), .I1 (g17942), .I2 (g18030));
OR3X1 gate19337(.O (I25588), .I1 (g17201), .I2 (g17192), .I3 (g17180));
OR3X1 gate19338(.O (g19281), .I1 (g17171), .I2 (g17150), .I3 (I25588));
OR2X1 gate19339(.O (g19283), .I1 (g14565), .I2 (g16586));
OR3X1 gate19340(.O (g19294), .I1 (g16895), .I2 (g16546), .I3 (g16507));
OR2X1 gate19341(.O (g19297), .I1 (g18115), .I2 (g18212));
OR2X1 gate19342(.O (g19298), .I1 (g18053), .I2 (g18147));
OR3X1 gate19343(.O (g19312), .I1 (g16924), .I2 (g16578), .I3 (g16529));
OR2X1 gate19344(.O (g19315), .I1 (g18231), .I2 (g18319));
OR3X1 gate19345(.O (g19333), .I1 (g16954), .I2 (g16602), .I3 (g16560));
OR2X1 gate19346(.O (g19450), .I1 (g14837), .I2 (g16682));
OR2X1 gate19347(.O (g19477), .I1 (g14910), .I2 (g16708));
OR2X1 gate19348(.O (g19500), .I1 (g14991), .I2 (g16739));
OR3X1 gate19349(.O (g19503), .I1 (g16884), .I2 (g16697), .I3 (g16665));
OR2X1 gate19350(.O (g19521), .I1 (g15080), .I2 (g16781));
OR3X1 gate19351(.O (g19522), .I1 (g16913), .I2 (g16728), .I3 (g16686));
OR3X1 gate19352(.O (g19532), .I1 (g16943), .I2 (g16770), .I3 (g16712));
OR3X1 gate19353(.O (g19542), .I1 (g16974), .I2 (g16797), .I3 (g16743));
OR3X1 gate19354(.O (I26429), .I1 (g17979), .I2 (g17887), .I3 (g17807));
OR3X1 gate19355(.O (g19981), .I1 (g17729), .I2 (g18419), .I3 (I26429));
OR3X1 gate19356(.O (I26455), .I1 (g18424), .I2 (g18346), .I3 (g18270));
OR3X1 gate19357(.O (g20015), .I1 (g18183), .I2 (g18079), .I3 (I26455));
OR3X1 gate19358(.O (I26461), .I1 (g18096), .I2 (g17998), .I3 (g17919));
OR3X1 gate19359(.O (g20019), .I1 (g17830), .I2 (g18492), .I3 (I26461));
OR3X1 gate19360(.O (I26491), .I1 (g18497), .I2 (g18441), .I3 (g18363));
OR3X1 gate19361(.O (g20057), .I1 (g18290), .I2 (g18195), .I3 (I26491));
OR3X1 gate19362(.O (I26497), .I1 (g18212), .I2 (g18115), .I3 (g18030));
OR3X1 gate19363(.O (g20061), .I1 (g17942), .I2 (g18556), .I3 (I26497));
OR3X1 gate19364(.O (I26532), .I1 (g18561), .I2 (g18514), .I3 (g18458));
OR3X1 gate19365(.O (g20098), .I1 (g18383), .I2 (g18302), .I3 (I26532));
OR3X1 gate19366(.O (I26538), .I1 (g18319), .I2 (g18231), .I3 (g18147));
OR3X1 gate19367(.O (g20102), .I1 (g18053), .I2 (g18606), .I3 (I26538));
OR3X1 gate19368(.O (I26571), .I1 (g18611), .I2 (g18578), .I3 (g18531));
OR3X1 gate19369(.O (g20123), .I1 (g18478), .I2 (g18395), .I3 (I26571));
OR3X1 gate19370(.O (g21120), .I1 (g19484), .I2 (g16515), .I3 (g14071));
OR3X1 gate19371(.O (g21139), .I1 (g19505), .I2 (g16546), .I3 (g14186));
OR3X1 gate19372(.O (g21159), .I1 (g19524), .I2 (g16578), .I3 (g14301));
OR3X1 gate19373(.O (g21179), .I1 (g19534), .I2 (g16602), .I3 (g14423));
OR3X1 gate19374(.O (g21244), .I1 (g19578), .I2 (g16697), .I3 (g14776));
OR3X1 gate19375(.O (g21253), .I1 (g19608), .I2 (g16728), .I3 (g14811));
OR3X1 gate19376(.O (g21261), .I1 (g19641), .I2 (g16770), .I3 (g14863));
OR3X1 gate19377(.O (g21269), .I1 (g19681), .I2 (g16797), .I3 (g14936));
OR3X1 gate19378(.O (g21501), .I1 (g20522), .I2 (g16867), .I3 (g14071));
OR3X1 gate19379(.O (g21536), .I1 (g20522), .I2 (g19484), .I3 (g19001));
OR3X1 gate19380(.O (g21540), .I1 (g20542), .I2 (g16895), .I3 (g14186));
OR3X1 gate19381(.O (g21572), .I1 (g20542), .I2 (g19505), .I3 (g16507));
OR3X1 gate19382(.O (g21576), .I1 (g19067), .I2 (g16924), .I3 (g14301));
OR3X1 gate19383(.O (g21605), .I1 (g19067), .I2 (g19524), .I3 (g16529));
OR3X1 gate19384(.O (g21609), .I1 (g19084), .I2 (g16954), .I3 (g14423));
OR3X1 gate19385(.O (g21634), .I1 (g19084), .I2 (g19534), .I3 (g16560));
OR3X1 gate19386(.O (g21774), .I1 (g19121), .I2 (g16884), .I3 (g14776));
OR3X1 gate19387(.O (g21787), .I1 (g19121), .I2 (g19578), .I3 (g16665));
OR3X1 gate19388(.O (I28305), .I1 (g20197), .I2 (g20177), .I3 (g20145));
OR3X1 gate19389(.O (g21788), .I1 (g20117), .I2 (g20094), .I3 (I28305));
OR3X1 gate19390(.O (g21789), .I1 (g19128), .I2 (g16913), .I3 (g14811));
OR3X1 gate19391(.O (I28318), .I1 (g19092), .I2 (g19088), .I3 (g19079));
OR4X1 gate19392(.O (g21799), .I1 (g16505), .I2 (g20538), .I3 (g18994), .I4 (I28318));
OR4X1 gate19393(.O (g21800), .I1 (g18665), .I2 (g20270), .I3 (g20248), .I4 (g18647));
OR3X1 gate19394(.O (g21801), .I1 (g19128), .I2 (g19608), .I3 (g16686));
OR3X1 gate19395(.O (I28323), .I1 (g20227), .I2 (g20211), .I3 (g20183));
OR3X1 gate19396(.O (g21802), .I1 (g20147), .I2 (g20119), .I3 (I28323));
OR3X1 gate19397(.O (g21803), .I1 (g19135), .I2 (g16943), .I3 (g14863));
OR4X1 gate19398(.O (g21806), .I1 (g20116), .I2 (g20093), .I3 (g18547), .I4 (g19097));
OR3X1 gate19399(.O (I28330), .I1 (g19099), .I2 (g19094), .I3 (g19089));
OR4X1 gate19400(.O (g21807), .I1 (g16527), .I2 (g19063), .I3 (g19007), .I4 (I28330));
OR4X1 gate19401(.O (g21808), .I1 (g18688), .I2 (g20282), .I3 (g20271), .I4 (g18650));
OR3X1 gate19402(.O (g21809), .I1 (g19135), .I2 (g19641), .I3 (g16712));
OR3X1 gate19403(.O (I28335), .I1 (g20254), .I2 (g20241), .I3 (g20217));
OR3X1 gate19404(.O (g21810), .I1 (g20185), .I2 (g20149), .I3 (I28335));
OR3X1 gate19405(.O (g21811), .I1 (g19138), .I2 (g16974), .I3 (g14936));
OR4X1 gate19406(.O (g21813), .I1 (g20146), .I2 (g20118), .I3 (g18597), .I4 (g19104));
OR3X1 gate19407(.O (I28341), .I1 (g19106), .I2 (g19101), .I3 (g19095));
OR4X1 gate19408(.O (g21814), .I1 (g16558), .I2 (g19080), .I3 (g16513), .I4 (I28341));
OR4X1 gate19409(.O (g21815), .I1 (g18717), .I2 (g20293), .I3 (g20283), .I4 (g18654));
OR3X1 gate19410(.O (g21816), .I1 (g19138), .I2 (g19681), .I3 (g16743));
OR3X1 gate19411(.O (I28346), .I1 (g20277), .I2 (g20268), .I3 (g20247));
OR3X1 gate19412(.O (g21817), .I1 (g20219), .I2 (g20187), .I3 (I28346));
OR4X1 gate19413(.O (g21819), .I1 (g20184), .I2 (g20148), .I3 (g18629), .I4 (g19109));
OR3X1 gate19414(.O (I28351), .I1 (g19111), .I2 (g19108), .I3 (g19102));
OR4X1 gate19415(.O (g21820), .I1 (g16590), .I2 (g19090), .I3 (g16535), .I4 (I28351));
OR4X1 gate19416(.O (g21821), .I1 (g18753), .I2 (g20309), .I3 (g20294), .I4 (g18668));
OR4X1 gate19417(.O (g21823), .I1 (g20218), .I2 (g20186), .I3 (g18638), .I4 (g19116));
OR3X1 gate19418(.O (I28365), .I1 (g20280), .I2 (g18652), .I3 (g18649));
OR3X1 gate19419(.O (g21844), .I1 (g20222), .I2 (g18645), .I3 (I28365));
OR3X1 gate19420(.O (I28369), .I1 (g20291), .I2 (g18666), .I3 (g18653));
OR3X1 gate19421(.O (g21846), .I1 (g20249), .I2 (g18648), .I3 (I28369));
OR3X1 gate19422(.O (I28374), .I1 (g20307), .I2 (g18689), .I3 (g18667));
OR3X1 gate19423(.O (g21849), .I1 (g20272), .I2 (g18651), .I3 (I28374));
OR3X1 gate19424(.O (I28380), .I1 (g20326), .I2 (g18718), .I3 (g18690));
OR3X1 gate19425(.O (g21856), .I1 (g20284), .I2 (g18655), .I3 (I28380));
OR2X1 gate19426(.O (g22175), .I1 (g16075), .I2 (g20842));
OR2X1 gate19427(.O (g22190), .I1 (g16113), .I2 (g20850));
OR2X1 gate19428(.O (g22199), .I1 (g16164), .I2 (g20858));
OR2X1 gate19429(.O (g22205), .I1 (g16223), .I2 (g20866));
OR4X1 gate19430(.O (g22811), .I1 (g562), .I2 (g559), .I3 (g12451), .I4 (g21851));
OR3X1 gate19431(.O (g23052), .I1 (g21800), .I2 (g21788), .I3 (g21844));
OR3X1 gate19432(.O (g23071), .I1 (g21808), .I2 (g21802), .I3 (g21846));
OR3X1 gate19433(.O (g23084), .I1 (g21815), .I2 (g21810), .I3 (g21849));
OR2X1 gate19434(.O (g23089), .I1 (g21806), .I2 (g21799));
OR3X1 gate19435(.O (g23100), .I1 (g21821), .I2 (g21817), .I3 (g21856));
OR2X1 gate19436(.O (g23107), .I1 (g21813), .I2 (g21807));
OR2X1 gate19437(.O (g23120), .I1 (g21819), .I2 (g21814));
OR2X1 gate19438(.O (g23129), .I1 (g21823), .I2 (g21820));
OR2X1 gate19439(.O (g23319), .I1 (g14493), .I2 (g22385));
OR2X1 gate19440(.O (g23688), .I1 (g23106), .I2 (g21906));
OR2X1 gate19441(.O (g23742), .I1 (g23119), .I2 (g21920));
OR2X1 gate19442(.O (g23797), .I1 (g23128), .I2 (g21938));
OR2X1 gate19443(.O (g23850), .I1 (g23139), .I2 (g20647));
OR2X1 gate19444(.O (g23919), .I1 (g22666), .I2 (g23140));
OR2X1 gate19445(.O (g24239), .I1 (g19387), .I2 (g22401));
OR2X1 gate19446(.O (g24244), .I1 (g14144), .I2 (g22317));
OR2X1 gate19447(.O (g24245), .I1 (g19417), .I2 (g22402));
OR2X1 gate19448(.O (g24252), .I1 (g14259), .I2 (g22342));
OR2X1 gate19449(.O (g24254), .I1 (g19454), .I2 (g22403));
OR2X1 gate19450(.O (g24257), .I1 (g14381), .I2 (g22365));
OR2X1 gate19451(.O (g24258), .I1 (g19481), .I2 (g22404));
OR2X1 gate19452(.O (g24633), .I1 (g24094), .I2 (g20842));
OR2X1 gate19453(.O (g24653), .I1 (g24095), .I2 (g20850));
OR2X1 gate19454(.O (g24672), .I1 (g24097), .I2 (g20858));
OR2X1 gate19455(.O (g24691), .I1 (g24103), .I2 (g20866));
OR2X1 gate19456(.O (g24890), .I1 (g23639), .I2 (g23144));
OR2X1 gate19457(.O (g24909), .I1 (g23726), .I2 (g23142));
OR2X1 gate19458(.O (g24925), .I1 (g23772), .I2 (g23141));
OR2X1 gate19459(.O (g24965), .I1 (g23922), .I2 (g23945));
OR2X1 gate19460(.O (g24978), .I1 (g23954), .I2 (g23974));
OR2X1 gate19461(.O (g24989), .I1 (g23983), .I2 (g24004));
OR2X1 gate19462(.O (g25000), .I1 (g24013), .I2 (g24038));
OR2X1 gate19463(.O (g25183), .I1 (g24958), .I2 (g24893));
OR2X1 gate19464(.O (g25186), .I1 (g24969), .I2 (g24916));
OR2X1 gate19465(.O (g25190), .I1 (g24982), .I2 (g24933));
OR2X1 gate19466(.O (g25195), .I1 (g24993), .I2 (g24945));
OR2X1 gate19467(.O (g25489), .I1 (g24795), .I2 (g16466));
OR2X1 gate19468(.O (g25490), .I1 (g24759), .I2 (g23146));
OR2X1 gate19469(.O (g25520), .I1 (g24813), .I2 (g23145));
OR2X1 gate19470(.O (g25566), .I1 (g24843), .I2 (g23143));
OR2X1 gate19471(.O (g26320), .I1 (g25852), .I2 (g25870));
OR2X1 gate19472(.O (g26367), .I1 (g25873), .I2 (g25882));
OR2X1 gate19473(.O (g26410), .I1 (g25885), .I2 (g25887));
OR2X1 gate19474(.O (g26451), .I1 (g25890), .I2 (g25892));
OR2X1 gate19475(.O (g26974), .I1 (g26157), .I2 (g23147));
OR3X1 gate19476(.O (g27113), .I1 (g1248), .I2 (g1245), .I3 (g26534));
OR2X1 gate19477(.O (g28501), .I1 (g27738), .I2 (g25764));
OR2X1 gate19478(.O (g28512), .I1 (g26481), .I2 (g27738));
OR2X1 gate19479(.O (g28529), .I1 (g27743), .I2 (g25818));
OR2X1 gate19480(.O (g28540), .I1 (g26497), .I2 (g27743));
OR2X1 gate19481(.O (g28556), .I1 (g27751), .I2 (g25853));
OR2X1 gate19482(.O (g28567), .I1 (g26512), .I2 (g27751));
OR2X1 gate19483(.O (g28584), .I1 (g27756), .I2 (g25874));
OR2X1 gate19484(.O (g28595), .I1 (g26520), .I2 (g27756));
OR3X1 gate19485(.O (g29348), .I1 (g1942), .I2 (g1939), .I3 (g29113));
OR3X1 gate19486(.O (g30305), .I1 (g2636), .I2 (g2633), .I3 (g30072));
ND2X1 gate19487(.O (I15167), .I1 (g2981), .I2 (g2874));
ND2X1 gate19488(.O (I15168), .I1 (g2981), .I2 (I15167));
ND2X1 gate19489(.O (I15169), .I1 (g2874), .I2 (I15167));
ND2X1 gate19490(.O (g7855), .I1 (I15168), .I2 (I15169));
ND2X1 gate19491(.O (I15183), .I1 (g2975), .I2 (g2978));
ND2X1 gate19492(.O (I15184), .I1 (g2975), .I2 (I15183));
ND2X1 gate19493(.O (I15185), .I1 (g2978), .I2 (I15183));
ND2X1 gate19494(.O (g7875), .I1 (I15184), .I2 (I15185));
ND2X1 gate19495(.O (I15190), .I1 (g2956), .I2 (g2959));
ND2X1 gate19496(.O (I15191), .I1 (g2956), .I2 (I15190));
ND2X1 gate19497(.O (I15192), .I1 (g2959), .I2 (I15190));
ND2X1 gate19498(.O (g7876), .I1 (I15191), .I2 (I15192));
ND2X1 gate19499(.O (I15204), .I1 (g2969), .I2 (g2972));
ND2X1 gate19500(.O (I15205), .I1 (g2969), .I2 (I15204));
ND2X1 gate19501(.O (I15206), .I1 (g2972), .I2 (I15204));
ND2X1 gate19502(.O (g7895), .I1 (I15205), .I2 (I15206));
ND2X1 gate19503(.O (I15211), .I1 (g2947), .I2 (g2953));
ND2X1 gate19504(.O (I15212), .I1 (g2947), .I2 (I15211));
ND2X1 gate19505(.O (I15213), .I1 (g2953), .I2 (I15211));
ND2X1 gate19506(.O (g7896), .I1 (I15212), .I2 (I15213));
ND2X1 gate19507(.O (I15237), .I1 (g2963), .I2 (g2966));
ND2X1 gate19508(.O (I15238), .I1 (g2963), .I2 (I15237));
ND2X1 gate19509(.O (I15239), .I1 (g2966), .I2 (I15237));
ND2X1 gate19510(.O (g7922), .I1 (I15238), .I2 (I15239));
ND2X1 gate19511(.O (I15244), .I1 (g2941), .I2 (g2944));
ND2X1 gate19512(.O (I15245), .I1 (g2941), .I2 (I15244));
ND2X1 gate19513(.O (I15246), .I1 (g2944), .I2 (I15244));
ND2X1 gate19514(.O (g7923), .I1 (I15245), .I2 (I15246));
ND2X1 gate19515(.O (I15276), .I1 (g2935), .I2 (g2938));
ND2X1 gate19516(.O (I15277), .I1 (g2935), .I2 (I15276));
ND2X1 gate19517(.O (I15278), .I1 (g2938), .I2 (I15276));
ND2X1 gate19518(.O (g7970), .I1 (I15277), .I2 (I15278));
ND4X1 gate19519(.O (g8381), .I1 (g8182), .I2 (g8120), .I3 (g8044), .I4 (g7989));
ND2X1 gate19520(.O (g8533), .I1 (g3398), .I2 (g3366));
ND2X1 gate19521(.O (g8547), .I1 (g3398), .I2 (g3366));
ND2X1 gate19522(.O (g8550), .I1 (g3554), .I2 (g3522));
ND2X1 gate19523(.O (g8560), .I1 (g3554), .I2 (g3522));
ND2X1 gate19524(.O (g8563), .I1 (g3710), .I2 (g3678));
ND2X1 gate19525(.O (g8571), .I1 (g3710), .I2 (g3678));
ND2X1 gate19526(.O (g8574), .I1 (g3866), .I2 (g3834));
ND2X1 gate19527(.O (g8577), .I1 (g3866), .I2 (g3834));
ND2X1 gate19528(.O (I16879), .I1 (g4203), .I2 (g3998));
ND2X1 gate19529(.O (I16880), .I1 (g4203), .I2 (I16879));
ND2X1 gate19530(.O (I16881), .I1 (g3998), .I2 (I16879));
ND2X1 gate19531(.O (g9883), .I1 (I16880), .I2 (I16881));
ND2X1 gate19532(.O (I16965), .I1 (g4734), .I2 (g4452));
ND2X1 gate19533(.O (I16966), .I1 (g4734), .I2 (I16965));
ND2X1 gate19534(.O (I16967), .I1 (g4452), .I2 (I16965));
ND2X1 gate19535(.O (g10003), .I1 (I16966), .I2 (I16967));
ND2X1 gate19536(.O (g10038), .I1 (g7772), .I2 (g3366));
ND2X1 gate19537(.O (I17059), .I1 (g6637), .I2 (g6309));
ND2X1 gate19538(.O (I17060), .I1 (g6637), .I2 (I17059));
ND2X1 gate19539(.O (I17061), .I1 (g6309), .I2 (I17059));
ND2X1 gate19540(.O (g10095), .I1 (I17060), .I2 (I17061));
ND2X1 gate19541(.O (g10147), .I1 (g7788), .I2 (g3522));
ND2X1 gate19542(.O (I17149), .I1 (g7465), .I2 (g7142));
ND2X1 gate19543(.O (I17150), .I1 (g7465), .I2 (I17149));
ND2X1 gate19544(.O (I17151), .I1 (g7142), .I2 (I17149));
ND2X1 gate19545(.O (g10185), .I1 (I17150), .I2 (I17151));
ND2X1 gate19546(.O (g10252), .I1 (g7802), .I2 (g3678));
ND2X1 gate19547(.O (g10354), .I1 (g7815), .I2 (g3834));
ND2X1 gate19548(.O (g10649), .I1 (g3398), .I2 (g6912));
ND2X1 gate19549(.O (g10676), .I1 (g3398), .I2 (g6678));
ND2X1 gate19550(.O (g10677), .I1 (g3398), .I2 (g6912));
ND2X1 gate19551(.O (g10679), .I1 (g3554), .I2 (g7162));
ND2X1 gate19552(.O (g10703), .I1 (g3398), .I2 (g6678));
ND2X1 gate19553(.O (g10705), .I1 (g3554), .I2 (g6980));
ND2X1 gate19554(.O (g10706), .I1 (g3554), .I2 (g7162));
ND2X1 gate19555(.O (g10708), .I1 (g3710), .I2 (g7358));
ND2X1 gate19556(.O (g10723), .I1 (g3554), .I2 (g6980));
ND2X1 gate19557(.O (g10725), .I1 (g3710), .I2 (g7230));
ND2X1 gate19558(.O (g10726), .I1 (g3710), .I2 (g7358));
ND2X1 gate19559(.O (g10728), .I1 (g3866), .I2 (g7488));
ND2X1 gate19560(.O (g10744), .I1 (g3710), .I2 (g7230));
ND2X1 gate19561(.O (g10746), .I1 (g3866), .I2 (g7426));
ND2X1 gate19562(.O (g10747), .I1 (g3866), .I2 (g7488));
ND2X1 gate19563(.O (g10763), .I1 (g3866), .I2 (g7426));
ND2X1 gate19564(.O (I18106), .I1 (g7875), .I2 (g7855));
ND2X1 gate19565(.O (I18107), .I1 (g7875), .I2 (I18106));
ND2X1 gate19566(.O (I18108), .I1 (g7855), .I2 (I18106));
ND2X1 gate19567(.O (g11188), .I1 (I18107), .I2 (I18108));
ND2X1 gate19568(.O (I18113), .I1 (g3997), .I2 (g8181));
ND2X1 gate19569(.O (I18114), .I1 (g3997), .I2 (I18113));
ND2X1 gate19570(.O (I18115), .I1 (g8181), .I2 (I18113));
ND2X1 gate19571(.O (g11189), .I1 (I18114), .I2 (I18115));
ND2X1 gate19572(.O (I18190), .I1 (g7922), .I2 (g7895));
ND2X1 gate19573(.O (I18191), .I1 (g7922), .I2 (I18190));
ND2X1 gate19574(.O (I18192), .I1 (g7895), .I2 (I18190));
ND2X1 gate19575(.O (g11262), .I1 (I18191), .I2 (I18192));
ND2X1 gate19576(.O (I18197), .I1 (g7896), .I2 (g7876));
ND2X1 gate19577(.O (I18198), .I1 (g7896), .I2 (I18197));
ND2X1 gate19578(.O (I18199), .I1 (g7876), .I2 (I18197));
ND2X1 gate19579(.O (g11263), .I1 (I18198), .I2 (I18199));
ND2X1 gate19580(.O (I18204), .I1 (g7975), .I2 (g4202));
ND2X1 gate19581(.O (I18205), .I1 (g7975), .I2 (I18204));
ND2X1 gate19582(.O (I18206), .I1 (g4202), .I2 (I18204));
ND2X1 gate19583(.O (g11264), .I1 (I18205), .I2 (I18206));
ND2X1 gate19584(.O (I18280), .I1 (g7970), .I2 (g7923));
ND2X1 gate19585(.O (I18281), .I1 (g7970), .I2 (I18280));
ND2X1 gate19586(.O (I18282), .I1 (g7923), .I2 (I18280));
ND2X1 gate19587(.O (g11330), .I1 (I18281), .I2 (I18282));
ND2X1 gate19588(.O (I18287), .I1 (g8256), .I2 (g8102));
ND2X1 gate19589(.O (I18288), .I1 (g8256), .I2 (I18287));
ND2X1 gate19590(.O (I18289), .I1 (g8102), .I2 (I18287));
ND2X1 gate19591(.O (g11331), .I1 (I18288), .I2 (I18289));
ND2X1 gate19592(.O (I18368), .I1 (g4325), .I2 (g4093));
ND2X1 gate19593(.O (I18369), .I1 (g4325), .I2 (I18368));
ND2X1 gate19594(.O (I18370), .I1 (g4093), .I2 (I18368));
ND2X1 gate19595(.O (g11410), .I1 (I18369), .I2 (I18370));
ND2X1 gate19596(.O (g11617), .I1 (g8313), .I2 (g2883));
ND2X1 gate19597(.O (I18799), .I1 (g11410), .I2 (g11331));
ND2X1 gate19598(.O (I18800), .I1 (g11410), .I2 (I18799));
ND2X1 gate19599(.O (I18801), .I1 (g11331), .I2 (I18799));
ND2X1 gate19600(.O (g11621), .I1 (I18800), .I2 (I18801));
ND2X1 gate19601(.O (g11661), .I1 (g9534), .I2 (g3366));
ND2X1 gate19602(.O (g11662), .I1 (g9534), .I2 (g3366));
ND2X1 gate19603(.O (g11672), .I1 (g9534), .I2 (g3366));
ND2X1 gate19604(.O (g11673), .I1 (g9676), .I2 (g3522));
ND2X1 gate19605(.O (g11674), .I1 (g9676), .I2 (g3522));
ND2X1 gate19606(.O (g11683), .I1 (g9534), .I2 (g3366));
ND2X1 gate19607(.O (g11684), .I1 (g9676), .I2 (g3522));
ND2X1 gate19608(.O (g11685), .I1 (g9822), .I2 (g3678));
ND2X1 gate19609(.O (g11686), .I1 (g9822), .I2 (g3678));
ND2X1 gate19610(.O (g11691), .I1 (g9534), .I2 (g3366));
ND2X1 gate19611(.O (g11692), .I1 (g9676), .I2 (g3522));
ND2X1 gate19612(.O (g11693), .I1 (g9822), .I2 (g3678));
ND2X1 gate19613(.O (g11694), .I1 (g9968), .I2 (g3834));
ND2X1 gate19614(.O (g11695), .I1 (g9968), .I2 (g3834));
ND2X1 gate19615(.O (g11696), .I1 (g9534), .I2 (g3366));
ND2X1 gate19616(.O (g11698), .I1 (g9676), .I2 (g3522));
ND2X1 gate19617(.O (g11699), .I1 (g9822), .I2 (g3678));
ND2X1 gate19618(.O (g11700), .I1 (g9968), .I2 (g3834));
ND2X1 gate19619(.O (g11701), .I1 (g9534), .I2 (g3366));
ND2X1 gate19620(.O (g11702), .I1 (g9676), .I2 (g3522));
ND2X1 gate19621(.O (g11704), .I1 (g9822), .I2 (g3678));
ND2X1 gate19622(.O (g11705), .I1 (g9968), .I2 (g3834));
ND2X1 gate19623(.O (g11707), .I1 (g9534), .I2 (g3366));
ND2X1 gate19624(.O (g11708), .I1 (g9534), .I2 (g3366));
ND2X1 gate19625(.O (g11709), .I1 (g9676), .I2 (g3522));
ND2X1 gate19626(.O (g11710), .I1 (g9822), .I2 (g3678));
ND2X1 gate19627(.O (g11712), .I1 (g9968), .I2 (g3834));
ND2X1 gate19628(.O (g11713), .I1 (g10481), .I2 (g9144));
ND2X1 gate19629(.O (g11716), .I1 (g9534), .I2 (g3366));
ND2X1 gate19630(.O (g11717), .I1 (g9676), .I2 (g3522));
ND2X1 gate19631(.O (g11718), .I1 (g9676), .I2 (g3522));
ND2X1 gate19632(.O (g11719), .I1 (g9822), .I2 (g3678));
ND2X1 gate19633(.O (g11720), .I1 (g9968), .I2 (g3834));
ND2X1 gate19634(.O (g11721), .I1 (g9534), .I2 (g3366));
ND2X1 gate19635(.O (g11722), .I1 (g9676), .I2 (g3522));
ND2X1 gate19636(.O (g11723), .I1 (g9822), .I2 (g3678));
ND2X1 gate19637(.O (g11724), .I1 (g9822), .I2 (g3678));
ND2X1 gate19638(.O (g11725), .I1 (g9968), .I2 (g3834));
ND2X1 gate19639(.O (g11726), .I1 (g9676), .I2 (g3522));
ND2X1 gate19640(.O (g11727), .I1 (g9822), .I2 (g3678));
ND2X1 gate19641(.O (g11728), .I1 (g9968), .I2 (g3834));
ND2X1 gate19642(.O (g11729), .I1 (g9968), .I2 (g3834));
ND2X1 gate19643(.O (g11730), .I1 (g9822), .I2 (g3678));
ND2X1 gate19644(.O (g11731), .I1 (g9968), .I2 (g3834));
ND2X1 gate19645(.O (g11733), .I1 (g9968), .I2 (g3834));
ND2X1 gate19646(.O (g12433), .I1 (g2879), .I2 (g10778));
ND2X1 gate19647(.O (g12486), .I1 (g8278), .I2 (g6448));
ND2X1 gate19648(.O (g12503), .I1 (g8278), .I2 (g5438));
ND2X1 gate19649(.O (g12506), .I1 (g8287), .I2 (g6713));
ND2X1 gate19650(.O (g12520), .I1 (g8287), .I2 (g5473));
ND2X1 gate19651(.O (g12523), .I1 (g8296), .I2 (g7015));
ND2X1 gate19652(.O (g12535), .I1 (g8296), .I2 (g5512));
ND2X1 gate19653(.O (g12538), .I1 (g8305), .I2 (g7265));
ND2X1 gate19654(.O (g12544), .I1 (g8305), .I2 (g5556));
ND2X1 gate19655(.O (I20031), .I1 (g10003), .I2 (g9883));
ND2X1 gate19656(.O (I20032), .I1 (g10003), .I2 (I20031));
ND2X1 gate19657(.O (I20033), .I1 (g9883), .I2 (I20031));
ND2X1 gate19658(.O (g12988), .I1 (I20032), .I2 (I20033));
ND2X1 gate19659(.O (I20048), .I1 (g10185), .I2 (g10095));
ND2X1 gate19660(.O (I20049), .I1 (g10185), .I2 (I20048));
ND2X1 gate19661(.O (I20050), .I1 (g10095), .I2 (I20048));
ND2X1 gate19662(.O (g12999), .I1 (I20049), .I2 (I20050));
ND2X1 gate19663(.O (g13020), .I1 (g9534), .I2 (g6912));
ND2X1 gate19664(.O (g13021), .I1 (g9534), .I2 (g6912));
ND2X1 gate19665(.O (g13026), .I1 (g9534), .I2 (g6678));
ND2X1 gate19666(.O (g13027), .I1 (g9534), .I2 (g6912));
ND2X1 gate19667(.O (g13028), .I1 (g9534), .I2 (g6678));
ND2X1 gate19668(.O (g13029), .I1 (g9676), .I2 (g7162));
ND2X1 gate19669(.O (g13030), .I1 (g9676), .I2 (g7162));
ND2X1 gate19670(.O (g13034), .I1 (g9534), .I2 (g6678));
ND2X1 gate19671(.O (g13035), .I1 (g9534), .I2 (g6912));
ND2X1 gate19672(.O (g13037), .I1 (g9676), .I2 (g6980));
ND2X1 gate19673(.O (g13038), .I1 (g9676), .I2 (g7162));
ND2X1 gate19674(.O (g13039), .I1 (g9676), .I2 (g6980));
ND2X1 gate19675(.O (g13040), .I1 (g9822), .I2 (g7358));
ND2X1 gate19676(.O (g13041), .I1 (g9822), .I2 (g7358));
ND2X1 gate19677(.O (g13044), .I1 (g9534), .I2 (g6678));
ND2X1 gate19678(.O (g13045), .I1 (g9534), .I2 (g6912));
ND2X1 gate19679(.O (g13047), .I1 (g9676), .I2 (g6980));
ND2X1 gate19680(.O (g13048), .I1 (g9676), .I2 (g7162));
ND2X1 gate19681(.O (g13050), .I1 (g9822), .I2 (g7230));
ND2X1 gate19682(.O (g13051), .I1 (g9822), .I2 (g7358));
ND2X1 gate19683(.O (g13052), .I1 (g9822), .I2 (g7230));
ND2X1 gate19684(.O (g13053), .I1 (g9968), .I2 (g7488));
ND2X1 gate19685(.O (g13054), .I1 (g9968), .I2 (g7488));
ND2X1 gate19686(.O (g13058), .I1 (g9534), .I2 (g6678));
ND2X1 gate19687(.O (g13059), .I1 (g9534), .I2 (g6912));
ND2X1 gate19688(.O (g13061), .I1 (g9676), .I2 (g6980));
ND2X1 gate19689(.O (g13062), .I1 (g9676), .I2 (g7162));
ND2X1 gate19690(.O (g13064), .I1 (g9822), .I2 (g7230));
ND2X1 gate19691(.O (g13065), .I1 (g9822), .I2 (g7358));
ND2X1 gate19692(.O (g13067), .I1 (g9968), .I2 (g7426));
ND2X1 gate19693(.O (g13068), .I1 (g9968), .I2 (g7488));
ND2X1 gate19694(.O (g13069), .I1 (g9968), .I2 (g7426));
ND2X1 gate19695(.O (g13071), .I1 (g9534), .I2 (g6678));
ND2X1 gate19696(.O (g13072), .I1 (g9534), .I2 (g6912));
ND2X1 gate19697(.O (g13074), .I1 (g9676), .I2 (g6980));
ND2X1 gate19698(.O (g13075), .I1 (g9676), .I2 (g7162));
ND2X1 gate19699(.O (g13077), .I1 (g9822), .I2 (g7230));
ND2X1 gate19700(.O (g13078), .I1 (g9822), .I2 (g7358));
ND2X1 gate19701(.O (g13080), .I1 (g9968), .I2 (g7426));
ND2X1 gate19702(.O (g13081), .I1 (g9968), .I2 (g7488));
ND2X1 gate19703(.O (g13087), .I1 (g9534), .I2 (g6678));
ND2X1 gate19704(.O (g13088), .I1 (g9534), .I2 (g6912));
ND2X1 gate19705(.O (g13089), .I1 (g9534), .I2 (g6912));
ND2X1 gate19706(.O (g13090), .I1 (g9676), .I2 (g6980));
ND2X1 gate19707(.O (g13091), .I1 (g9676), .I2 (g7162));
ND2X1 gate19708(.O (g13093), .I1 (g9822), .I2 (g7230));
ND2X1 gate19709(.O (g13094), .I1 (g9822), .I2 (g7358));
ND2X1 gate19710(.O (g13096), .I1 (g9968), .I2 (g7426));
ND2X1 gate19711(.O (g13097), .I1 (g9968), .I2 (g7488));
ND2X1 gate19712(.O (g13098), .I1 (g9534), .I2 (g6678));
ND2X1 gate19713(.O (g13099), .I1 (g9534), .I2 (g6912));
ND2X1 gate19714(.O (g13100), .I1 (g9534), .I2 (g6678));
ND2X1 gate19715(.O (g13102), .I1 (g9676), .I2 (g6980));
ND2X1 gate19716(.O (g13103), .I1 (g9676), .I2 (g7162));
ND2X1 gate19717(.O (g13104), .I1 (g9676), .I2 (g7162));
ND2X1 gate19718(.O (g13105), .I1 (g9822), .I2 (g7230));
ND2X1 gate19719(.O (g13106), .I1 (g9822), .I2 (g7358));
ND2X1 gate19720(.O (g13108), .I1 (g9968), .I2 (g7426));
ND2X1 gate19721(.O (g13109), .I1 (g9968), .I2 (g7488));
ND2X1 gate19722(.O (g13112), .I1 (g9534), .I2 (g6678));
ND2X1 gate19723(.O (g13113), .I1 (g9534), .I2 (g6912));
ND2X1 gate19724(.O (g13114), .I1 (g9676), .I2 (g6980));
ND2X1 gate19725(.O (g13115), .I1 (g9676), .I2 (g7162));
ND2X1 gate19726(.O (g13116), .I1 (g9676), .I2 (g6980));
ND2X1 gate19727(.O (g13118), .I1 (g9822), .I2 (g7230));
ND2X1 gate19728(.O (g13119), .I1 (g9822), .I2 (g7358));
ND2X1 gate19729(.O (g13120), .I1 (g9822), .I2 (g7358));
ND2X1 gate19730(.O (g13121), .I1 (g9968), .I2 (g7426));
ND2X1 gate19731(.O (g13122), .I1 (g9968), .I2 (g7488));
ND2X1 gate19732(.O (g13123), .I1 (g9534), .I2 (g6678));
ND2X1 gate19733(.O (g13125), .I1 (g9676), .I2 (g6980));
ND2X1 gate19734(.O (g13126), .I1 (g9676), .I2 (g7162));
ND2X1 gate19735(.O (g13127), .I1 (g9822), .I2 (g7230));
ND2X1 gate19736(.O (g13128), .I1 (g9822), .I2 (g7358));
ND2X1 gate19737(.O (g13129), .I1 (g9822), .I2 (g7230));
ND2X1 gate19738(.O (g13131), .I1 (g9968), .I2 (g7426));
ND2X1 gate19739(.O (g13132), .I1 (g9968), .I2 (g7488));
ND2X1 gate19740(.O (g13133), .I1 (g9968), .I2 (g7488));
ND2X1 gate19741(.O (g13134), .I1 (g9676), .I2 (g6980));
ND2X1 gate19742(.O (g13136), .I1 (g9822), .I2 (g7230));
ND2X1 gate19743(.O (g13137), .I1 (g9822), .I2 (g7358));
ND2X1 gate19744(.O (g13138), .I1 (g9968), .I2 (g7426));
ND2X1 gate19745(.O (g13139), .I1 (g9968), .I2 (g7488));
ND2X1 gate19746(.O (g13140), .I1 (g9968), .I2 (g7426));
ND2X1 gate19747(.O (g13142), .I1 (g9822), .I2 (g7230));
ND2X1 gate19748(.O (g13144), .I1 (g9968), .I2 (g7426));
ND2X1 gate19749(.O (g13145), .I1 (g9968), .I2 (g7488));
ND2X1 gate19750(.O (g13146), .I1 (g9968), .I2 (g7426));
ND2X1 gate19751(.O (g13147), .I1 (g8278), .I2 (g3306));
ND2X1 gate19752(.O (g13150), .I1 (g8287), .I2 (g3462));
ND2X1 gate19753(.O (g13156), .I1 (g8296), .I2 (g3618));
ND2X1 gate19754(.O (g13165), .I1 (g8305), .I2 (g3774));
ND2X1 gate19755(.O (g13245), .I1 (g10779), .I2 (g7901));
ND2X1 gate19756(.O (g13305), .I1 (g8317), .I2 (g2993));
ND2X1 gate19757(.O (I20429), .I1 (g11262), .I2 (g11188));
ND2X1 gate19758(.O (I20430), .I1 (g11262), .I2 (I20429));
ND2X1 gate19759(.O (I20431), .I1 (g11188), .I2 (I20429));
ND2X1 gate19760(.O (g13348), .I1 (I20430), .I2 (I20431));
ND2X1 gate19761(.O (I20465), .I1 (g11330), .I2 (g11263));
ND2X1 gate19762(.O (I20466), .I1 (g11330), .I2 (I20465));
ND2X1 gate19763(.O (I20467), .I1 (g11263), .I2 (I20465));
ND2X1 gate19764(.O (g13370), .I1 (I20466), .I2 (I20467));
ND2X1 gate19765(.O (I20504), .I1 (g11264), .I2 (g11189));
ND2X1 gate19766(.O (I20505), .I1 (g11264), .I2 (I20504));
ND2X1 gate19767(.O (I20506), .I1 (g11189), .I2 (I20504));
ND2X1 gate19768(.O (g13399), .I1 (I20505), .I2 (I20506));
ND2X1 gate19769(.O (g13476), .I1 (g12565), .I2 (g3254));
ND2X1 gate19770(.O (g13478), .I1 (g12611), .I2 (g3410));
ND2X1 gate19771(.O (g13482), .I1 (g12657), .I2 (g3566));
ND2X1 gate19772(.O (g13494), .I1 (g12565), .I2 (g3254));
ND2X1 gate19773(.O (g13495), .I1 (g12611), .I2 (g3410));
ND2X1 gate19774(.O (g13497), .I1 (g12657), .I2 (g3566));
ND2X1 gate19775(.O (g13501), .I1 (g12711), .I2 (g3722));
ND2X1 gate19776(.O (I20743), .I1 (g11621), .I2 (g13399));
ND2X1 gate19777(.O (I20744), .I1 (g11621), .I2 (I20743));
ND2X1 gate19778(.O (I20745), .I1 (g13399), .I2 (I20743));
ND2X1 gate19779(.O (g13507), .I1 (I20744), .I2 (I20745));
ND2X1 gate19780(.O (g13510), .I1 (g12565), .I2 (g3254));
ND2X1 gate19781(.O (g13511), .I1 (g12611), .I2 (g3410));
ND2X1 gate19782(.O (g13512), .I1 (g12657), .I2 (g3566));
ND2X1 gate19783(.O (g13514), .I1 (g12711), .I2 (g3722));
ND2X1 gate19784(.O (g13518), .I1 (g12565), .I2 (g3254));
ND2X1 gate19785(.O (g13524), .I1 (g12611), .I2 (g3410));
ND2X1 gate19786(.O (g13525), .I1 (g12657), .I2 (g3566));
ND2X1 gate19787(.O (g13526), .I1 (g12711), .I2 (g3722));
ND2X1 gate19788(.O (g13528), .I1 (g12565), .I2 (g3254));
ND2X1 gate19789(.O (g13529), .I1 (g12611), .I2 (g3410));
ND2X1 gate19790(.O (g13535), .I1 (g12657), .I2 (g3566));
ND2X1 gate19791(.O (g13536), .I1 (g12711), .I2 (g3722));
ND2X1 gate19792(.O (g13537), .I1 (g12565), .I2 (g3254));
ND2X1 gate19793(.O (g13538), .I1 (g12565), .I2 (g3254));
ND2X1 gate19794(.O (g13539), .I1 (g12611), .I2 (g3410));
ND2X1 gate19795(.O (g13540), .I1 (g12657), .I2 (g3566));
ND2X1 gate19796(.O (g13546), .I1 (g12711), .I2 (g3722));
ND2X1 gate19797(.O (g13547), .I1 (g12565), .I2 (g3254));
ND2X1 gate19798(.O (g13548), .I1 (g12611), .I2 (g3410));
ND2X1 gate19799(.O (g13549), .I1 (g12611), .I2 (g3410));
ND2X1 gate19800(.O (g13550), .I1 (g12657), .I2 (g3566));
ND2X1 gate19801(.O (g13551), .I1 (g12711), .I2 (g3722));
ND2X1 gate19802(.O (g13557), .I1 (g12611), .I2 (g3410));
ND2X1 gate19803(.O (g13558), .I1 (g12657), .I2 (g3566));
ND2X1 gate19804(.O (g13559), .I1 (g12657), .I2 (g3566));
ND2X1 gate19805(.O (g13560), .I1 (g12711), .I2 (g3722));
ND2X1 gate19806(.O (g13561), .I1 (g12657), .I2 (g3566));
ND2X1 gate19807(.O (g13562), .I1 (g12711), .I2 (g3722));
ND2X1 gate19808(.O (g13563), .I1 (g12711), .I2 (g3722));
ND2X1 gate19809(.O (g13564), .I1 (g12711), .I2 (g3722));
ND2X1 gate19810(.O (g13599), .I1 (g12886), .I2 (g3366));
ND2X1 gate19811(.O (g13611), .I1 (g12926), .I2 (g3522));
ND2X1 gate19812(.O (g13621), .I1 (g12955), .I2 (g3678));
ND2X1 gate19813(.O (g13633), .I1 (g12984), .I2 (g3834));
ND2X1 gate19814(.O (g13893), .I1 (g8580), .I2 (g12463));
ND3X1 gate19815(.O (g13915), .I1 (g8822), .I2 (g12473), .I3 (g12463));
ND2X1 gate19816(.O (g13934), .I1 (g8587), .I2 (g12478));
ND2X1 gate19817(.O (g13957), .I1 (g10730), .I2 (g12473));
ND3X1 gate19818(.O (g13971), .I1 (g8846), .I2 (g12490), .I3 (g12478));
ND2X1 gate19819(.O (g13990), .I1 (g8594), .I2 (g12495));
ND2X1 gate19820(.O (g14027), .I1 (g10749), .I2 (g12490));
ND3X1 gate19821(.O (g14041), .I1 (g8873), .I2 (g12510), .I3 (g12495));
ND2X1 gate19822(.O (g14060), .I1 (g8605), .I2 (g12515));
ND2X1 gate19823(.O (g14118), .I1 (g10767), .I2 (g12510));
ND3X1 gate19824(.O (g14132), .I1 (g8911), .I2 (g12527), .I3 (g12515));
ND2X1 gate19825(.O (g14233), .I1 (g10773), .I2 (g12527));
ND3X1 gate19826(.O (g15454), .I1 (g9232), .I2 (g9150), .I3 (g12780));
ND3X1 gate19827(.O (g15540), .I1 (g9310), .I2 (g9174), .I3 (g12819));
ND3X1 gate19828(.O (g15618), .I1 (g9391), .I2 (g9216), .I3 (g12857));
ND2X1 gate19829(.O (g15660), .I1 (g13401), .I2 (g12354));
ND2X1 gate19830(.O (g15664), .I1 (g12565), .I2 (g6314));
ND3X1 gate19831(.O (g15694), .I1 (g9488), .I2 (g9277), .I3 (g12898));
ND2X1 gate19832(.O (g15718), .I1 (g13286), .I2 (g12354));
ND2X1 gate19833(.O (g15719), .I1 (g13401), .I2 (g12392));
ND2X1 gate19834(.O (g15720), .I1 (g12565), .I2 (g6232));
ND2X1 gate19835(.O (g15721), .I1 (g12565), .I2 (g6314));
ND2X1 gate19836(.O (g15723), .I1 (g12611), .I2 (g6519));
ND2X1 gate19837(.O (g15756), .I1 (g13313), .I2 (g12354));
ND2X1 gate19838(.O (g15757), .I1 (g11622), .I2 (g12392));
ND2X1 gate19839(.O (g15758), .I1 (g12565), .I2 (g6232));
ND2X1 gate19840(.O (g15759), .I1 (g12565), .I2 (g6314));
ND2X1 gate19841(.O (g15760), .I1 (g12611), .I2 (g6369));
ND2X1 gate19842(.O (g15761), .I1 (g12611), .I2 (g6519));
ND2X1 gate19843(.O (g15763), .I1 (g12657), .I2 (g6783));
ND2X1 gate19844(.O (g15782), .I1 (g13332), .I2 (g12354));
ND2X1 gate19845(.O (g15783), .I1 (g11643), .I2 (g12392));
ND2X1 gate19846(.O (g15784), .I1 (g12565), .I2 (g6232));
ND2X1 gate19847(.O (g15785), .I1 (g12565), .I2 (g6314));
ND2X1 gate19848(.O (g15786), .I1 (g12611), .I2 (g6369));
ND2X1 gate19849(.O (g15787), .I1 (g12611), .I2 (g6519));
ND2X1 gate19850(.O (g15788), .I1 (g12657), .I2 (g6574));
ND2X1 gate19851(.O (g15789), .I1 (g12657), .I2 (g6783));
ND2X1 gate19852(.O (g15791), .I1 (g12711), .I2 (g7085));
ND2X1 gate19853(.O (g15803), .I1 (g13375), .I2 (g12354));
ND2X1 gate19854(.O (g15804), .I1 (g11660), .I2 (g12392));
ND2X1 gate19855(.O (g15805), .I1 (g12565), .I2 (g6232));
ND2X1 gate19856(.O (g15806), .I1 (g12565), .I2 (g6314));
ND2X1 gate19857(.O (g15807), .I1 (g12611), .I2 (g6369));
ND2X1 gate19858(.O (g15808), .I1 (g12611), .I2 (g6519));
ND2X1 gate19859(.O (g15809), .I1 (g12657), .I2 (g6574));
ND2X1 gate19860(.O (g15810), .I1 (g12657), .I2 (g6783));
ND2X1 gate19861(.O (g15811), .I1 (g12711), .I2 (g6838));
ND2X1 gate19862(.O (g15812), .I1 (g12711), .I2 (g7085));
ND2X1 gate19863(.O (I22062), .I1 (g12999), .I2 (g12988));
ND2X1 gate19864(.O (I22063), .I1 (g12999), .I2 (I22062));
ND2X1 gate19865(.O (I22064), .I1 (g12988), .I2 (I22062));
ND2X1 gate19866(.O (g15814), .I1 (I22063), .I2 (I22064));
ND2X1 gate19867(.O (g15818), .I1 (g13024), .I2 (g12354));
ND2X1 gate19868(.O (g15819), .I1 (g13286), .I2 (g12392));
ND2X1 gate19869(.O (g15820), .I1 (g12565), .I2 (g6232));
ND2X1 gate19870(.O (g15821), .I1 (g12565), .I2 (g6314));
ND2X1 gate19871(.O (g15822), .I1 (g12611), .I2 (g6369));
ND2X1 gate19872(.O (g15823), .I1 (g12611), .I2 (g6519));
ND2X1 gate19873(.O (g15824), .I1 (g12657), .I2 (g6574));
ND2X1 gate19874(.O (g15825), .I1 (g12657), .I2 (g6783));
ND2X1 gate19875(.O (g15826), .I1 (g12711), .I2 (g6838));
ND2X1 gate19876(.O (g15827), .I1 (g12711), .I2 (g7085));
ND2X1 gate19877(.O (g15830), .I1 (g13310), .I2 (g12392));
ND2X1 gate19878(.O (g15831), .I1 (g13313), .I2 (g12392));
ND2X1 gate19879(.O (g15832), .I1 (g12565), .I2 (g6232));
ND2X1 gate19880(.O (g15833), .I1 (g12565), .I2 (g6314));
ND2X1 gate19881(.O (g15834), .I1 (g12611), .I2 (g6369));
ND2X1 gate19882(.O (g15835), .I1 (g12611), .I2 (g6519));
ND2X1 gate19883(.O (g15836), .I1 (g12657), .I2 (g6574));
ND2X1 gate19884(.O (g15837), .I1 (g12657), .I2 (g6783));
ND2X1 gate19885(.O (g15838), .I1 (g12711), .I2 (g6838));
ND2X1 gate19886(.O (g15839), .I1 (g12711), .I2 (g7085));
ND2X1 gate19887(.O (g15841), .I1 (g13331), .I2 (g12392));
ND2X1 gate19888(.O (g15842), .I1 (g13332), .I2 (g12392));
ND2X1 gate19889(.O (g15843), .I1 (g12565), .I2 (g6314));
ND2X1 gate19890(.O (g15844), .I1 (g12565), .I2 (g6232));
ND2X1 gate19891(.O (g15845), .I1 (g12565), .I2 (g6314));
ND2X1 gate19892(.O (g15846), .I1 (g12611), .I2 (g6369));
ND2X1 gate19893(.O (g15847), .I1 (g12611), .I2 (g6519));
ND2X1 gate19894(.O (g15848), .I1 (g12657), .I2 (g6574));
ND2X1 gate19895(.O (g15849), .I1 (g12657), .I2 (g6783));
ND2X1 gate19896(.O (g15850), .I1 (g12711), .I2 (g6838));
ND2X1 gate19897(.O (g15851), .I1 (g12711), .I2 (g7085));
ND2X1 gate19898(.O (g15853), .I1 (g13310), .I2 (g12354));
ND2X1 gate19899(.O (g15854), .I1 (g13353), .I2 (g12392));
ND2X1 gate19900(.O (g15855), .I1 (g13354), .I2 (g12392));
ND2X1 gate19901(.O (g15856), .I1 (g12565), .I2 (g6232));
ND2X1 gate19902(.O (g15857), .I1 (g12565), .I2 (g6314));
ND2X1 gate19903(.O (g15858), .I1 (g12565), .I2 (g6232));
ND2X1 gate19904(.O (g15866), .I1 (g12611), .I2 (g6519));
ND2X1 gate19905(.O (g15867), .I1 (g12611), .I2 (g6369));
ND2X1 gate19906(.O (g15868), .I1 (g12611), .I2 (g6519));
ND2X1 gate19907(.O (g15869), .I1 (g12657), .I2 (g6574));
ND2X1 gate19908(.O (g15870), .I1 (g12657), .I2 (g6783));
ND2X1 gate19909(.O (g15871), .I1 (g12711), .I2 (g6838));
ND2X1 gate19910(.O (g15872), .I1 (g12711), .I2 (g7085));
ND2X1 gate19911(.O (g15877), .I1 (g13374), .I2 (g12392));
ND2X1 gate19912(.O (g15878), .I1 (g13375), .I2 (g12392));
ND2X1 gate19913(.O (g15879), .I1 (g12565), .I2 (g6232));
ND2X1 gate19914(.O (g15887), .I1 (g12611), .I2 (g6369));
ND2X1 gate19915(.O (g15888), .I1 (g12611), .I2 (g6519));
ND2X1 gate19916(.O (g15889), .I1 (g12611), .I2 (g6369));
ND2X1 gate19917(.O (g15897), .I1 (g12657), .I2 (g6783));
ND2X1 gate19918(.O (g15898), .I1 (g12657), .I2 (g6574));
ND2X1 gate19919(.O (g15899), .I1 (g12657), .I2 (g6783));
ND2X1 gate19920(.O (g15900), .I1 (g12711), .I2 (g6838));
ND2X1 gate19921(.O (g15901), .I1 (g12711), .I2 (g7085));
ND2X1 gate19922(.O (g15903), .I1 (g13404), .I2 (g12392));
ND2X1 gate19923(.O (g15912), .I1 (g12611), .I2 (g6369));
ND2X1 gate19924(.O (g15920), .I1 (g12657), .I2 (g6574));
ND2X1 gate19925(.O (g15921), .I1 (g12657), .I2 (g6783));
ND2X1 gate19926(.O (g15922), .I1 (g12657), .I2 (g6574));
ND2X1 gate19927(.O (g15930), .I1 (g12711), .I2 (g7085));
ND2X1 gate19928(.O (g15931), .I1 (g12711), .I2 (g6838));
ND2X1 gate19929(.O (g15932), .I1 (g12711), .I2 (g7085));
ND2X1 gate19930(.O (g15941), .I1 (g12657), .I2 (g6574));
ND2X1 gate19931(.O (g15949), .I1 (g12711), .I2 (g6838));
ND2X1 gate19932(.O (g15950), .I1 (g12711), .I2 (g7085));
ND2X1 gate19933(.O (g15951), .I1 (g12711), .I2 (g6838));
ND2X1 gate19934(.O (g15970), .I1 (g12711), .I2 (g6838));
ND2X1 gate19935(.O (g15990), .I1 (g12886), .I2 (g6912));
ND2X1 gate19936(.O (g15992), .I1 (g12886), .I2 (g6678));
ND2X1 gate19937(.O (g15993), .I1 (g12926), .I2 (g7162));
ND2X1 gate19938(.O (g15995), .I1 (g12926), .I2 (g6980));
ND2X1 gate19939(.O (g15996), .I1 (g12955), .I2 (g7358));
ND2X1 gate19940(.O (g15999), .I1 (g12955), .I2 (g7230));
ND2X1 gate19941(.O (g16000), .I1 (g12984), .I2 (g7488));
ND2X1 gate19942(.O (g16006), .I1 (g12984), .I2 (g7426));
ND2X1 gate19943(.O (g16085), .I1 (g12883), .I2 (g633));
ND2X1 gate19944(.O (g16123), .I1 (g12923), .I2 (g1319));
ND2X1 gate19945(.O (I22282), .I1 (g2962), .I2 (g13348));
ND2X1 gate19946(.O (I22283), .I1 (g2962), .I2 (I22282));
ND2X1 gate19947(.O (I22284), .I1 (g13348), .I2 (I22282));
ND2X1 gate19948(.O (g16132), .I1 (I22283), .I2 (I22284));
ND2X1 gate19949(.O (g16174), .I1 (g12952), .I2 (g2013));
ND2X1 gate19950(.O (I22316), .I1 (g2934), .I2 (g13370));
ND2X1 gate19951(.O (I22317), .I1 (g2934), .I2 (I22316));
ND2X1 gate19952(.O (I22318), .I1 (g13370), .I2 (I22316));
ND2X1 gate19953(.O (g16181), .I1 (I22317), .I2 (I22318));
ND2X1 gate19954(.O (g16233), .I1 (g12981), .I2 (g2707));
ND2X1 gate19955(.O (g16341), .I1 (g12377), .I2 (g12407));
ND2X1 gate19956(.O (g16412), .I1 (g12565), .I2 (g3254));
ND2X1 gate19957(.O (g16439), .I1 (g13082), .I2 (g2912));
ND2X1 gate19958(.O (g16442), .I1 (g12565), .I2 (g3254));
ND2X1 gate19959(.O (g16446), .I1 (g12611), .I2 (g3410));
ND2X1 gate19960(.O (g16463), .I1 (g13004), .I2 (g3018));
ND2X1 gate19961(.O (g16536), .I1 (g15873), .I2 (g2896));
ND2X1 gate19962(.O (I22630), .I1 (g13507), .I2 (g15978));
ND2X1 gate19963(.O (I22631), .I1 (g13507), .I2 (I22630));
ND2X1 gate19964(.O (I22632), .I1 (g15978), .I2 (I22630));
ND2X1 gate19965(.O (g16566), .I1 (I22631), .I2 (I22632));
ND2X1 gate19966(.O (I22705), .I1 (g13348), .I2 (g15661));
ND2X1 gate19967(.O (I22706), .I1 (g13348), .I2 (I22705));
ND2X1 gate19968(.O (I22707), .I1 (g15661), .I2 (I22705));
ND2X1 gate19969(.O (g16662), .I1 (I22706), .I2 (I22707));
ND2X1 gate19970(.O (I22884), .I1 (g13370), .I2 (g15661));
ND2X1 gate19971(.O (I22885), .I1 (g13370), .I2 (I22884));
ND2X1 gate19972(.O (I22886), .I1 (g15661), .I2 (I22884));
ND2X1 gate19973(.O (g16935), .I1 (I22885), .I2 (I22886));
ND2X1 gate19974(.O (I22900), .I1 (g15022), .I2 (g14000));
ND2X1 gate19975(.O (I22901), .I1 (g15022), .I2 (I22900));
ND2X1 gate19976(.O (I22902), .I1 (g14000), .I2 (I22900));
ND2X1 gate19977(.O (g16965), .I1 (I22901), .I2 (I22902));
ND2X1 gate19978(.O (I22917), .I1 (g15096), .I2 (g13945));
ND2X1 gate19979(.O (I22918), .I1 (g15096), .I2 (I22917));
ND2X1 gate19980(.O (I22919), .I1 (g13945), .I2 (I22917));
ND2X1 gate19981(.O (g16985), .I1 (I22918), .I2 (I22919));
ND2X1 gate19982(.O (I22924), .I1 (g15118), .I2 (g14091));
ND2X1 gate19983(.O (I22925), .I1 (g15118), .I2 (I22924));
ND2X1 gate19984(.O (I22926), .I1 (g14091), .I2 (I22924));
ND2X1 gate19985(.O (g16986), .I1 (I22925), .I2 (I22926));
ND2X1 gate19986(.O (I22936), .I1 (g9150), .I2 (g13906));
ND2X1 gate19987(.O (I22937), .I1 (g9150), .I2 (I22936));
ND2X1 gate19988(.O (I22938), .I1 (g13906), .I2 (I22936));
ND2X1 gate19989(.O (g16992), .I1 (I22937), .I2 (I22938));
ND2X1 gate19990(.O (I22945), .I1 (g15188), .I2 (g14015));
ND2X1 gate19991(.O (I22946), .I1 (g15188), .I2 (I22945));
ND2X1 gate19992(.O (I22947), .I1 (g14015), .I2 (I22945));
ND2X1 gate19993(.O (g16995), .I1 (I22946), .I2 (I22947));
ND2X1 gate19994(.O (I22952), .I1 (g15210), .I2 (g14206));
ND2X1 gate19995(.O (I22953), .I1 (g15210), .I2 (I22952));
ND2X1 gate19996(.O (I22954), .I1 (g14206), .I2 (I22952));
ND2X1 gate19997(.O (g16996), .I1 (I22953), .I2 (I22954));
ND2X1 gate19998(.O (I22962), .I1 (g9161), .I2 (g13885));
ND2X1 gate19999(.O (I22963), .I1 (g9161), .I2 (I22962));
ND2X1 gate20000(.O (I22964), .I1 (g13885), .I2 (I22962));
ND2X1 gate20001(.O (g17000), .I1 (I22963), .I2 (I22964));
ND2X1 gate20002(.O (I22972), .I1 (g9174), .I2 (g13962));
ND2X1 gate20003(.O (I22973), .I1 (g9174), .I2 (I22972));
ND2X1 gate20004(.O (I22974), .I1 (g13962), .I2 (I22972));
ND2X1 gate20005(.O (g17016), .I1 (I22973), .I2 (I22974));
ND2X1 gate20006(.O (I22981), .I1 (g15274), .I2 (g14106));
ND2X1 gate20007(.O (I22982), .I1 (g15274), .I2 (I22981));
ND2X1 gate20008(.O (I22983), .I1 (g14106), .I2 (I22981));
ND2X1 gate20009(.O (g17019), .I1 (I22982), .I2 (I22983));
ND2X1 gate20010(.O (I22988), .I1 (g15296), .I2 (g14321));
ND2X1 gate20011(.O (I22989), .I1 (g15296), .I2 (I22988));
ND2X1 gate20012(.O (I22990), .I1 (g14321), .I2 (I22988));
ND2X1 gate20013(.O (g17020), .I1 (I22989), .I2 (I22990));
ND2X1 gate20014(.O (I22998), .I1 (g9187), .I2 (g13872));
ND2X1 gate20015(.O (I22999), .I1 (g9187), .I2 (I22998));
ND2X1 gate20016(.O (I23000), .I1 (g13872), .I2 (I22998));
ND2X1 gate20017(.O (g17024), .I1 (I22999), .I2 (I23000));
ND2X1 gate20018(.O (I23008), .I1 (g9203), .I2 (g13926));
ND2X1 gate20019(.O (I23009), .I1 (g9203), .I2 (I23008));
ND2X1 gate20020(.O (I23010), .I1 (g13926), .I2 (I23008));
ND2X1 gate20021(.O (g17030), .I1 (I23009), .I2 (I23010));
ND2X1 gate20022(.O (I23018), .I1 (g9216), .I2 (g14032));
ND2X1 gate20023(.O (I23019), .I1 (g9216), .I2 (I23018));
ND2X1 gate20024(.O (I23020), .I1 (g14032), .I2 (I23018));
ND2X1 gate20025(.O (g17046), .I1 (I23019), .I2 (I23020));
ND2X1 gate20026(.O (I23027), .I1 (g15366), .I2 (g14221));
ND2X1 gate20027(.O (I23028), .I1 (g15366), .I2 (I23027));
ND2X1 gate20028(.O (I23029), .I1 (g14221), .I2 (I23027));
ND2X1 gate20029(.O (g17049), .I1 (I23028), .I2 (I23029));
ND2X1 gate20030(.O (I23034), .I1 (g9232), .I2 (g13864));
ND2X1 gate20031(.O (I23035), .I1 (g9232), .I2 (I23034));
ND2X1 gate20032(.O (I23036), .I1 (g13864), .I2 (I23034));
ND2X1 gate20033(.O (g17050), .I1 (I23035), .I2 (I23036));
ND2X1 gate20034(.O (I23045), .I1 (g9248), .I2 (g13894));
ND2X1 gate20035(.O (I23046), .I1 (g9248), .I2 (I23045));
ND2X1 gate20036(.O (I23047), .I1 (g13894), .I2 (I23045));
ND2X1 gate20037(.O (g17058), .I1 (I23046), .I2 (I23047));
ND2X1 gate20038(.O (I23055), .I1 (g9264), .I2 (g13982));
ND2X1 gate20039(.O (I23056), .I1 (g9264), .I2 (I23055));
ND2X1 gate20040(.O (I23057), .I1 (g13982), .I2 (I23055));
ND2X1 gate20041(.O (g17064), .I1 (I23056), .I2 (I23057));
ND2X1 gate20042(.O (I23065), .I1 (g9277), .I2 (g14123));
ND2X1 gate20043(.O (I23066), .I1 (g9277), .I2 (I23065));
ND2X1 gate20044(.O (I23067), .I1 (g14123), .I2 (I23065));
ND2X1 gate20045(.O (g17080), .I1 (I23066), .I2 (I23067));
ND2X1 gate20046(.O (I23074), .I1 (g9293), .I2 (g13856));
ND2X1 gate20047(.O (I23075), .I1 (g9293), .I2 (I23074));
ND2X1 gate20048(.O (I23076), .I1 (g13856), .I2 (I23074));
ND2X1 gate20049(.O (g17083), .I1 (I23075), .I2 (I23076));
ND2X1 gate20050(.O (I23082), .I1 (g9310), .I2 (g13879));
ND2X1 gate20051(.O (I23083), .I1 (g9310), .I2 (I23082));
ND2X1 gate20052(.O (I23084), .I1 (g13879), .I2 (I23082));
ND2X1 gate20053(.O (g17085), .I1 (I23083), .I2 (I23084));
ND2X1 gate20054(.O (I23093), .I1 (g9326), .I2 (g13935));
ND2X1 gate20055(.O (I23094), .I1 (g9326), .I2 (I23093));
ND2X1 gate20056(.O (I23095), .I1 (g13935), .I2 (I23093));
ND2X1 gate20057(.O (g17093), .I1 (I23094), .I2 (I23095));
ND2X1 gate20058(.O (I23103), .I1 (g9342), .I2 (g14052));
ND2X1 gate20059(.O (I23104), .I1 (g9342), .I2 (I23103));
ND2X1 gate20060(.O (I23105), .I1 (g14052), .I2 (I23103));
ND2X1 gate20061(.O (g17099), .I1 (I23104), .I2 (I23105));
ND2X1 gate20062(.O (I23113), .I1 (g9356), .I2 (g13848));
ND2X1 gate20063(.O (I23114), .I1 (g9356), .I2 (I23113));
ND2X1 gate20064(.O (I23115), .I1 (g13848), .I2 (I23113));
ND2X1 gate20065(.O (g17115), .I1 (I23114), .I2 (I23115));
ND2X1 gate20066(.O (g17118), .I1 (g13915), .I2 (g13893));
ND2X1 gate20067(.O (I23123), .I1 (g9374), .I2 (g13866));
ND2X1 gate20068(.O (I23124), .I1 (g9374), .I2 (I23123));
ND2X1 gate20069(.O (I23125), .I1 (g13866), .I2 (I23123));
ND2X1 gate20070(.O (g17121), .I1 (I23124), .I2 (I23125));
ND2X1 gate20071(.O (I23131), .I1 (g9391), .I2 (g13901));
ND2X1 gate20072(.O (I23132), .I1 (g9391), .I2 (I23131));
ND2X1 gate20073(.O (I23133), .I1 (g13901), .I2 (I23131));
ND2X1 gate20074(.O (g17123), .I1 (I23132), .I2 (I23133));
ND2X1 gate20075(.O (I23142), .I1 (g9407), .I2 (g13991));
ND2X1 gate20076(.O (I23143), .I1 (g9407), .I2 (I23142));
ND2X1 gate20077(.O (I23144), .I1 (g13991), .I2 (I23142));
ND2X1 gate20078(.O (g17131), .I1 (I23143), .I2 (I23144));
ND2X1 gate20079(.O (I23152), .I1 (g9427), .I2 (g14061));
ND2X1 gate20080(.O (I23153), .I1 (g9427), .I2 (I23152));
ND2X1 gate20081(.O (I23154), .I1 (g14061), .I2 (I23152));
ND2X1 gate20082(.O (g17137), .I1 (I23153), .I2 (I23154));
ND2X1 gate20083(.O (g17139), .I1 (g13957), .I2 (g13915));
ND2X1 gate20084(.O (I23161), .I1 (g9453), .I2 (g13857));
ND2X1 gate20085(.O (I23162), .I1 (g9453), .I2 (I23161));
ND2X1 gate20086(.O (I23163), .I1 (g13857), .I2 (I23161));
ND2X1 gate20087(.O (g17142), .I1 (I23162), .I2 (I23163));
ND2X1 gate20088(.O (g17145), .I1 (g13971), .I2 (g13934));
ND2X1 gate20089(.O (I23171), .I1 (g9471), .I2 (g13881));
ND2X1 gate20090(.O (I23172), .I1 (g9471), .I2 (I23171));
ND2X1 gate20091(.O (I23173), .I1 (g13881), .I2 (I23171));
ND2X1 gate20092(.O (g17148), .I1 (I23172), .I2 (I23173));
ND2X1 gate20093(.O (I23179), .I1 (g9488), .I2 (g13942));
ND2X1 gate20094(.O (I23180), .I1 (g9488), .I2 (I23179));
ND2X1 gate20095(.O (I23181), .I1 (g13942), .I2 (I23179));
ND2X1 gate20096(.O (g17150), .I1 (I23180), .I2 (I23181));
ND2X1 gate20097(.O (I23190), .I1 (g9507), .I2 (g13999));
ND2X1 gate20098(.O (I23191), .I1 (g9507), .I2 (I23190));
ND2X1 gate20099(.O (I23192), .I1 (g13999), .I2 (I23190));
ND2X1 gate20100(.O (g17158), .I1 (I23191), .I2 (I23192));
ND2X1 gate20101(.O (g17159), .I1 (g14642), .I2 (g14657));
ND2X1 gate20102(.O (I23198), .I1 (g9569), .I2 (g14176));
ND2X1 gate20103(.O (I23199), .I1 (g9569), .I2 (I23198));
ND2X1 gate20104(.O (I23200), .I1 (g14176), .I2 (I23198));
ND2X1 gate20105(.O (g17160), .I1 (I23199), .I2 (I23200));
ND2X1 gate20106(.O (g17162), .I1 (g14027), .I2 (g13971));
ND2X1 gate20107(.O (I23207), .I1 (g9595), .I2 (g13867));
ND2X1 gate20108(.O (I23208), .I1 (g9595), .I2 (I23207));
ND2X1 gate20109(.O (I23209), .I1 (g13867), .I2 (I23207));
ND2X1 gate20110(.O (g17165), .I1 (I23208), .I2 (I23209));
ND2X1 gate20111(.O (g17168), .I1 (g14041), .I2 (g13990));
ND2X1 gate20112(.O (I23217), .I1 (g9613), .I2 (g13903));
ND2X1 gate20113(.O (I23218), .I1 (g9613), .I2 (I23217));
ND2X1 gate20114(.O (I23219), .I1 (g13903), .I2 (I23217));
ND2X1 gate20115(.O (g17171), .I1 (I23218), .I2 (I23219));
ND2X1 gate20116(.O (I23225), .I1 (g9649), .I2 (g14090));
ND2X1 gate20117(.O (I23226), .I1 (g9649), .I2 (I23225));
ND2X1 gate20118(.O (I23227), .I1 (g14090), .I2 (I23225));
ND2X1 gate20119(.O (g17173), .I1 (I23226), .I2 (I23227));
ND2X1 gate20120(.O (g17174), .I1 (g14669), .I2 (g14691));
ND2X1 gate20121(.O (I23233), .I1 (g9711), .I2 (g14291));
ND2X1 gate20122(.O (I23234), .I1 (g9711), .I2 (I23233));
ND2X1 gate20123(.O (I23235), .I1 (g14291), .I2 (I23233));
ND2X1 gate20124(.O (g17175), .I1 (I23234), .I2 (I23235));
ND2X1 gate20125(.O (g17177), .I1 (g14118), .I2 (g14041));
ND2X1 gate20126(.O (I23242), .I1 (g9737), .I2 (g13882));
ND2X1 gate20127(.O (I23243), .I1 (g9737), .I2 (I23242));
ND2X1 gate20128(.O (I23244), .I1 (g13882), .I2 (I23242));
ND2X1 gate20129(.O (g17180), .I1 (I23243), .I2 (I23244));
ND2X1 gate20130(.O (g17183), .I1 (g14132), .I2 (g14060));
ND2X1 gate20131(.O (I23256), .I1 (g9795), .I2 (g14205));
ND2X1 gate20132(.O (I23257), .I1 (g9795), .I2 (I23256));
ND2X1 gate20133(.O (I23258), .I1 (g14205), .I2 (I23256));
ND2X1 gate20134(.O (g17190), .I1 (I23257), .I2 (I23258));
ND2X1 gate20135(.O (g17191), .I1 (g14703), .I2 (g14725));
ND2X1 gate20136(.O (I23264), .I1 (g9857), .I2 (g14413));
ND2X1 gate20137(.O (I23265), .I1 (g9857), .I2 (I23264));
ND2X1 gate20138(.O (I23266), .I1 (g14413), .I2 (I23264));
ND2X1 gate20139(.O (g17192), .I1 (I23265), .I2 (I23266));
ND2X1 gate20140(.O (g17194), .I1 (g14233), .I2 (g14132));
ND2X1 gate20141(.O (I23277), .I1 (g9941), .I2 (g14320));
ND2X1 gate20142(.O (I23278), .I1 (g9941), .I2 (I23277));
ND2X1 gate20143(.O (I23279), .I1 (g14320), .I2 (I23277));
ND2X1 gate20144(.O (g17201), .I1 (I23278), .I2 (I23279));
ND2X1 gate20145(.O (g17202), .I1 (g14737), .I2 (g14753));
ND2X1 gate20146(.O (I23806), .I1 (g14062), .I2 (g9150));
ND2X1 gate20147(.O (I23807), .I1 (g14062), .I2 (I23806));
ND2X1 gate20148(.O (I23808), .I1 (g9150), .I2 (I23806));
ND2X1 gate20149(.O (g17729), .I1 (I23807), .I2 (I23808));
ND2X1 gate20150(.O (I23878), .I1 (g14001), .I2 (g9187));
ND2X1 gate20151(.O (I23879), .I1 (g14001), .I2 (I23878));
ND2X1 gate20152(.O (I23880), .I1 (g9187), .I2 (I23878));
ND2X1 gate20153(.O (g17807), .I1 (I23879), .I2 (I23880));
ND2X1 gate20154(.O (I23893), .I1 (g14177), .I2 (g9174));
ND2X1 gate20155(.O (I23894), .I1 (g14177), .I2 (I23893));
ND2X1 gate20156(.O (I23895), .I1 (g9174), .I2 (I23893));
ND2X1 gate20157(.O (g17830), .I1 (I23894), .I2 (I23895));
ND2X1 gate20158(.O (I23941), .I1 (g13946), .I2 (g9293));
ND2X1 gate20159(.O (I23942), .I1 (g13946), .I2 (I23941));
ND2X1 gate20160(.O (I23943), .I1 (g9293), .I2 (I23941));
ND2X1 gate20161(.O (g17887), .I1 (I23942), .I2 (I23943));
ND2X1 gate20162(.O (I23958), .I1 (g6513), .I2 (g14171));
ND2X1 gate20163(.O (I23959), .I1 (g6513), .I2 (I23958));
ND2X1 gate20164(.O (I23960), .I1 (g14171), .I2 (I23958));
ND2X1 gate20165(.O (g17913), .I1 (I23959), .I2 (I23960));
ND2X1 gate20166(.O (I23966), .I1 (g14092), .I2 (g9248));
ND2X1 gate20167(.O (I23967), .I1 (g14092), .I2 (I23966));
ND2X1 gate20168(.O (I23968), .I1 (g9248), .I2 (I23966));
ND2X1 gate20169(.O (g17919), .I1 (I23967), .I2 (I23968));
ND2X1 gate20170(.O (I23981), .I1 (g14292), .I2 (g9216));
ND2X1 gate20171(.O (I23982), .I1 (g14292), .I2 (I23981));
ND2X1 gate20172(.O (I23983), .I1 (g9216), .I2 (I23981));
ND2X1 gate20173(.O (g17942), .I1 (I23982), .I2 (I23983));
ND2X1 gate20174(.O (I24005), .I1 (g7548), .I2 (g15814));
ND2X1 gate20175(.O (I24006), .I1 (g7548), .I2 (I24005));
ND2X1 gate20176(.O (I24007), .I1 (g15814), .I2 (I24005));
ND2X1 gate20177(.O (g17968), .I1 (I24006), .I2 (I24007));
ND2X1 gate20178(.O (I24015), .I1 (g13907), .I2 (g9427));
ND2X1 gate20179(.O (I24016), .I1 (g13907), .I2 (I24015));
ND2X1 gate20180(.O (I24017), .I1 (g9427), .I2 (I24015));
ND2X1 gate20181(.O (g17979), .I1 (I24016), .I2 (I24017));
ND2X1 gate20182(.O (g17985), .I1 (g14641), .I2 (g9636));
ND2X1 gate20183(.O (I24028), .I1 (g6201), .I2 (g14086));
ND2X1 gate20184(.O (I24029), .I1 (g6201), .I2 (I24028));
ND2X1 gate20185(.O (I24030), .I1 (g14086), .I2 (I24028));
ND2X1 gate20186(.O (g17992), .I1 (I24029), .I2 (I24030));
ND2X1 gate20187(.O (I24036), .I1 (g14016), .I2 (g9374));
ND2X1 gate20188(.O (I24037), .I1 (g14016), .I2 (I24036));
ND2X1 gate20189(.O (I24038), .I1 (g9374), .I2 (I24036));
ND2X1 gate20190(.O (g17998), .I1 (I24037), .I2 (I24038));
ND2X1 gate20191(.O (I24053), .I1 (g6777), .I2 (g14286));
ND2X1 gate20192(.O (I24054), .I1 (g6777), .I2 (I24053));
ND2X1 gate20193(.O (I24055), .I1 (g14286), .I2 (I24053));
ND2X1 gate20194(.O (g18024), .I1 (I24054), .I2 (I24055));
ND2X1 gate20195(.O (I24061), .I1 (g14207), .I2 (g9326));
ND2X1 gate20196(.O (I24062), .I1 (g14207), .I2 (I24061));
ND2X1 gate20197(.O (I24063), .I1 (g9326), .I2 (I24061));
ND2X1 gate20198(.O (g18030), .I1 (I24062), .I2 (I24063));
ND2X1 gate20199(.O (I24076), .I1 (g14414), .I2 (g9277));
ND2X1 gate20200(.O (I24077), .I1 (g14414), .I2 (I24076));
ND2X1 gate20201(.O (I24078), .I1 (g9277), .I2 (I24076));
ND2X1 gate20202(.O (g18053), .I1 (I24077), .I2 (I24078));
ND2X1 gate20203(.O (I24091), .I1 (g13886), .I2 (g15096));
ND2X1 gate20204(.O (I24092), .I1 (g13886), .I2 (I24091));
ND2X1 gate20205(.O (I24093), .I1 (g15096), .I2 (I24091));
ND2X1 gate20206(.O (g18079), .I1 (I24092), .I2 (I24093));
ND2X1 gate20207(.O (I24102), .I1 (g6363), .I2 (g14011));
ND2X1 gate20208(.O (I24103), .I1 (g6363), .I2 (I24102));
ND2X1 gate20209(.O (I24104), .I1 (g14011), .I2 (I24102));
ND2X1 gate20210(.O (g18090), .I1 (I24103), .I2 (I24104));
ND2X1 gate20211(.O (I24110), .I1 (g13963), .I2 (g9569));
ND2X1 gate20212(.O (I24111), .I1 (g13963), .I2 (I24110));
ND2X1 gate20213(.O (I24112), .I1 (g9569), .I2 (I24110));
ND2X1 gate20214(.O (g18096), .I1 (I24111), .I2 (I24112));
ND2X1 gate20215(.O (g18102), .I1 (g14668), .I2 (g9782));
ND2X1 gate20216(.O (I24123), .I1 (g6290), .I2 (g14201));
ND2X1 gate20217(.O (I24124), .I1 (g6290), .I2 (I24123));
ND2X1 gate20218(.O (I24125), .I1 (g14201), .I2 (I24123));
ND2X1 gate20219(.O (g18109), .I1 (I24124), .I2 (I24125));
ND2X1 gate20220(.O (I24131), .I1 (g14107), .I2 (g9471));
ND2X1 gate20221(.O (I24132), .I1 (g14107), .I2 (I24131));
ND2X1 gate20222(.O (I24133), .I1 (g9471), .I2 (I24131));
ND2X1 gate20223(.O (g18115), .I1 (I24132), .I2 (I24133));
ND2X1 gate20224(.O (I24148), .I1 (g7079), .I2 (g14408));
ND2X1 gate20225(.O (I24149), .I1 (g7079), .I2 (I24148));
ND2X1 gate20226(.O (I24150), .I1 (g14408), .I2 (I24148));
ND2X1 gate20227(.O (g18141), .I1 (I24149), .I2 (I24150));
ND2X1 gate20228(.O (I24156), .I1 (g14322), .I2 (g9407));
ND2X1 gate20229(.O (I24157), .I1 (g14322), .I2 (I24156));
ND2X1 gate20230(.O (I24158), .I1 (g9407), .I2 (I24156));
ND2X1 gate20231(.O (g18147), .I1 (I24157), .I2 (I24158));
ND2X1 gate20232(.O (I24178), .I1 (g13873), .I2 (g9161));
ND2X1 gate20233(.O (I24179), .I1 (g13873), .I2 (I24178));
ND2X1 gate20234(.O (I24180), .I1 (g9161), .I2 (I24178));
ND2X1 gate20235(.O (g18183), .I1 (I24179), .I2 (I24180));
ND2X1 gate20236(.O (I24186), .I1 (g6177), .I2 (g13958));
ND2X1 gate20237(.O (I24187), .I1 (g6177), .I2 (I24186));
ND2X1 gate20238(.O (I24188), .I1 (g13958), .I2 (I24186));
ND2X1 gate20239(.O (g18189), .I1 (I24187), .I2 (I24188));
ND2X1 gate20240(.O (I24194), .I1 (g13927), .I2 (g15188));
ND2X1 gate20241(.O (I24195), .I1 (g13927), .I2 (I24194));
ND2X1 gate20242(.O (I24196), .I1 (g15188), .I2 (I24194));
ND2X1 gate20243(.O (g18195), .I1 (I24195), .I2 (I24196));
ND2X1 gate20244(.O (I24205), .I1 (g6568), .I2 (g14102));
ND2X1 gate20245(.O (I24206), .I1 (g6568), .I2 (I24205));
ND2X1 gate20246(.O (I24207), .I1 (g14102), .I2 (I24205));
ND2X1 gate20247(.O (g18206), .I1 (I24206), .I2 (I24207));
ND2X1 gate20248(.O (I24213), .I1 (g14033), .I2 (g9711));
ND2X1 gate20249(.O (I24214), .I1 (g14033), .I2 (I24213));
ND2X1 gate20250(.O (I24215), .I1 (g9711), .I2 (I24213));
ND2X1 gate20251(.O (g18212), .I1 (I24214), .I2 (I24215));
ND2X1 gate20252(.O (g18218), .I1 (g14702), .I2 (g9928));
ND2X1 gate20253(.O (I24226), .I1 (g6427), .I2 (g14316));
ND2X1 gate20254(.O (I24227), .I1 (g6427), .I2 (I24226));
ND2X1 gate20255(.O (I24228), .I1 (g14316), .I2 (I24226));
ND2X1 gate20256(.O (g18225), .I1 (I24227), .I2 (I24228));
ND2X1 gate20257(.O (I24234), .I1 (g14222), .I2 (g9613));
ND2X1 gate20258(.O (I24235), .I1 (g14222), .I2 (I24234));
ND2X1 gate20259(.O (I24236), .I1 (g9613), .I2 (I24234));
ND2X1 gate20260(.O (g18231), .I1 (I24235), .I2 (I24236));
ND2X1 gate20261(.O (I24251), .I1 (g7329), .I2 (g14520));
ND2X1 gate20262(.O (I24252), .I1 (g7329), .I2 (I24251));
ND2X1 gate20263(.O (I24253), .I1 (g14520), .I2 (I24251));
ND2X1 gate20264(.O (g18257), .I1 (I24252), .I2 (I24253));
ND2X1 gate20265(.O (I24263), .I1 (g14342), .I2 (g9232));
ND2X1 gate20266(.O (I24264), .I1 (g14342), .I2 (I24263));
ND2X1 gate20267(.O (I24265), .I1 (g9232), .I2 (I24263));
ND2X1 gate20268(.O (g18270), .I1 (I24264), .I2 (I24265));
ND2X1 gate20269(.O (I24271), .I1 (g6180), .I2 (g13922));
ND2X1 gate20270(.O (I24272), .I1 (g6180), .I2 (I24271));
ND2X1 gate20271(.O (I24273), .I1 (g13922), .I2 (I24271));
ND2X1 gate20272(.O (g18276), .I1 (I24272), .I2 (I24273));
ND2X1 gate20273(.O (I24278), .I1 (g6284), .I2 (g13918));
ND2X1 gate20274(.O (I24279), .I1 (g6284), .I2 (I24278));
ND2X1 gate20275(.O (I24280), .I1 (g13918), .I2 (I24278));
ND2X1 gate20276(.O (g18277), .I1 (I24279), .I2 (I24280));
ND2X1 gate20277(.O (I24290), .I1 (g13895), .I2 (g9203));
ND2X1 gate20278(.O (I24291), .I1 (g13895), .I2 (I24290));
ND2X1 gate20279(.O (I24292), .I1 (g9203), .I2 (I24290));
ND2X1 gate20280(.O (g18290), .I1 (I24291), .I2 (I24292));
ND2X1 gate20281(.O (I24298), .I1 (g6209), .I2 (g14028));
ND2X1 gate20282(.O (I24299), .I1 (g6209), .I2 (I24298));
ND2X1 gate20283(.O (I24300), .I1 (g14028), .I2 (I24298));
ND2X1 gate20284(.O (g18296), .I1 (I24299), .I2 (I24300));
ND2X1 gate20285(.O (I24306), .I1 (g13983), .I2 (g15274));
ND2X1 gate20286(.O (I24307), .I1 (g13983), .I2 (I24306));
ND2X1 gate20287(.O (I24308), .I1 (g15274), .I2 (I24306));
ND2X1 gate20288(.O (g18302), .I1 (I24307), .I2 (I24308));
ND2X1 gate20289(.O (I24317), .I1 (g6832), .I2 (g14217));
ND2X1 gate20290(.O (I24318), .I1 (g6832), .I2 (I24317));
ND2X1 gate20291(.O (I24319), .I1 (g14217), .I2 (I24317));
ND2X1 gate20292(.O (g18313), .I1 (I24318), .I2 (I24319));
ND2X1 gate20293(.O (I24325), .I1 (g14124), .I2 (g9857));
ND2X1 gate20294(.O (I24326), .I1 (g14124), .I2 (I24325));
ND2X1 gate20295(.O (I24327), .I1 (g9857), .I2 (I24325));
ND2X1 gate20296(.O (g18319), .I1 (I24326), .I2 (I24327));
ND2X1 gate20297(.O (g18325), .I1 (g14736), .I2 (g10082));
ND2X1 gate20298(.O (I24338), .I1 (g6632), .I2 (g14438));
ND2X1 gate20299(.O (I24339), .I1 (g6632), .I2 (I24338));
ND2X1 gate20300(.O (I24340), .I1 (g14438), .I2 (I24338));
ND2X1 gate20301(.O (g18332), .I1 (I24339), .I2 (I24340));
ND2X1 gate20302(.O (I24351), .I1 (g14238), .I2 (g9356));
ND2X1 gate20303(.O (I24352), .I1 (g14238), .I2 (I24351));
ND2X1 gate20304(.O (I24353), .I1 (g9356), .I2 (I24351));
ND2X1 gate20305(.O (g18346), .I1 (I24352), .I2 (I24353));
ND2X1 gate20306(.O (I24361), .I1 (g6157), .I2 (g14525));
ND2X1 gate20307(.O (I24362), .I1 (g6157), .I2 (I24361));
ND2X1 gate20308(.O (I24363), .I1 (g14525), .I2 (I24361));
ND2X1 gate20309(.O (g18354), .I1 (I24362), .I2 (I24363));
ND2X1 gate20310(.O (I24372), .I1 (g14454), .I2 (g9310));
ND2X1 gate20311(.O (I24373), .I1 (g14454), .I2 (I24372));
ND2X1 gate20312(.O (I24374), .I1 (g9310), .I2 (I24372));
ND2X1 gate20313(.O (g18363), .I1 (I24373), .I2 (I24374));
ND2X1 gate20314(.O (I24380), .I1 (g6212), .I2 (g13978));
ND2X1 gate20315(.O (I24381), .I1 (g6212), .I2 (I24380));
ND2X1 gate20316(.O (I24382), .I1 (g13978), .I2 (I24380));
ND2X1 gate20317(.O (g18369), .I1 (I24381), .I2 (I24382));
ND2X1 gate20318(.O (I24387), .I1 (g6421), .I2 (g13974));
ND2X1 gate20319(.O (I24388), .I1 (g6421), .I2 (I24387));
ND2X1 gate20320(.O (I24389), .I1 (g13974), .I2 (I24387));
ND2X1 gate20321(.O (g18370), .I1 (I24388), .I2 (I24389));
ND2X1 gate20322(.O (I24399), .I1 (g13936), .I2 (g9264));
ND2X1 gate20323(.O (I24400), .I1 (g13936), .I2 (I24399));
ND2X1 gate20324(.O (I24401), .I1 (g9264), .I2 (I24399));
ND2X1 gate20325(.O (g18383), .I1 (I24400), .I2 (I24401));
ND2X1 gate20326(.O (I24407), .I1 (g6298), .I2 (g14119));
ND2X1 gate20327(.O (I24408), .I1 (g6298), .I2 (I24407));
ND2X1 gate20328(.O (I24409), .I1 (g14119), .I2 (I24407));
ND2X1 gate20329(.O (g18389), .I1 (I24408), .I2 (I24409));
ND2X1 gate20330(.O (I24415), .I1 (g14053), .I2 (g15366));
ND2X1 gate20331(.O (I24416), .I1 (g14053), .I2 (I24415));
ND2X1 gate20332(.O (I24417), .I1 (g15366), .I2 (I24415));
ND2X1 gate20333(.O (g18395), .I1 (I24416), .I2 (I24417));
ND2X1 gate20334(.O (I24426), .I1 (g7134), .I2 (g14332));
ND2X1 gate20335(.O (I24427), .I1 (g7134), .I2 (I24426));
ND2X1 gate20336(.O (I24428), .I1 (g14332), .I2 (I24426));
ND2X1 gate20337(.O (g18406), .I1 (I24427), .I2 (I24428));
ND2X1 gate20338(.O (I24436), .I1 (g14153), .I2 (g15022));
ND2X1 gate20339(.O (I24437), .I1 (g14153), .I2 (I24436));
ND2X1 gate20340(.O (I24438), .I1 (g15022), .I2 (I24436));
ND2X1 gate20341(.O (g18419), .I1 (I24437), .I2 (I24438));
ND2X1 gate20342(.O (I24443), .I1 (g14148), .I2 (g9507));
ND2X1 gate20343(.O (I24444), .I1 (g14148), .I2 (I24443));
ND2X1 gate20344(.O (I24445), .I1 (g9507), .I2 (I24443));
ND2X1 gate20345(.O (g18424), .I1 (I24444), .I2 (I24445));
ND2X1 gate20346(.O (I24452), .I1 (g6142), .I2 (g14450));
ND2X1 gate20347(.O (I24453), .I1 (g6142), .I2 (I24452));
ND2X1 gate20348(.O (I24454), .I1 (g14450), .I2 (I24452));
ND2X1 gate20349(.O (g18431), .I1 (I24453), .I2 (I24454));
ND2X1 gate20350(.O (I24464), .I1 (g14360), .I2 (g9453));
ND2X1 gate20351(.O (I24465), .I1 (g14360), .I2 (I24464));
ND2X1 gate20352(.O (I24466), .I1 (g9453), .I2 (I24464));
ND2X1 gate20353(.O (g18441), .I1 (I24465), .I2 (I24466));
ND2X1 gate20354(.O (I24474), .I1 (g6184), .I2 (g14580));
ND2X1 gate20355(.O (I24475), .I1 (g6184), .I2 (I24474));
ND2X1 gate20356(.O (I24476), .I1 (g14580), .I2 (I24474));
ND2X1 gate20357(.O (g18449), .I1 (I24475), .I2 (I24476));
ND2X1 gate20358(.O (I24485), .I1 (g14541), .I2 (g9391));
ND2X1 gate20359(.O (I24486), .I1 (g14541), .I2 (I24485));
ND2X1 gate20360(.O (I24487), .I1 (g9391), .I2 (I24485));
ND2X1 gate20361(.O (g18458), .I1 (I24486), .I2 (I24487));
ND2X1 gate20362(.O (I24493), .I1 (g6301), .I2 (g14048));
ND2X1 gate20363(.O (I24494), .I1 (g6301), .I2 (I24493));
ND2X1 gate20364(.O (I24495), .I1 (g14048), .I2 (I24493));
ND2X1 gate20365(.O (g18464), .I1 (I24494), .I2 (I24495));
ND2X1 gate20366(.O (I24500), .I1 (g6626), .I2 (g14044));
ND2X1 gate20367(.O (I24501), .I1 (g6626), .I2 (I24500));
ND2X1 gate20368(.O (I24502), .I1 (g14044), .I2 (I24500));
ND2X1 gate20369(.O (g18465), .I1 (I24501), .I2 (I24502));
ND2X1 gate20370(.O (I24512), .I1 (g13992), .I2 (g9342));
ND2X1 gate20371(.O (I24513), .I1 (g13992), .I2 (I24512));
ND2X1 gate20372(.O (I24514), .I1 (g9342), .I2 (I24512));
ND2X1 gate20373(.O (g18478), .I1 (I24513), .I2 (I24514));
ND2X1 gate20374(.O (I24520), .I1 (g6435), .I2 (g14234));
ND2X1 gate20375(.O (I24521), .I1 (g6435), .I2 (I24520));
ND2X1 gate20376(.O (I24522), .I1 (g14234), .I2 (I24520));
ND2X1 gate20377(.O (g18484), .I1 (I24521), .I2 (I24522));
ND2X1 gate20378(.O (I24530), .I1 (g6707), .I2 (g14355));
ND2X1 gate20379(.O (I24531), .I1 (g6707), .I2 (I24530));
ND2X1 gate20380(.O (I24532), .I1 (g14355), .I2 (I24530));
ND2X1 gate20381(.O (g18491), .I1 (I24531), .I2 (I24532));
ND2X1 gate20382(.O (I24537), .I1 (g14268), .I2 (g15118));
ND2X1 gate20383(.O (I24538), .I1 (g14268), .I2 (I24537));
ND2X1 gate20384(.O (I24539), .I1 (g15118), .I2 (I24537));
ND2X1 gate20385(.O (g18492), .I1 (I24538), .I2 (I24539));
ND2X1 gate20386(.O (I24544), .I1 (g14263), .I2 (g9649));
ND2X1 gate20387(.O (I24545), .I1 (g14263), .I2 (I24544));
ND2X1 gate20388(.O (I24546), .I1 (g9649), .I2 (I24544));
ND2X1 gate20389(.O (g18497), .I1 (I24545), .I2 (I24546));
ND2X1 gate20390(.O (I24553), .I1 (g6163), .I2 (g14537));
ND2X1 gate20391(.O (I24554), .I1 (g6163), .I2 (I24553));
ND2X1 gate20392(.O (I24555), .I1 (g14537), .I2 (I24553));
ND2X1 gate20393(.O (g18504), .I1 (I24554), .I2 (I24555));
ND2X1 gate20394(.O (I24565), .I1 (g14472), .I2 (g9595));
ND2X1 gate20395(.O (I24566), .I1 (g14472), .I2 (I24565));
ND2X1 gate20396(.O (I24567), .I1 (g9595), .I2 (I24565));
ND2X1 gate20397(.O (g18514), .I1 (I24566), .I2 (I24567));
ND2X1 gate20398(.O (I24575), .I1 (g6216), .I2 (g14614));
ND2X1 gate20399(.O (I24576), .I1 (g6216), .I2 (I24575));
ND2X1 gate20400(.O (I24577), .I1 (g14614), .I2 (I24575));
ND2X1 gate20401(.O (g18522), .I1 (I24576), .I2 (I24577));
ND2X1 gate20402(.O (I24586), .I1 (g14596), .I2 (g9488));
ND2X1 gate20403(.O (I24587), .I1 (g14596), .I2 (I24586));
ND2X1 gate20404(.O (I24588), .I1 (g9488), .I2 (I24586));
ND2X1 gate20405(.O (g18531), .I1 (I24587), .I2 (I24588));
ND2X1 gate20406(.O (I24594), .I1 (g6438), .I2 (g14139));
ND2X1 gate20407(.O (I24595), .I1 (g6438), .I2 (I24594));
ND2X1 gate20408(.O (I24596), .I1 (g14139), .I2 (I24594));
ND2X1 gate20409(.O (g18537), .I1 (I24595), .I2 (I24596));
ND2X1 gate20410(.O (I24601), .I1 (g6890), .I2 (g14135));
ND2X1 gate20411(.O (I24602), .I1 (g6890), .I2 (I24601));
ND2X1 gate20412(.O (I24603), .I1 (g14135), .I2 (I24601));
ND2X1 gate20413(.O (g18538), .I1 (I24602), .I2 (I24603));
ND2X1 gate20414(.O (I24611), .I1 (g15814), .I2 (g15978));
ND2X1 gate20415(.O (I24612), .I1 (g15814), .I2 (I24611));
ND2X1 gate20416(.O (I24613), .I1 (g15978), .I2 (I24611));
ND2X1 gate20417(.O (g18542), .I1 (I24612), .I2 (I24613));
ND2X1 gate20418(.O (I24624), .I1 (g6136), .I2 (g14252));
ND2X1 gate20419(.O (I24625), .I1 (g6136), .I2 (I24624));
ND2X1 gate20420(.O (I24626), .I1 (g14252), .I2 (I24624));
ND2X1 gate20421(.O (g18553), .I1 (I24625), .I2 (I24626));
ND2X1 gate20422(.O (I24632), .I1 (g7009), .I2 (g14467));
ND2X1 gate20423(.O (I24633), .I1 (g7009), .I2 (I24632));
ND2X1 gate20424(.O (I24634), .I1 (g14467), .I2 (I24632));
ND2X1 gate20425(.O (g18555), .I1 (I24633), .I2 (I24634));
ND2X1 gate20426(.O (I24639), .I1 (g14390), .I2 (g15210));
ND2X1 gate20427(.O (I24640), .I1 (g14390), .I2 (I24639));
ND2X1 gate20428(.O (I24641), .I1 (g15210), .I2 (I24639));
ND2X1 gate20429(.O (g18556), .I1 (I24640), .I2 (I24641));
ND2X1 gate20430(.O (I24646), .I1 (g14385), .I2 (g9795));
ND2X1 gate20431(.O (I24647), .I1 (g14385), .I2 (I24646));
ND2X1 gate20432(.O (I24648), .I1 (g9795), .I2 (I24646));
ND2X1 gate20433(.O (g18561), .I1 (I24647), .I2 (I24648));
ND2X1 gate20434(.O (I24655), .I1 (g6190), .I2 (g14592));
ND2X1 gate20435(.O (I24656), .I1 (g6190), .I2 (I24655));
ND2X1 gate20436(.O (I24657), .I1 (g14592), .I2 (I24655));
ND2X1 gate20437(.O (g18568), .I1 (I24656), .I2 (I24657));
ND2X1 gate20438(.O (I24667), .I1 (g14559), .I2 (g9737));
ND2X1 gate20439(.O (I24668), .I1 (g14559), .I2 (I24667));
ND2X1 gate20440(.O (I24669), .I1 (g9737), .I2 (I24667));
ND2X1 gate20441(.O (g18578), .I1 (I24668), .I2 (I24669));
ND2X1 gate20442(.O (I24677), .I1 (g6305), .I2 (g14637));
ND2X1 gate20443(.O (I24678), .I1 (g6305), .I2 (I24677));
ND2X1 gate20444(.O (I24679), .I1 (g14637), .I2 (I24677));
ND2X1 gate20445(.O (g18586), .I1 (I24678), .I2 (I24679));
ND2X1 gate20446(.O (I24694), .I1 (g6146), .I2 (g14374));
ND2X1 gate20447(.O (I24695), .I1 (g6146), .I2 (I24694));
ND2X1 gate20448(.O (I24696), .I1 (g14374), .I2 (I24694));
ND2X1 gate20449(.O (g18603), .I1 (I24695), .I2 (I24696));
ND2X1 gate20450(.O (I24702), .I1 (g7259), .I2 (g14554));
ND2X1 gate20451(.O (I24703), .I1 (g7259), .I2 (I24702));
ND2X1 gate20452(.O (I24704), .I1 (g14554), .I2 (I24702));
ND2X1 gate20453(.O (g18605), .I1 (I24703), .I2 (I24704));
ND2X1 gate20454(.O (I24709), .I1 (g14502), .I2 (g15296));
ND2X1 gate20455(.O (I24710), .I1 (g14502), .I2 (I24709));
ND2X1 gate20456(.O (I24711), .I1 (g15296), .I2 (I24709));
ND2X1 gate20457(.O (g18606), .I1 (I24710), .I2 (I24711));
ND2X1 gate20458(.O (I24716), .I1 (g14497), .I2 (g9941));
ND2X1 gate20459(.O (I24717), .I1 (g14497), .I2 (I24716));
ND2X1 gate20460(.O (I24718), .I1 (g9941), .I2 (I24716));
ND2X1 gate20461(.O (g18611), .I1 (I24717), .I2 (I24718));
ND2X1 gate20462(.O (I24725), .I1 (g6222), .I2 (g14626));
ND2X1 gate20463(.O (I24726), .I1 (g6222), .I2 (I24725));
ND2X1 gate20464(.O (I24727), .I1 (g14626), .I2 (I24725));
ND2X1 gate20465(.O (g18618), .I1 (I24726), .I2 (I24727));
ND2X1 gate20466(.O (I24743), .I1 (g6167), .I2 (g14486));
ND2X1 gate20467(.O (I24744), .I1 (g6167), .I2 (I24743));
ND2X1 gate20468(.O (I24745), .I1 (g14486), .I2 (I24743));
ND2X1 gate20469(.O (g18635), .I1 (I24744), .I2 (I24745));
ND2X1 gate20470(.O (I24751), .I1 (g7455), .I2 (g14609));
ND2X1 gate20471(.O (I24752), .I1 (g7455), .I2 (I24751));
ND2X1 gate20472(.O (I24753), .I1 (g14609), .I2 (I24751));
ND2X1 gate20473(.O (g18637), .I1 (I24752), .I2 (I24753));
ND2X1 gate20474(.O (I24763), .I1 (g6194), .I2 (g14573));
ND2X1 gate20475(.O (I24764), .I1 (g6194), .I2 (I24763));
ND2X1 gate20476(.O (I24765), .I1 (g14573), .I2 (I24763));
ND2X1 gate20477(.O (g18644), .I1 (I24764), .I2 (I24765));
ND2X1 gate20478(.O (g18977), .I1 (g15797), .I2 (g3006));
ND2X1 gate20479(.O (I25030), .I1 (g8029), .I2 (g13507));
ND2X1 gate20480(.O (I25031), .I1 (g8029), .I2 (I25030));
ND2X1 gate20481(.O (I25032), .I1 (g13507), .I2 (I25030));
ND2X1 gate20482(.O (g18980), .I1 (I25031), .I2 (I25032));
ND2X1 gate20483(.O (g19067), .I1 (g16554), .I2 (g16578));
ND2X1 gate20484(.O (g19084), .I1 (g16586), .I2 (g16602));
ND2X1 gate20485(.O (g19103), .I1 (g18590), .I2 (g2924));
ND2X1 gate20486(.O (g19121), .I1 (g16682), .I2 (g16697));
ND2X1 gate20487(.O (g19128), .I1 (g16708), .I2 (g16728));
ND2X1 gate20488(.O (g19135), .I1 (g16739), .I2 (g16770));
ND2X1 gate20489(.O (g19138), .I1 (g16781), .I2 (g16797));
ND2X1 gate20490(.O (g19141), .I1 (g3088), .I2 (g16825));
ND2X1 gate20491(.O (g19152), .I1 (g5378), .I2 (g18884));
ND2X1 gate20492(.O (I25532), .I1 (g52), .I2 (g18179));
ND2X1 gate20493(.O (I25533), .I1 (g52), .I2 (I25532));
ND2X1 gate20494(.O (I25534), .I1 (g18179), .I2 (I25532));
ND2X1 gate20495(.O (g19261), .I1 (I25533), .I2 (I25534));
ND2X1 gate20496(.O (I25539), .I1 (g92), .I2 (g18174));
ND2X1 gate20497(.O (I25540), .I1 (g92), .I2 (I25539));
ND2X1 gate20498(.O (I25541), .I1 (g18174), .I2 (I25539));
ND2X1 gate20499(.O (g19262), .I1 (I25540), .I2 (I25541));
ND2X1 gate20500(.O (I25560), .I1 (g56), .I2 (g17724));
ND2X1 gate20501(.O (I25561), .I1 (g56), .I2 (I25560));
ND2X1 gate20502(.O (I25562), .I1 (g17724), .I2 (I25560));
ND2X1 gate20503(.O (g19271), .I1 (I25561), .I2 (I25562));
ND2X1 gate20504(.O (I25571), .I1 (g740), .I2 (g18286));
ND2X1 gate20505(.O (I25572), .I1 (g740), .I2 (I25571));
ND2X1 gate20506(.O (I25573), .I1 (g18286), .I2 (I25571));
ND2X1 gate20507(.O (g19276), .I1 (I25572), .I2 (I25573));
ND2X1 gate20508(.O (I25578), .I1 (g780), .I2 (g18281));
ND2X1 gate20509(.O (I25579), .I1 (g780), .I2 (I25578));
ND2X1 gate20510(.O (I25580), .I1 (g18281), .I2 (I25578));
ND2X1 gate20511(.O (g19277), .I1 (I25579), .I2 (I25580));
ND2X1 gate20512(.O (I25595), .I1 (g61), .I2 (g18074));
ND2X1 gate20513(.O (I25596), .I1 (g61), .I2 (I25595));
ND2X1 gate20514(.O (I25597), .I1 (g18074), .I2 (I25595));
ND2X1 gate20515(.O (g19286), .I1 (I25596), .I2 (I25597));
ND3X1 gate20516(.O (g19288), .I1 (g14685), .I2 (g8580), .I3 (g17057));
ND2X1 gate20517(.O (I25605), .I1 (g744), .I2 (g17825));
ND2X1 gate20518(.O (I25606), .I1 (g744), .I2 (I25605));
ND2X1 gate20519(.O (I25607), .I1 (g17825), .I2 (I25605));
ND2X1 gate20520(.O (g19290), .I1 (I25606), .I2 (I25607));
ND2X1 gate20521(.O (I25616), .I1 (g1426), .I2 (g18379));
ND2X1 gate20522(.O (I25617), .I1 (g1426), .I2 (I25616));
ND2X1 gate20523(.O (I25618), .I1 (g18379), .I2 (I25616));
ND2X1 gate20524(.O (g19295), .I1 (I25617), .I2 (I25618));
ND2X1 gate20525(.O (I25623), .I1 (g1466), .I2 (g18374));
ND2X1 gate20526(.O (I25624), .I1 (g1466), .I2 (I25623));
ND2X1 gate20527(.O (I25625), .I1 (g18374), .I2 (I25623));
ND2X1 gate20528(.O (g19296), .I1 (I25624), .I2 (I25625));
ND2X1 gate20529(.O (I25633), .I1 (g65), .I2 (g17640));
ND2X1 gate20530(.O (I25634), .I1 (g65), .I2 (I25633));
ND2X1 gate20531(.O (I25635), .I1 (g17640), .I2 (I25633));
ND2X1 gate20532(.O (g19300), .I1 (I25634), .I2 (I25635));
ND2X1 gate20533(.O (I25643), .I1 (g749), .I2 (g18190));
ND2X1 gate20534(.O (I25644), .I1 (g749), .I2 (I25643));
ND2X1 gate20535(.O (I25645), .I1 (g18190), .I2 (I25643));
ND2X1 gate20536(.O (g19304), .I1 (I25644), .I2 (I25645));
ND3X1 gate20537(.O (g19306), .I1 (g14719), .I2 (g8587), .I3 (g17092));
ND2X1 gate20538(.O (I25653), .I1 (g1430), .I2 (g17937));
ND2X1 gate20539(.O (I25654), .I1 (g1430), .I2 (I25653));
ND2X1 gate20540(.O (I25655), .I1 (g17937), .I2 (I25653));
ND2X1 gate20541(.O (g19308), .I1 (I25654), .I2 (I25655));
ND2X1 gate20542(.O (I25664), .I1 (g2120), .I2 (g18474));
ND2X1 gate20543(.O (I25665), .I1 (g2120), .I2 (I25664));
ND2X1 gate20544(.O (I25666), .I1 (g18474), .I2 (I25664));
ND2X1 gate20545(.O (g19313), .I1 (I25665), .I2 (I25666));
ND2X1 gate20546(.O (I25671), .I1 (g2160), .I2 (g18469));
ND2X1 gate20547(.O (I25672), .I1 (g2160), .I2 (I25671));
ND2X1 gate20548(.O (I25673), .I1 (g18469), .I2 (I25671));
ND2X1 gate20549(.O (g19314), .I1 (I25672), .I2 (I25673));
ND2X1 gate20550(.O (I25681), .I1 (g70), .I2 (g17974));
ND2X1 gate20551(.O (I25682), .I1 (g70), .I2 (I25681));
ND2X1 gate20552(.O (I25683), .I1 (g17974), .I2 (I25681));
ND2X1 gate20553(.O (g19318), .I1 (I25682), .I2 (I25683));
ND2X1 gate20554(.O (I25690), .I1 (g753), .I2 (g17741));
ND2X1 gate20555(.O (I25691), .I1 (g753), .I2 (I25690));
ND2X1 gate20556(.O (I25692), .I1 (g17741), .I2 (I25690));
ND2X1 gate20557(.O (g19321), .I1 (I25691), .I2 (I25692));
ND2X1 gate20558(.O (I25700), .I1 (g1435), .I2 (g18297));
ND2X1 gate20559(.O (I25701), .I1 (g1435), .I2 (I25700));
ND2X1 gate20560(.O (I25702), .I1 (g18297), .I2 (I25700));
ND2X1 gate20561(.O (g19325), .I1 (I25701), .I2 (I25702));
ND3X1 gate20562(.O (g19327), .I1 (g14747), .I2 (g8594), .I3 (g17130));
ND2X1 gate20563(.O (I25710), .I1 (g2124), .I2 (g18048));
ND2X1 gate20564(.O (I25711), .I1 (g2124), .I2 (I25710));
ND2X1 gate20565(.O (I25712), .I1 (g18048), .I2 (I25710));
ND2X1 gate20566(.O (g19329), .I1 (I25711), .I2 (I25712));
ND2X1 gate20567(.O (I25721), .I1 (g74), .I2 (g18341));
ND2X1 gate20568(.O (I25722), .I1 (g74), .I2 (I25721));
ND2X1 gate20569(.O (I25723), .I1 (g18341), .I2 (I25721));
ND2X1 gate20570(.O (g19334), .I1 (I25722), .I2 (I25723));
ND2X1 gate20571(.O (I25731), .I1 (g758), .I2 (g18091));
ND2X1 gate20572(.O (I25732), .I1 (g758), .I2 (I25731));
ND2X1 gate20573(.O (I25733), .I1 (g18091), .I2 (I25731));
ND2X1 gate20574(.O (g19345), .I1 (I25732), .I2 (I25733));
ND2X1 gate20575(.O (I25740), .I1 (g1439), .I2 (g17842));
ND2X1 gate20576(.O (I25741), .I1 (g1439), .I2 (I25740));
ND2X1 gate20577(.O (I25742), .I1 (g17842), .I2 (I25740));
ND2X1 gate20578(.O (g19348), .I1 (I25741), .I2 (I25742));
ND2X1 gate20579(.O (I25750), .I1 (g2129), .I2 (g18390));
ND2X1 gate20580(.O (I25751), .I1 (g2129), .I2 (I25750));
ND2X1 gate20581(.O (I25752), .I1 (g18390), .I2 (I25750));
ND2X1 gate20582(.O (g19352), .I1 (I25751), .I2 (I25752));
ND3X1 gate20583(.O (g19354), .I1 (g14768), .I2 (g8605), .I3 (g17157));
ND2X1 gate20584(.O (I25761), .I1 (g79), .I2 (g17882));
ND2X1 gate20585(.O (I25762), .I1 (g79), .I2 (I25761));
ND2X1 gate20586(.O (I25763), .I1 (g17882), .I2 (I25761));
ND2X1 gate20587(.O (g19357), .I1 (I25762), .I2 (I25763));
ND2X1 gate20588(.O (I25771), .I1 (g762), .I2 (g18436));
ND2X1 gate20589(.O (I25772), .I1 (g762), .I2 (I25771));
ND2X1 gate20590(.O (I25773), .I1 (g18436), .I2 (I25771));
ND2X1 gate20591(.O (g19368), .I1 (I25772), .I2 (I25773));
ND2X1 gate20592(.O (I25781), .I1 (g1444), .I2 (g18207));
ND2X1 gate20593(.O (I25782), .I1 (g1444), .I2 (I25781));
ND2X1 gate20594(.O (I25783), .I1 (g18207), .I2 (I25781));
ND2X1 gate20595(.O (g19379), .I1 (I25782), .I2 (I25783));
ND2X1 gate20596(.O (I25790), .I1 (g2133), .I2 (g17954));
ND2X1 gate20597(.O (I25791), .I1 (g2133), .I2 (I25790));
ND2X1 gate20598(.O (I25792), .I1 (g17954), .I2 (I25790));
ND2X1 gate20599(.O (g19382), .I1 (I25791), .I2 (I25792));
ND2X1 gate20600(.O (I25800), .I1 (g83), .I2 (g18265));
ND2X1 gate20601(.O (I25801), .I1 (g83), .I2 (I25800));
ND2X1 gate20602(.O (I25802), .I1 (g18265), .I2 (I25800));
ND2X1 gate20603(.O (g19386), .I1 (I25801), .I2 (I25802));
ND2X1 gate20604(.O (I25809), .I1 (g767), .I2 (g17993));
ND2X1 gate20605(.O (I25810), .I1 (g767), .I2 (I25809));
ND2X1 gate20606(.O (I25811), .I1 (g17993), .I2 (I25809));
ND2X1 gate20607(.O (g19389), .I1 (I25810), .I2 (I25811));
ND2X1 gate20608(.O (I25819), .I1 (g1448), .I2 (g18509));
ND2X1 gate20609(.O (I25820), .I1 (g1448), .I2 (I25819));
ND2X1 gate20610(.O (I25821), .I1 (g18509), .I2 (I25819));
ND2X1 gate20611(.O (g19400), .I1 (I25820), .I2 (I25821));
ND2X1 gate20612(.O (I25829), .I1 (g2138), .I2 (g18314));
ND2X1 gate20613(.O (I25830), .I1 (g2138), .I2 (I25829));
ND2X1 gate20614(.O (I25831), .I1 (g18314), .I2 (I25829));
ND2X1 gate20615(.O (g19411), .I1 (I25830), .I2 (I25831));
ND2X1 gate20616(.O (I25838), .I1 (g88), .I2 (g17802));
ND2X1 gate20617(.O (I25839), .I1 (g88), .I2 (I25838));
ND2X1 gate20618(.O (I25840), .I1 (g17802), .I2 (I25838));
ND2X1 gate20619(.O (g19414), .I1 (I25839), .I2 (I25840));
ND2X1 gate20620(.O (I25846), .I1 (g771), .I2 (g18358));
ND2X1 gate20621(.O (I25847), .I1 (g771), .I2 (I25846));
ND2X1 gate20622(.O (I25848), .I1 (g18358), .I2 (I25846));
ND2X1 gate20623(.O (g19416), .I1 (I25847), .I2 (I25848));
ND2X1 gate20624(.O (I25855), .I1 (g1453), .I2 (g18110));
ND2X1 gate20625(.O (I25856), .I1 (g1453), .I2 (I25855));
ND2X1 gate20626(.O (I25857), .I1 (g18110), .I2 (I25855));
ND2X1 gate20627(.O (g19419), .I1 (I25856), .I2 (I25857));
ND2X1 gate20628(.O (I25865), .I1 (g2142), .I2 (g18573));
ND2X1 gate20629(.O (I25866), .I1 (g2142), .I2 (I25865));
ND2X1 gate20630(.O (I25867), .I1 (g18573), .I2 (I25865));
ND2X1 gate20631(.O (g19430), .I1 (I25866), .I2 (I25867));
ND2X1 gate20632(.O (I25880), .I1 (g776), .I2 (g17914));
ND2X1 gate20633(.O (I25881), .I1 (g776), .I2 (I25880));
ND2X1 gate20634(.O (I25882), .I1 (g17914), .I2 (I25880));
ND2X1 gate20635(.O (g19451), .I1 (I25881), .I2 (I25882));
ND2X1 gate20636(.O (I25888), .I1 (g1457), .I2 (g18453));
ND2X1 gate20637(.O (I25889), .I1 (g1457), .I2 (I25888));
ND2X1 gate20638(.O (I25890), .I1 (g18453), .I2 (I25888));
ND2X1 gate20639(.O (g19453), .I1 (I25889), .I2 (I25890));
ND2X1 gate20640(.O (I25897), .I1 (g2147), .I2 (g18226));
ND2X1 gate20641(.O (I25898), .I1 (g2147), .I2 (I25897));
ND2X1 gate20642(.O (I25899), .I1 (g18226), .I2 (I25897));
ND2X1 gate20643(.O (g19456), .I1 (I25898), .I2 (I25899));
ND2X1 gate20644(.O (I25913), .I1 (g1462), .I2 (g18025));
ND2X1 gate20645(.O (I25914), .I1 (g1462), .I2 (I25913));
ND2X1 gate20646(.O (I25915), .I1 (g18025), .I2 (I25913));
ND2X1 gate20647(.O (g19478), .I1 (I25914), .I2 (I25915));
ND2X1 gate20648(.O (I25921), .I1 (g2151), .I2 (g18526));
ND2X1 gate20649(.O (I25922), .I1 (g2151), .I2 (I25921));
ND2X1 gate20650(.O (I25923), .I1 (g18526), .I2 (I25921));
ND2X1 gate20651(.O (g19480), .I1 (I25922), .I2 (I25923));
ND2X1 gate20652(.O (I25938), .I1 (g2156), .I2 (g18142));
ND2X1 gate20653(.O (I25939), .I1 (g2156), .I2 (I25938));
ND2X1 gate20654(.O (I25940), .I1 (g18142), .I2 (I25938));
ND2X1 gate20655(.O (g19501), .I1 (I25939), .I2 (I25940));
ND2X1 gate20656(.O (g19865), .I1 (g16607), .I2 (g9636));
ND2X1 gate20657(.O (g19896), .I1 (g16625), .I2 (g9782));
ND2X1 gate20658(.O (g19921), .I1 (g16639), .I2 (g9928));
ND2X1 gate20659(.O (g19936), .I1 (g16650), .I2 (g10082));
ND2X1 gate20660(.O (g19954), .I1 (g17186), .I2 (g92));
ND2X1 gate20661(.O (g19984), .I1 (g17197), .I2 (g780));
ND2X1 gate20662(.O (g20022), .I1 (g17204), .I2 (g1466));
ND2X1 gate20663(.O (g20064), .I1 (g17209), .I2 (g2160));
ND2X1 gate20664(.O (g20473), .I1 (g18085), .I2 (g646));
ND2X1 gate20665(.O (g20481), .I1 (g18201), .I2 (g1332));
ND2X1 gate20666(.O (g20487), .I1 (g18308), .I2 (g2026));
ND2X1 gate20667(.O (g20493), .I1 (g18401), .I2 (g2720));
ND2X1 gate20668(.O (g20497), .I1 (g5410), .I2 (g18886));
ND2X1 gate20669(.O (g20522), .I1 (g16501), .I2 (g16515));
ND2X1 gate20670(.O (g20537), .I1 (g18626), .I2 (g3036));
ND2X1 gate20671(.O (g20542), .I1 (g16523), .I2 (g16546));
ND2X1 gate20672(.O (g20633), .I1 (g20164), .I2 (g3254));
ND2X1 gate20673(.O (g20648), .I1 (g20164), .I2 (g3254));
ND2X1 gate20674(.O (g20658), .I1 (g20198), .I2 (g3410));
ND2X1 gate20675(.O (g20672), .I1 (g20164), .I2 (g3254));
ND2X1 gate20676(.O (g20683), .I1 (g20198), .I2 (g3410));
ND2X1 gate20677(.O (g20693), .I1 (g20228), .I2 (g3566));
ND2X1 gate20678(.O (g20700), .I1 (g20153), .I2 (g2903));
ND2X1 gate20679(.O (g20703), .I1 (g20164), .I2 (g3254));
ND2X1 gate20680(.O (g20707), .I1 (g20198), .I2 (g3410));
ND2X1 gate20681(.O (g20718), .I1 (g20228), .I2 (g3566));
ND2X1 gate20682(.O (g20728), .I1 (g20255), .I2 (g3722));
ND2X1 gate20683(.O (g20738), .I1 (g20198), .I2 (g3410));
ND2X1 gate20684(.O (g20742), .I1 (g20228), .I2 (g3566));
ND2X1 gate20685(.O (g20753), .I1 (g20255), .I2 (g3722));
ND2X1 gate20686(.O (g20775), .I1 (g20228), .I2 (g3566));
ND2X1 gate20687(.O (g20779), .I1 (g20255), .I2 (g3722));
ND2X1 gate20688(.O (g20805), .I1 (g20255), .I2 (g3722));
ND2X1 gate20689(.O (g20825), .I1 (g19219), .I2 (g15959));
ND2X1 gate20690(.O (g21659), .I1 (g20164), .I2 (g6314));
ND2X1 gate20691(.O (I28189), .I1 (g14079), .I2 (g19444));
ND2X1 gate20692(.O (I28190), .I1 (g14079), .I2 (I28189));
ND2X1 gate20693(.O (I28191), .I1 (g19444), .I2 (I28189));
ND2X1 gate20694(.O (g21660), .I1 (I28190), .I2 (I28191));
ND2X1 gate20695(.O (g21685), .I1 (g20164), .I2 (g6232));
ND2X1 gate20696(.O (g21686), .I1 (g20164), .I2 (g6314));
ND2X1 gate20697(.O (g21688), .I1 (g20198), .I2 (g6519));
ND2X1 gate20698(.O (I28217), .I1 (g14194), .I2 (g19471));
ND2X1 gate20699(.O (I28218), .I1 (g14194), .I2 (I28217));
ND2X1 gate20700(.O (I28219), .I1 (g19471), .I2 (I28217));
ND2X1 gate20701(.O (g21689), .I1 (I28218), .I2 (I28219));
ND2X1 gate20702(.O (g21714), .I1 (g20164), .I2 (g6232));
ND2X1 gate20703(.O (g21715), .I1 (g20164), .I2 (g6314));
ND4X1 gate20704(.O (g21720), .I1 (g14256), .I2 (g15177), .I3 (g19871), .I4 (g19842));
ND2X1 gate20705(.O (g21721), .I1 (g20198), .I2 (g6369));
ND2X1 gate20706(.O (g21722), .I1 (g20198), .I2 (g6519));
ND2X1 gate20707(.O (g21724), .I1 (g20228), .I2 (g6783));
ND2X1 gate20708(.O (I28247), .I1 (g14309), .I2 (g19494));
ND2X1 gate20709(.O (I28248), .I1 (g14309), .I2 (I28247));
ND2X1 gate20710(.O (I28249), .I1 (g19494), .I2 (I28247));
ND2X1 gate20711(.O (g21725), .I1 (I28248), .I2 (I28249));
ND2X1 gate20712(.O (g21736), .I1 (g20164), .I2 (g6232));
ND2X1 gate20713(.O (g21737), .I1 (g20164), .I2 (g6314));
ND2X1 gate20714(.O (g21740), .I1 (g20198), .I2 (g6369));
ND2X1 gate20715(.O (g21741), .I1 (g20198), .I2 (g6519));
ND4X1 gate20716(.O (g21746), .I1 (g14378), .I2 (g15263), .I3 (g19902), .I4 (g19875));
ND2X1 gate20717(.O (g21747), .I1 (g20228), .I2 (g6574));
ND2X1 gate20718(.O (g21748), .I1 (g20228), .I2 (g6783));
ND2X1 gate20719(.O (g21750), .I1 (g20255), .I2 (g7085));
ND2X1 gate20720(.O (I28271), .I1 (g14431), .I2 (g19515));
ND2X1 gate20721(.O (I28272), .I1 (g14431), .I2 (I28271));
ND2X1 gate20722(.O (I28273), .I1 (g19515), .I2 (I28271));
ND2X1 gate20723(.O (g21751), .I1 (I28272), .I2 (I28273));
ND2X1 gate20724(.O (g21759), .I1 (g20164), .I2 (g6232));
ND2X1 gate20725(.O (g21760), .I1 (g20198), .I2 (g6369));
ND2X1 gate20726(.O (g21761), .I1 (g20198), .I2 (g6519));
ND2X1 gate20727(.O (g21764), .I1 (g20228), .I2 (g6574));
ND2X1 gate20728(.O (g21765), .I1 (g20228), .I2 (g6783));
ND4X1 gate20729(.O (g21770), .I1 (g14490), .I2 (g15355), .I3 (g19927), .I4 (g19906));
ND2X1 gate20730(.O (g21771), .I1 (g20255), .I2 (g6838));
ND2X1 gate20731(.O (g21772), .I1 (g20255), .I2 (g7085));
ND2X1 gate20732(.O (g21775), .I1 (g20198), .I2 (g6369));
ND2X1 gate20733(.O (g21776), .I1 (g20228), .I2 (g6574));
ND2X1 gate20734(.O (g21777), .I1 (g20228), .I2 (g6783));
ND2X1 gate20735(.O (g21780), .I1 (g20255), .I2 (g6838));
ND2X1 gate20736(.O (g21781), .I1 (g20255), .I2 (g7085));
ND4X1 gate20737(.O (g21786), .I1 (g14577), .I2 (g15441), .I3 (g19942), .I4 (g19931));
ND2X1 gate20738(.O (g21790), .I1 (g20228), .I2 (g6574));
ND2X1 gate20739(.O (g21791), .I1 (g20255), .I2 (g6838));
ND2X1 gate20740(.O (g21792), .I1 (g20255), .I2 (g7085));
ND2X1 gate20741(.O (g21804), .I1 (g20255), .I2 (g6838));
ND3X1 gate20742(.O (g21848), .I1 (g17807), .I2 (g19181), .I3 (g19186));
ND3X1 gate20743(.O (g21850), .I1 (g17979), .I2 (g19187), .I3 (g19191));
ND3X1 gate20744(.O (g21855), .I1 (g17919), .I2 (g19188), .I3 (g19193));
ND3X1 gate20745(.O (g21857), .I1 (g18079), .I2 (g19192), .I3 (g19200));
ND3X1 gate20746(.O (g21858), .I1 (g18096), .I2 (g19194), .I3 (g19202));
ND3X1 gate20747(.O (g21859), .I1 (g18030), .I2 (g19195), .I3 (g19204));
ND3X1 gate20748(.O (g21860), .I1 (g18270), .I2 (g19201), .I3 (g19209));
ND3X1 gate20749(.O (g21862), .I1 (g18195), .I2 (g19203), .I3 (g19211));
ND3X1 gate20750(.O (g21863), .I1 (g18212), .I2 (g19205), .I3 (g19213));
ND3X1 gate20751(.O (g21864), .I1 (g18147), .I2 (g19206), .I3 (g19215));
ND3X1 gate20752(.O (g21865), .I1 (g18424), .I2 (g19210), .I3 (g19221));
ND3X1 gate20753(.O (g21866), .I1 (g18363), .I2 (g19212), .I3 (g19222));
ND3X1 gate20754(.O (g21868), .I1 (g18302), .I2 (g19214), .I3 (g19224));
ND3X1 gate20755(.O (g21869), .I1 (g18319), .I2 (g19216), .I3 (g19226));
ND3X1 gate20756(.O (g21870), .I1 (g18497), .I2 (g19223), .I3 (g19231));
ND3X1 gate20757(.O (g21871), .I1 (g18458), .I2 (g19225), .I3 (g19232));
ND3X1 gate20758(.O (g21873), .I1 (g18395), .I2 (g19227), .I3 (g19234));
ND3X1 gate20759(.O (g21874), .I1 (g18561), .I2 (g19233), .I3 (g19244));
ND3X1 gate20760(.O (g21875), .I1 (g18531), .I2 (g19235), .I3 (g19245));
ND3X1 gate20761(.O (g21877), .I1 (g18611), .I2 (g19246), .I3 (g19257));
ND3X1 gate20762(.O (g21879), .I1 (g18419), .I2 (g19250), .I3 (g19263));
ND3X1 gate20763(.O (g21881), .I1 (g18492), .I2 (g19264), .I3 (g19278));
ND3X1 gate20764(.O (g21885), .I1 (g18556), .I2 (g19279), .I3 (g19297));
ND3X1 gate20765(.O (g21888), .I1 (g18606), .I2 (g19298), .I3 (g19315));
ND2X1 gate20766(.O (g21903), .I1 (g20008), .I2 (g3013));
ND3X1 gate20767(.O (g21976), .I1 (g19242), .I2 (g21120), .I3 (g19275));
ND3X1 gate20768(.O (g21983), .I1 (g19255), .I2 (g21139), .I3 (g19294));
ND2X1 gate20769(.O (g21989), .I1 (g21048), .I2 (g18623));
ND2X1 gate20770(.O (g21991), .I1 (g21501), .I2 (g21536));
ND3X1 gate20771(.O (g21996), .I1 (g19268), .I2 (g21159), .I3 (g19312));
ND2X1 gate20772(.O (g22002), .I1 (g21065), .I2 (g21711));
ND2X1 gate20773(.O (g22005), .I1 (g21540), .I2 (g21572));
ND3X1 gate20774(.O (g22009), .I1 (g19283), .I2 (g21179), .I3 (g19333));
ND2X1 gate20775(.O (g22016), .I1 (g21576), .I2 (g21605));
ND2X1 gate20776(.O (g22021), .I1 (g21609), .I2 (g21634));
ND3X1 gate20777(.O (g22050), .I1 (g19450), .I2 (g21244), .I3 (g19503));
ND3X1 gate20778(.O (g22069), .I1 (g19477), .I2 (g21253), .I3 (g19522));
ND2X1 gate20779(.O (g22083), .I1 (g21774), .I2 (g21787));
ND3X1 gate20780(.O (g22093), .I1 (g19500), .I2 (g21261), .I3 (g19532));
ND2X1 gate20781(.O (g22108), .I1 (g21789), .I2 (g21801));
ND3X1 gate20782(.O (g22118), .I1 (g19521), .I2 (g21269), .I3 (g19542));
ND2X1 gate20783(.O (g22134), .I1 (g21803), .I2 (g21809));
ND2X1 gate20784(.O (g22157), .I1 (g21811), .I2 (g21816));
ND2X1 gate20785(.O (I28726), .I1 (g21887), .I2 (g13519));
ND2X1 gate20786(.O (I28727), .I1 (g21887), .I2 (I28726));
ND2X1 gate20787(.O (I28728), .I1 (g13519), .I2 (I28726));
ND2X1 gate20788(.O (g22188), .I1 (I28727), .I2 (I28728));
ND2X1 gate20789(.O (I28741), .I1 (g21890), .I2 (g13530));
ND2X1 gate20790(.O (I28742), .I1 (g21890), .I2 (I28741));
ND2X1 gate20791(.O (I28743), .I1 (g13530), .I2 (I28741));
ND2X1 gate20792(.O (g22197), .I1 (I28742), .I2 (I28743));
ND2X1 gate20793(.O (I28753), .I1 (g21893), .I2 (g13541));
ND2X1 gate20794(.O (I28754), .I1 (g21893), .I2 (I28753));
ND2X1 gate20795(.O (I28755), .I1 (g13541), .I2 (I28753));
ND2X1 gate20796(.O (g22203), .I1 (I28754), .I2 (I28755));
ND2X1 gate20797(.O (I28765), .I1 (g21901), .I2 (g13552));
ND2X1 gate20798(.O (I28766), .I1 (g21901), .I2 (I28765));
ND2X1 gate20799(.O (I28767), .I1 (g13552), .I2 (I28765));
ND2X1 gate20800(.O (g22209), .I1 (I28766), .I2 (I28767));
ND3X1 gate20801(.O (g22317), .I1 (g21152), .I2 (g21241), .I3 (g21136));
ND3X1 gate20802(.O (g22339), .I1 (g14442), .I2 (g21149), .I3 (g10694));
ND3X1 gate20803(.O (g22342), .I1 (g21172), .I2 (g21249), .I3 (g21156));
ND3X1 gate20804(.O (g22362), .I1 (g14529), .I2 (g21169), .I3 (g10714));
ND3X1 gate20805(.O (g22365), .I1 (g21192), .I2 (g21258), .I3 (g21176));
ND3X1 gate20806(.O (g22381), .I1 (g21211), .I2 (g14442), .I3 (g10694));
ND3X1 gate20807(.O (g22382), .I1 (g14584), .I2 (g21189), .I3 (g10735));
ND3X1 gate20808(.O (g22385), .I1 (g21207), .I2 (g21266), .I3 (g21196));
ND3X1 gate20809(.O (g22396), .I1 (g21219), .I2 (g14529), .I3 (g10714));
ND3X1 gate20810(.O (g22397), .I1 (g14618), .I2 (g21204), .I3 (g10754));
ND3X1 gate20811(.O (g22399), .I1 (g21230), .I2 (g14584), .I3 (g10735));
ND3X1 gate20812(.O (g22400), .I1 (g21235), .I2 (g14618), .I3 (g10754));
ND2X1 gate20813(.O (g22608), .I1 (g20842), .I2 (g20885));
ND2X1 gate20814(.O (g22644), .I1 (g20850), .I2 (g20904));
ND2X1 gate20815(.O (g22668), .I1 (g16075), .I2 (g21271));
ND2X1 gate20816(.O (g22680), .I1 (g20858), .I2 (g20928));
ND2X1 gate20817(.O (g22708), .I1 (g16113), .I2 (g21278));
ND2X1 gate20818(.O (g22720), .I1 (g20866), .I2 (g20956));
ND2X1 gate20819(.O (g22739), .I1 (g16164), .I2 (g21285));
ND2X1 gate20820(.O (g22771), .I1 (g16223), .I2 (g21293));
ND3X1 gate20821(.O (g22809), .I1 (g21850), .I2 (g21848), .I3 (g21879));
ND3X1 gate20822(.O (g22844), .I1 (g21865), .I2 (g21860), .I3 (g21857));
ND2X1 gate20823(.O (g22845), .I1 (g19441), .I2 (g20885));
ND2X1 gate20824(.O (g22846), .I1 (g8278), .I2 (g21660));
ND3X1 gate20825(.O (g22850), .I1 (g21858), .I2 (g21855), .I3 (g21881));
ND2X1 gate20826(.O (g22876), .I1 (g21238), .I2 (g83));
ND3X1 gate20827(.O (g22879), .I1 (g21870), .I2 (g21866), .I3 (g21862));
ND2X1 gate20828(.O (g22880), .I1 (g19468), .I2 (g20904));
ND2X1 gate20829(.O (g22881), .I1 (g8287), .I2 (g21689));
ND3X1 gate20830(.O (g22885), .I1 (g21863), .I2 (g21859), .I3 (g21885));
ND2X1 gate20831(.O (g22911), .I1 (g21246), .I2 (g771));
ND3X1 gate20832(.O (g22914), .I1 (g21874), .I2 (g21871), .I3 (g21868));
ND2X1 gate20833(.O (g22915), .I1 (g19491), .I2 (g20928));
ND2X1 gate20834(.O (g22916), .I1 (g8296), .I2 (g21725));
ND3X1 gate20835(.O (g22920), .I1 (g21869), .I2 (g21864), .I3 (g21888));
ND2X1 gate20836(.O (g22936), .I1 (g21255), .I2 (g1457));
ND3X1 gate20837(.O (g22939), .I1 (g21877), .I2 (g21875), .I3 (g21873));
ND2X1 gate20838(.O (g22940), .I1 (g19512), .I2 (g20956));
ND2X1 gate20839(.O (g22941), .I1 (g8305), .I2 (g21751));
ND2X1 gate20840(.O (g22942), .I1 (g21263), .I2 (g2151));
ND2X1 gate20841(.O (g22992), .I1 (g21636), .I2 (g672));
ND2X1 gate20842(.O (g23003), .I1 (g21667), .I2 (g1358));
ND2X1 gate20843(.O (g23017), .I1 (g21696), .I2 (g2052));
ND2X1 gate20844(.O (g23033), .I1 (g21732), .I2 (g2746));
ND2X1 gate20845(.O (g23320), .I1 (g23066), .I2 (g23051));
ND2X1 gate20846(.O (g23325), .I1 (g23080), .I2 (g23070));
ND2X1 gate20847(.O (g23331), .I1 (g22999), .I2 (g22174));
ND2X1 gate20848(.O (g23335), .I1 (g23096), .I2 (g23083));
ND2X1 gate20849(.O (g23340), .I1 (g23013), .I2 (g22189));
ND2X1 gate20850(.O (g23344), .I1 (g23113), .I2 (g23099));
ND2X1 gate20851(.O (g23349), .I1 (g23029), .I2 (g22198));
ND2X1 gate20852(.O (g23353), .I1 (g23046), .I2 (g22204));
ND2X1 gate20853(.O (g23360), .I1 (g21980), .I2 (g21975));
ND2X1 gate20854(.O (g23364), .I1 (g21987), .I2 (g21981));
ND2X1 gate20855(.O (g23368), .I1 (g23135), .I2 (g22288));
ND2X1 gate20856(.O (g23372), .I1 (g22000), .I2 (g21988));
ND2X1 gate20857(.O (g23376), .I1 (g18435), .I2 (g22812));
ND2X1 gate20858(.O (g23377), .I1 (g21968), .I2 (g22308));
ND2X1 gate20859(.O (g23381), .I1 (g22013), .I2 (g22001));
ND2X1 gate20860(.O (g23387), .I1 (g18508), .I2 (g22852));
ND2X1 gate20861(.O (g23388), .I1 (g21971), .I2 (g22336));
ND2X1 gate20862(.O (g23394), .I1 (g18572), .I2 (g22887));
ND2X1 gate20863(.O (g23395), .I1 (g21973), .I2 (g22361));
ND2X1 gate20864(.O (g23402), .I1 (g18622), .I2 (g22922));
ND3X1 gate20865(.O (g23478), .I1 (g22809), .I2 (g14442), .I3 (g10694));
ND3X1 gate20866(.O (g23486), .I1 (g22844), .I2 (g14442), .I3 (g10694));
ND3X1 gate20867(.O (g23489), .I1 (g22850), .I2 (g14529), .I3 (g10714));
ND3X1 gate20868(.O (g23495), .I1 (g10694), .I2 (g14442), .I3 (g22316));
ND3X1 gate20869(.O (g23502), .I1 (g22879), .I2 (g14529), .I3 (g10714));
ND3X1 gate20870(.O (g23505), .I1 (g22885), .I2 (g14584), .I3 (g10735));
ND3X1 gate20871(.O (g23511), .I1 (g10714), .I2 (g14529), .I3 (g22341));
ND3X1 gate20872(.O (g23518), .I1 (g22914), .I2 (g14584), .I3 (g10735));
ND3X1 gate20873(.O (g23521), .I1 (g22920), .I2 (g14618), .I3 (g10754));
ND3X1 gate20874(.O (g23526), .I1 (g10735), .I2 (g14584), .I3 (g22364));
ND3X1 gate20875(.O (g23533), .I1 (g22939), .I2 (g14618), .I3 (g10754));
ND3X1 gate20876(.O (g23537), .I1 (g10754), .I2 (g14618), .I3 (g22384));
ND2X1 gate20877(.O (I30790), .I1 (g22846), .I2 (g14079));
ND2X1 gate20878(.O (I30791), .I1 (g22846), .I2 (I30790));
ND2X1 gate20879(.O (I30792), .I1 (g14079), .I2 (I30790));
ND2X1 gate20880(.O (g23660), .I1 (I30791), .I2 (I30792));
ND2X1 gate20881(.O (I30868), .I1 (g22881), .I2 (g14194));
ND2X1 gate20882(.O (I30869), .I1 (g22881), .I2 (I30868));
ND2X1 gate20883(.O (I30870), .I1 (g14194), .I2 (I30868));
ND2X1 gate20884(.O (g23710), .I1 (I30869), .I2 (I30870));
ND2X1 gate20885(.O (I30952), .I1 (g22916), .I2 (g14309));
ND2X1 gate20886(.O (I30953), .I1 (g22916), .I2 (I30952));
ND2X1 gate20887(.O (I30954), .I1 (g14309), .I2 (I30952));
ND2X1 gate20888(.O (g23764), .I1 (I30953), .I2 (I30954));
ND2X1 gate20889(.O (I31035), .I1 (g22941), .I2 (g14431));
ND2X1 gate20890(.O (I31036), .I1 (g22941), .I2 (I31035));
ND2X1 gate20891(.O (I31037), .I1 (g14431), .I2 (I31035));
ND2X1 gate20892(.O (g23819), .I1 (I31036), .I2 (I31037));
ND2X1 gate20893(.O (g23906), .I1 (g22812), .I2 (g13958));
ND2X1 gate20894(.O (g23936), .I1 (g22812), .I2 (g13922));
ND2X1 gate20895(.O (g23937), .I1 (g22812), .I2 (g13918));
ND2X1 gate20896(.O (g23938), .I1 (g22852), .I2 (g14028));
ND2X1 gate20897(.O (g23953), .I1 (g22812), .I2 (g14525));
ND2X1 gate20898(.O (g23968), .I1 (g22852), .I2 (g13978));
ND2X1 gate20899(.O (g23969), .I1 (g22852), .I2 (g13974));
ND2X1 gate20900(.O (g23970), .I1 (g22887), .I2 (g14119));
ND2X1 gate20901(.O (g23973), .I1 (g22812), .I2 (g14450));
ND2X1 gate20902(.O (g23982), .I1 (g22852), .I2 (g14580));
ND2X1 gate20903(.O (g23997), .I1 (g22887), .I2 (g14048));
ND2X1 gate20904(.O (g23998), .I1 (g22887), .I2 (g14044));
ND2X1 gate20905(.O (g23999), .I1 (g22922), .I2 (g14234));
ND2X1 gate20906(.O (g24002), .I1 (g22812), .I2 (g14355));
ND2X1 gate20907(.O (g24003), .I1 (g22852), .I2 (g14537));
ND2X1 gate20908(.O (g24012), .I1 (g22887), .I2 (g14614));
ND2X1 gate20909(.O (g24027), .I1 (g22922), .I2 (g14139));
ND2X1 gate20910(.O (g24028), .I1 (g22922), .I2 (g14135));
ND2X1 gate20911(.O (g24034), .I1 (g22812), .I2 (g14252));
ND2X1 gate20912(.O (g24036), .I1 (g22852), .I2 (g14467));
ND2X1 gate20913(.O (g24037), .I1 (g22887), .I2 (g14592));
ND2X1 gate20914(.O (g24046), .I1 (g22922), .I2 (g14637));
ND2X1 gate20915(.O (g24052), .I1 (g22812), .I2 (g14171));
ND2X1 gate20916(.O (g24054), .I1 (g22852), .I2 (g14374));
ND2X1 gate20917(.O (g24056), .I1 (g22887), .I2 (g14554));
ND2X1 gate20918(.O (g24057), .I1 (g22922), .I2 (g14626));
ND2X1 gate20919(.O (g24058), .I1 (g22812), .I2 (g14086));
ND2X1 gate20920(.O (g24065), .I1 (g22852), .I2 (g14286));
ND2X1 gate20921(.O (g24067), .I1 (g22887), .I2 (g14486));
ND2X1 gate20922(.O (g24069), .I1 (g22922), .I2 (g14609));
ND2X1 gate20923(.O (g24070), .I1 (g22812), .I2 (g14011));
ND2X1 gate20924(.O (g24071), .I1 (g22852), .I2 (g14201));
ND2X1 gate20925(.O (g24078), .I1 (g22887), .I2 (g14408));
ND2X1 gate20926(.O (g24080), .I1 (g22922), .I2 (g14573));
ND2X1 gate20927(.O (g24081), .I1 (g22852), .I2 (g14102));
ND2X1 gate20928(.O (g24082), .I1 (g22887), .I2 (g14316));
ND2X1 gate20929(.O (g24089), .I1 (g22922), .I2 (g14520));
ND2X1 gate20930(.O (g24090), .I1 (g22887), .I2 (g14217));
ND2X1 gate20931(.O (g24091), .I1 (g22922), .I2 (g14438));
ND2X1 gate20932(.O (g24093), .I1 (g22922), .I2 (g14332));
ND2X1 gate20933(.O (g24100), .I1 (g20885), .I2 (g22175));
ND2X1 gate20934(.O (g24109), .I1 (g20904), .I2 (g22190));
ND2X1 gate20935(.O (g24126), .I1 (g20928), .I2 (g22199));
ND2X1 gate20936(.O (g24145), .I1 (g20956), .I2 (g22205));
ND2X1 gate20937(.O (g24442), .I1 (g23644), .I2 (g3306));
ND2X1 gate20938(.O (g24443), .I1 (g23644), .I2 (g3306));
ND2X1 gate20939(.O (g24444), .I1 (g23694), .I2 (g3462));
ND2X1 gate20940(.O (g24447), .I1 (g23644), .I2 (g3306));
ND2X1 gate20941(.O (g24448), .I1 (g23923), .I2 (g3338));
ND2X1 gate20942(.O (g24449), .I1 (g23694), .I2 (g3462));
ND2X1 gate20943(.O (g24450), .I1 (g23748), .I2 (g3618));
ND2X1 gate20944(.O (g24451), .I1 (g23644), .I2 (g3306));
ND2X1 gate20945(.O (g24452), .I1 (g23923), .I2 (g3338));
ND2X1 gate20946(.O (g24453), .I1 (g23694), .I2 (g3462));
ND2X1 gate20947(.O (g24454), .I1 (g23955), .I2 (g3494));
ND2X1 gate20948(.O (g24455), .I1 (g23748), .I2 (g3618));
ND2X1 gate20949(.O (g24456), .I1 (g23803), .I2 (g3774));
ND2X1 gate20950(.O (g24457), .I1 (g23923), .I2 (g3338));
ND2X1 gate20951(.O (g24458), .I1 (g23694), .I2 (g3462));
ND2X1 gate20952(.O (g24459), .I1 (g23955), .I2 (g3494));
ND2X1 gate20953(.O (g24460), .I1 (g23748), .I2 (g3618));
ND2X1 gate20954(.O (g24461), .I1 (g23984), .I2 (g3650));
ND2X1 gate20955(.O (g24462), .I1 (g23803), .I2 (g3774));
ND2X1 gate20956(.O (g24463), .I1 (g23923), .I2 (g3338));
ND2X1 gate20957(.O (g24464), .I1 (g23955), .I2 (g3494));
ND2X1 gate20958(.O (g24465), .I1 (g23748), .I2 (g3618));
ND2X1 gate20959(.O (g24466), .I1 (g23984), .I2 (g3650));
ND2X1 gate20960(.O (g24467), .I1 (g23803), .I2 (g3774));
ND2X1 gate20961(.O (g24468), .I1 (g24014), .I2 (g3806));
ND2X1 gate20962(.O (g24469), .I1 (g23955), .I2 (g3494));
ND2X1 gate20963(.O (g24470), .I1 (g23984), .I2 (g3650));
ND2X1 gate20964(.O (g24471), .I1 (g23803), .I2 (g3774));
ND2X1 gate20965(.O (g24472), .I1 (g24014), .I2 (g3806));
ND2X1 gate20966(.O (g24474), .I1 (g23984), .I2 (g3650));
ND2X1 gate20967(.O (g24475), .I1 (g24014), .I2 (g3806));
ND2X1 gate20968(.O (g24477), .I1 (g24014), .I2 (g3806));
ND2X1 gate20969(.O (g24616), .I1 (g499), .I2 (g23376));
ND2X1 gate20970(.O (g24627), .I1 (g1186), .I2 (g23387));
ND2X1 gate20971(.O (g24641), .I1 (g1880), .I2 (g23394));
ND2X1 gate20972(.O (g24660), .I1 (g2574), .I2 (g23402));
ND2X1 gate20973(.O (I32265), .I1 (g17903), .I2 (g23936));
ND2X1 gate20974(.O (I32266), .I1 (g17903), .I2 (I32265));
ND2X1 gate20975(.O (I32267), .I1 (g23936), .I2 (I32265));
ND2X1 gate20976(.O (g24753), .I1 (I32266), .I2 (I32267));
ND2X1 gate20977(.O (I32284), .I1 (g17815), .I2 (g23953));
ND2X1 gate20978(.O (I32285), .I1 (g17815), .I2 (I32284));
ND2X1 gate20979(.O (I32286), .I1 (g23953), .I2 (I32284));
ND2X1 gate20980(.O (g24766), .I1 (I32285), .I2 (I32286));
ND2X1 gate20981(.O (I32295), .I1 (g18014), .I2 (g23968));
ND2X1 gate20982(.O (I32296), .I1 (g18014), .I2 (I32295));
ND2X1 gate20983(.O (I32297), .I1 (g23968), .I2 (I32295));
ND2X1 gate20984(.O (g24771), .I1 (I32296), .I2 (I32297));
ND2X1 gate20985(.O (I32308), .I1 (g17903), .I2 (g23973));
ND2X1 gate20986(.O (I32309), .I1 (g17903), .I2 (I32308));
ND2X1 gate20987(.O (I32310), .I1 (g23973), .I2 (I32308));
ND2X1 gate20988(.O (g24778), .I1 (I32309), .I2 (I32310));
ND2X1 gate20989(.O (I32323), .I1 (g17927), .I2 (g23982));
ND2X1 gate20990(.O (I32324), .I1 (g17927), .I2 (I32323));
ND2X1 gate20991(.O (I32325), .I1 (g23982), .I2 (I32323));
ND2X1 gate20992(.O (g24787), .I1 (I32324), .I2 (I32325));
ND2X1 gate20993(.O (I32333), .I1 (g18131), .I2 (g23997));
ND2X1 gate20994(.O (I32334), .I1 (g18131), .I2 (I32333));
ND2X1 gate20995(.O (I32335), .I1 (g23997), .I2 (I32333));
ND2X1 gate20996(.O (g24791), .I1 (I32334), .I2 (I32335));
ND2X1 gate20997(.O (I32345), .I1 (g17815), .I2 (g24002));
ND2X1 gate20998(.O (I32346), .I1 (g17815), .I2 (I32345));
ND2X1 gate20999(.O (I32347), .I1 (g24002), .I2 (I32345));
ND2X1 gate21000(.O (g24797), .I1 (I32346), .I2 (I32347));
ND2X1 gate21001(.O (I32355), .I1 (g18014), .I2 (g24003));
ND2X1 gate21002(.O (I32356), .I1 (g18014), .I2 (I32355));
ND2X1 gate21003(.O (I32357), .I1 (g24003), .I2 (I32355));
ND2X1 gate21004(.O (g24801), .I1 (I32356), .I2 (I32357));
ND2X1 gate21005(.O (I32368), .I1 (g18038), .I2 (g24012));
ND2X1 gate21006(.O (I32369), .I1 (g18038), .I2 (I32368));
ND2X1 gate21007(.O (I32370), .I1 (g24012), .I2 (I32368));
ND2X1 gate21008(.O (g24808), .I1 (I32369), .I2 (I32370));
ND2X1 gate21009(.O (I32378), .I1 (g18247), .I2 (g24027));
ND2X1 gate21010(.O (I32379), .I1 (g18247), .I2 (I32378));
ND2X1 gate21011(.O (I32380), .I1 (g24027), .I2 (I32378));
ND2X1 gate21012(.O (g24812), .I1 (I32379), .I2 (I32380));
ND2X1 gate21013(.O (g24814), .I1 (g24239), .I2 (g24244));
ND2X1 gate21014(.O (I32391), .I1 (g17903), .I2 (g24034));
ND2X1 gate21015(.O (I32392), .I1 (g17903), .I2 (I32391));
ND2X1 gate21016(.O (I32393), .I1 (g24034), .I2 (I32391));
ND2X1 gate21017(.O (g24817), .I1 (I32392), .I2 (I32393));
ND2X1 gate21018(.O (I32400), .I1 (g17927), .I2 (g24036));
ND2X1 gate21019(.O (I32401), .I1 (g17927), .I2 (I32400));
ND2X1 gate21020(.O (I32402), .I1 (g24036), .I2 (I32400));
ND2X1 gate21021(.O (g24820), .I1 (I32401), .I2 (I32402));
ND2X1 gate21022(.O (I32409), .I1 (g18131), .I2 (g24037));
ND2X1 gate21023(.O (I32410), .I1 (g18131), .I2 (I32409));
ND2X1 gate21024(.O (I32411), .I1 (g24037), .I2 (I32409));
ND2X1 gate21025(.O (g24823), .I1 (I32410), .I2 (I32411));
ND2X1 gate21026(.O (I32422), .I1 (g18155), .I2 (g24046));
ND2X1 gate21027(.O (I32423), .I1 (g18155), .I2 (I32422));
ND2X1 gate21028(.O (I32424), .I1 (g24046), .I2 (I32422));
ND2X1 gate21029(.O (g24830), .I1 (I32423), .I2 (I32424));
ND2X1 gate21030(.O (I32430), .I1 (g17815), .I2 (g24052));
ND2X1 gate21031(.O (I32431), .I1 (g17815), .I2 (I32430));
ND2X1 gate21032(.O (I32432), .I1 (g24052), .I2 (I32430));
ND2X1 gate21033(.O (g24832), .I1 (I32431), .I2 (I32432));
ND2X1 gate21034(.O (g24833), .I1 (g24245), .I2 (g24252));
ND2X1 gate21035(.O (I32443), .I1 (g18014), .I2 (g24054));
ND2X1 gate21036(.O (I32444), .I1 (g18014), .I2 (I32443));
ND2X1 gate21037(.O (I32445), .I1 (g24054), .I2 (I32443));
ND2X1 gate21038(.O (g24837), .I1 (I32444), .I2 (I32445));
ND2X1 gate21039(.O (I32451), .I1 (g18038), .I2 (g24056));
ND2X1 gate21040(.O (I32452), .I1 (g18038), .I2 (I32451));
ND2X1 gate21041(.O (I32453), .I1 (g24056), .I2 (I32451));
ND2X1 gate21042(.O (g24839), .I1 (I32452), .I2 (I32453));
ND2X1 gate21043(.O (I32460), .I1 (g18247), .I2 (g24057));
ND2X1 gate21044(.O (I32461), .I1 (g18247), .I2 (I32460));
ND2X1 gate21045(.O (I32462), .I1 (g24057), .I2 (I32460));
ND2X1 gate21046(.O (g24842), .I1 (I32461), .I2 (I32462));
ND2X1 gate21047(.O (I32468), .I1 (g17903), .I2 (g24058));
ND2X1 gate21048(.O (I32469), .I1 (g17903), .I2 (I32468));
ND2X1 gate21049(.O (I32470), .I1 (g24058), .I2 (I32468));
ND2X1 gate21050(.O (g24844), .I1 (I32469), .I2 (I32470));
ND2X1 gate21051(.O (I32478), .I1 (g17927), .I2 (g24065));
ND2X1 gate21052(.O (I32479), .I1 (g17927), .I2 (I32478));
ND2X1 gate21053(.O (I32480), .I1 (g24065), .I2 (I32478));
ND2X1 gate21054(.O (g24848), .I1 (I32479), .I2 (I32480));
ND2X1 gate21055(.O (g24849), .I1 (g24254), .I2 (g24257));
ND2X1 gate21056(.O (I32490), .I1 (g18131), .I2 (g24067));
ND2X1 gate21057(.O (I32491), .I1 (g18131), .I2 (I32490));
ND2X1 gate21058(.O (I32492), .I1 (g24067), .I2 (I32490));
ND2X1 gate21059(.O (g24852), .I1 (I32491), .I2 (I32492));
ND2X1 gate21060(.O (I32498), .I1 (g18155), .I2 (g24069));
ND2X1 gate21061(.O (I32499), .I1 (g18155), .I2 (I32498));
ND2X1 gate21062(.O (I32500), .I1 (g24069), .I2 (I32498));
ND2X1 gate21063(.O (g24854), .I1 (I32499), .I2 (I32500));
ND2X1 gate21064(.O (I32509), .I1 (g17815), .I2 (g24070));
ND2X1 gate21065(.O (I32510), .I1 (g17815), .I2 (I32509));
ND2X1 gate21066(.O (I32511), .I1 (g24070), .I2 (I32509));
ND2X1 gate21067(.O (g24857), .I1 (I32510), .I2 (I32511));
ND2X1 gate21068(.O (I32518), .I1 (g18014), .I2 (g24071));
ND2X1 gate21069(.O (I32519), .I1 (g18014), .I2 (I32518));
ND2X1 gate21070(.O (I32520), .I1 (g24071), .I2 (I32518));
ND2X1 gate21071(.O (g24860), .I1 (I32519), .I2 (I32520));
ND2X1 gate21072(.O (I32526), .I1 (g18038), .I2 (g24078));
ND2X1 gate21073(.O (I32527), .I1 (g18038), .I2 (I32526));
ND2X1 gate21074(.O (I32528), .I1 (g24078), .I2 (I32526));
ND2X1 gate21075(.O (g24862), .I1 (I32527), .I2 (I32528));
ND2X1 gate21076(.O (g24863), .I1 (g24258), .I2 (g23319));
ND2X1 gate21077(.O (I32538), .I1 (g18247), .I2 (g24080));
ND2X1 gate21078(.O (I32539), .I1 (g18247), .I2 (I32538));
ND2X1 gate21079(.O (I32540), .I1 (g24080), .I2 (I32538));
ND2X1 gate21080(.O (g24866), .I1 (I32539), .I2 (I32540));
ND2X1 gate21081(.O (I32546), .I1 (g17903), .I2 (g23906));
ND2X1 gate21082(.O (I32547), .I1 (g17903), .I2 (I32546));
ND2X1 gate21083(.O (I32548), .I1 (g23906), .I2 (I32546));
ND2X1 gate21084(.O (g24868), .I1 (I32547), .I2 (I32548));
ND2X1 gate21085(.O (I32559), .I1 (g17927), .I2 (g24081));
ND2X1 gate21086(.O (I32560), .I1 (g17927), .I2 (I32559));
ND2X1 gate21087(.O (I32561), .I1 (g24081), .I2 (I32559));
ND2X1 gate21088(.O (g24873), .I1 (I32560), .I2 (I32561));
ND2X1 gate21089(.O (I32567), .I1 (g18131), .I2 (g24082));
ND2X1 gate21090(.O (I32568), .I1 (g18131), .I2 (I32567));
ND2X1 gate21091(.O (I32569), .I1 (g24082), .I2 (I32567));
ND2X1 gate21092(.O (g24875), .I1 (I32568), .I2 (I32569));
ND2X1 gate21093(.O (I32575), .I1 (g18155), .I2 (g24089));
ND2X1 gate21094(.O (I32576), .I1 (g18155), .I2 (I32575));
ND2X1 gate21095(.O (I32577), .I1 (g24089), .I2 (I32575));
ND2X1 gate21096(.O (g24877), .I1 (I32576), .I2 (I32577));
ND2X1 gate21097(.O (I32586), .I1 (g17815), .I2 (g23937));
ND2X1 gate21098(.O (I32587), .I1 (g17815), .I2 (I32586));
ND2X1 gate21099(.O (I32588), .I1 (g23937), .I2 (I32586));
ND2X1 gate21100(.O (g24880), .I1 (I32587), .I2 (I32588));
ND2X1 gate21101(.O (I32595), .I1 (g18014), .I2 (g23938));
ND2X1 gate21102(.O (I32596), .I1 (g18014), .I2 (I32595));
ND2X1 gate21103(.O (I32597), .I1 (g23938), .I2 (I32595));
ND2X1 gate21104(.O (g24883), .I1 (I32596), .I2 (I32597));
ND2X1 gate21105(.O (I32607), .I1 (g18038), .I2 (g24090));
ND2X1 gate21106(.O (I32608), .I1 (g18038), .I2 (I32607));
ND2X1 gate21107(.O (I32609), .I1 (g24090), .I2 (I32607));
ND2X1 gate21108(.O (g24887), .I1 (I32608), .I2 (I32609));
ND2X1 gate21109(.O (I32615), .I1 (g18247), .I2 (g24091));
ND2X1 gate21110(.O (I32616), .I1 (g18247), .I2 (I32615));
ND2X1 gate21111(.O (I32617), .I1 (g24091), .I2 (I32615));
ND2X1 gate21112(.O (g24889), .I1 (I32616), .I2 (I32617));
ND2X1 gate21113(.O (I32624), .I1 (g17927), .I2 (g23969));
ND2X1 gate21114(.O (I32625), .I1 (g17927), .I2 (I32624));
ND2X1 gate21115(.O (I32626), .I1 (g23969), .I2 (I32624));
ND2X1 gate21116(.O (g24897), .I1 (I32625), .I2 (I32626));
ND2X1 gate21117(.O (I32633), .I1 (g18131), .I2 (g23970));
ND2X1 gate21118(.O (I32634), .I1 (g18131), .I2 (I32633));
ND2X1 gate21119(.O (I32635), .I1 (g23970), .I2 (I32633));
ND2X1 gate21120(.O (g24900), .I1 (I32634), .I2 (I32635));
ND2X1 gate21121(.O (I32645), .I1 (g18155), .I2 (g24093));
ND2X1 gate21122(.O (I32646), .I1 (g18155), .I2 (I32645));
ND2X1 gate21123(.O (I32647), .I1 (g24093), .I2 (I32645));
ND2X1 gate21124(.O (g24904), .I1 (I32646), .I2 (I32647));
ND2X1 gate21125(.O (I32659), .I1 (g18038), .I2 (g23998));
ND2X1 gate21126(.O (I32660), .I1 (g18038), .I2 (I32659));
ND2X1 gate21127(.O (I32661), .I1 (g23998), .I2 (I32659));
ND2X1 gate21128(.O (g24920), .I1 (I32660), .I2 (I32661));
ND2X1 gate21129(.O (I32668), .I1 (g18247), .I2 (g23999));
ND2X1 gate21130(.O (I32669), .I1 (g18247), .I2 (I32668));
ND2X1 gate21131(.O (I32670), .I1 (g23999), .I2 (I32668));
ND2X1 gate21132(.O (g24923), .I1 (I32669), .I2 (I32670));
ND2X1 gate21133(.O (I32677), .I1 (g23823), .I2 (g14165));
ND2X1 gate21134(.O (I32678), .I1 (g23823), .I2 (I32677));
ND2X1 gate21135(.O (I32679), .I1 (g14165), .I2 (I32677));
ND2X1 gate21136(.O (g24928), .I1 (I32678), .I2 (I32679));
ND2X1 gate21137(.O (I32686), .I1 (g18155), .I2 (g24028));
ND2X1 gate21138(.O (I32687), .I1 (g18155), .I2 (I32686));
ND2X1 gate21139(.O (I32688), .I1 (g24028), .I2 (I32686));
ND2X1 gate21140(.O (g24937), .I1 (I32687), .I2 (I32688));
ND2X1 gate21141(.O (I32695), .I1 (g23858), .I2 (g14280));
ND2X1 gate21142(.O (I32696), .I1 (g23858), .I2 (I32695));
ND2X1 gate21143(.O (I32697), .I1 (g14280), .I2 (I32695));
ND2X1 gate21144(.O (g24940), .I1 (I32696), .I2 (I32697));
ND2X1 gate21145(.O (I32708), .I1 (g23892), .I2 (g14402));
ND2X1 gate21146(.O (I32709), .I1 (g23892), .I2 (I32708));
ND2X1 gate21147(.O (I32710), .I1 (g14402), .I2 (I32708));
ND2X1 gate21148(.O (g24951), .I1 (I32709), .I2 (I32710));
ND2X1 gate21149(.O (I32724), .I1 (g23913), .I2 (g14514));
ND2X1 gate21150(.O (I32725), .I1 (g23913), .I2 (I32724));
ND2X1 gate21151(.O (I32726), .I1 (g14514), .I2 (I32724));
ND2X1 gate21152(.O (g24963), .I1 (I32725), .I2 (I32726));
ND2X1 gate21153(.O (g24975), .I1 (g23497), .I2 (g74));
ND2X1 gate21154(.O (g24986), .I1 (g23513), .I2 (g762));
ND2X1 gate21155(.O (g24997), .I1 (g23528), .I2 (g1448));
ND2X1 gate21156(.O (g25004), .I1 (g23644), .I2 (g6448));
ND2X1 gate21157(.O (g25005), .I1 (g23539), .I2 (g2142));
ND2X1 gate21158(.O (g25008), .I1 (g23644), .I2 (g5438));
ND2X1 gate21159(.O (g25009), .I1 (g23644), .I2 (g6448));
ND2X1 gate21160(.O (g25010), .I1 (g23694), .I2 (g6713));
ND2X1 gate21161(.O (g25011), .I1 (g23644), .I2 (g5438));
ND2X1 gate21162(.O (g25012), .I1 (g23644), .I2 (g6448));
ND2X1 gate21163(.O (g25013), .I1 (g23923), .I2 (g6643));
ND2X1 gate21164(.O (g25014), .I1 (g23694), .I2 (g5473));
ND2X1 gate21165(.O (g25015), .I1 (g23694), .I2 (g6713));
ND2X1 gate21166(.O (g25016), .I1 (g23748), .I2 (g7015));
ND2X1 gate21167(.O (g25017), .I1 (g23644), .I2 (g5438));
ND2X1 gate21168(.O (g25018), .I1 (g23644), .I2 (g6448));
ND2X1 gate21169(.O (g25019), .I1 (g23923), .I2 (g6486));
ND2X1 gate21170(.O (g25020), .I1 (g23923), .I2 (g6643));
ND2X1 gate21171(.O (g25021), .I1 (g23694), .I2 (g5473));
ND2X1 gate21172(.O (g25022), .I1 (g23694), .I2 (g6713));
ND2X1 gate21173(.O (g25023), .I1 (g23955), .I2 (g6945));
ND2X1 gate21174(.O (g25024), .I1 (g23748), .I2 (g5512));
ND2X1 gate21175(.O (g25025), .I1 (g23748), .I2 (g7015));
ND2X1 gate21176(.O (g25026), .I1 (g23803), .I2 (g7265));
ND2X1 gate21177(.O (g25028), .I1 (g23644), .I2 (g5438));
ND2X1 gate21178(.O (g25029), .I1 (g23923), .I2 (g6486));
ND2X1 gate21179(.O (g25030), .I1 (g23923), .I2 (g6643));
ND2X1 gate21180(.O (g25031), .I1 (g23694), .I2 (g5473));
ND2X1 gate21181(.O (g25032), .I1 (g23694), .I2 (g6713));
ND2X1 gate21182(.O (g25033), .I1 (g23955), .I2 (g6751));
ND2X1 gate21183(.O (g25034), .I1 (g23955), .I2 (g6945));
ND2X1 gate21184(.O (g25035), .I1 (g23748), .I2 (g5512));
ND2X1 gate21185(.O (g25036), .I1 (g23748), .I2 (g7015));
ND2X1 gate21186(.O (g25037), .I1 (g23984), .I2 (g7195));
ND2X1 gate21187(.O (g25038), .I1 (g23803), .I2 (g5556));
ND2X1 gate21188(.O (g25039), .I1 (g23803), .I2 (g7265));
ND2X1 gate21189(.O (g25040), .I1 (g23923), .I2 (g6486));
ND2X1 gate21190(.O (g25041), .I1 (g23923), .I2 (g6643));
ND2X1 gate21191(.O (g25043), .I1 (g23694), .I2 (g5473));
ND2X1 gate21192(.O (g25044), .I1 (g23955), .I2 (g6751));
ND2X1 gate21193(.O (g25045), .I1 (g23955), .I2 (g6945));
ND2X1 gate21194(.O (g25046), .I1 (g23748), .I2 (g5512));
ND2X1 gate21195(.O (g25047), .I1 (g23748), .I2 (g7015));
ND2X1 gate21196(.O (g25048), .I1 (g23984), .I2 (g7053));
ND2X1 gate21197(.O (g25049), .I1 (g23984), .I2 (g7195));
ND2X1 gate21198(.O (g25050), .I1 (g23803), .I2 (g5556));
ND2X1 gate21199(.O (g25051), .I1 (g23803), .I2 (g7265));
ND2X1 gate21200(.O (g25052), .I1 (g24014), .I2 (g7391));
ND2X1 gate21201(.O (g25053), .I1 (g23923), .I2 (g6486));
ND2X1 gate21202(.O (g25054), .I1 (g23955), .I2 (g6751));
ND2X1 gate21203(.O (g25055), .I1 (g23955), .I2 (g6945));
ND2X1 gate21204(.O (g25057), .I1 (g23748), .I2 (g5512));
ND2X1 gate21205(.O (g25058), .I1 (g23984), .I2 (g7053));
ND2X1 gate21206(.O (g25059), .I1 (g23984), .I2 (g7195));
ND2X1 gate21207(.O (g25060), .I1 (g23803), .I2 (g5556));
ND2X1 gate21208(.O (g25061), .I1 (g23803), .I2 (g7265));
ND2X1 gate21209(.O (g25062), .I1 (g24014), .I2 (g7303));
ND2X1 gate21210(.O (g25063), .I1 (g24014), .I2 (g7391));
ND2X1 gate21211(.O (g25064), .I1 (g23955), .I2 (g6751));
ND2X1 gate21212(.O (g25065), .I1 (g23984), .I2 (g7053));
ND2X1 gate21213(.O (g25066), .I1 (g23984), .I2 (g7195));
ND2X1 gate21214(.O (g25068), .I1 (g23803), .I2 (g5556));
ND2X1 gate21215(.O (g25069), .I1 (g24014), .I2 (g7303));
ND2X1 gate21216(.O (g25070), .I1 (g24014), .I2 (g7391));
ND2X1 gate21217(.O (g25071), .I1 (g23984), .I2 (g7053));
ND2X1 gate21218(.O (g25072), .I1 (g24014), .I2 (g7303));
ND2X1 gate21219(.O (g25073), .I1 (g24014), .I2 (g7391));
ND2X1 gate21220(.O (g25074), .I1 (g24014), .I2 (g7303));
ND2X1 gate21221(.O (g25088), .I1 (g23950), .I2 (g679));
ND2X1 gate21222(.O (g25096), .I1 (g23979), .I2 (g1365));
ND2X1 gate21223(.O (g25106), .I1 (g24009), .I2 (g2059));
ND2X1 gate21224(.O (g25112), .I1 (g24043), .I2 (g2753));
ND2X1 gate21225(.O (g25200), .I1 (g24965), .I2 (g3306));
ND2X1 gate21226(.O (g25203), .I1 (g24978), .I2 (g3462));
ND2X1 gate21227(.O (g25205), .I1 (g24989), .I2 (g3618));
ND2X1 gate21228(.O (g25210), .I1 (g25000), .I2 (g3774));
ND4X1 gate21229(.O (g25312), .I1 (g21211), .I2 (g14442), .I3 (g10694), .I4 (g24590));
ND4X1 gate21230(.O (g25320), .I1 (g21219), .I2 (g14529), .I3 (g10714), .I4 (g24595));
ND4X1 gate21231(.O (g25331), .I1 (g21230), .I2 (g14584), .I3 (g10735), .I4 (g24603));
ND4X1 gate21232(.O (g25340), .I1 (g21235), .I2 (g14618), .I3 (g10754), .I4 (g24610));
ND2X1 gate21233(.O (g25927), .I1 (g24965), .I2 (g6448));
ND2X1 gate21234(.O (g25928), .I1 (g24965), .I2 (g5438));
ND2X1 gate21235(.O (g25929), .I1 (g24978), .I2 (g6713));
ND2X1 gate21236(.O (g25930), .I1 (g24978), .I2 (g5473));
ND2X1 gate21237(.O (g25931), .I1 (g24989), .I2 (g7015));
ND2X1 gate21238(.O (g25933), .I1 (g24989), .I2 (g5512));
ND2X1 gate21239(.O (g25934), .I1 (g25000), .I2 (g7265));
ND2X1 gate21240(.O (g25936), .I1 (g25000), .I2 (g5556));
ND2X1 gate21241(.O (g25954), .I1 (g22806), .I2 (g24517));
ND2X1 gate21242(.O (g25958), .I1 (g22847), .I2 (g24530));
ND2X1 gate21243(.O (g25964), .I1 (g22882), .I2 (g24543));
ND2X1 gate21244(.O (g25969), .I1 (g22917), .I2 (g24555));
ND3X1 gate21245(.O (g26059), .I1 (g25422), .I2 (g25379), .I3 (g25274));
ND3X1 gate21246(.O (g26066), .I1 (g25431), .I2 (g25395), .I3 (g25283));
ND3X1 gate21247(.O (g26073), .I1 (g25438), .I2 (g25405), .I3 (g25291));
ND3X1 gate21248(.O (g26079), .I1 (g25445), .I2 (g25413), .I3 (g25301));
ND2X1 gate21249(.O (g26106), .I1 (g23644), .I2 (g25354));
ND4X1 gate21250(.O (g26119), .I1 (g8278), .I2 (g14657), .I3 (g25422), .I4 (g25379));
ND2X1 gate21251(.O (g26120), .I1 (g23694), .I2 (g25369));
ND4X1 gate21252(.O (g26129), .I1 (g8287), .I2 (g14691), .I3 (g25431), .I4 (g25395));
ND2X1 gate21253(.O (g26130), .I1 (g23748), .I2 (g25386));
ND4X1 gate21254(.O (g26143), .I1 (g8296), .I2 (g14725), .I3 (g25438), .I4 (g25405));
ND2X1 gate21255(.O (g26144), .I1 (g23803), .I2 (g25402));
ND4X1 gate21256(.O (g26148), .I1 (g8305), .I2 (g14753), .I3 (g25445), .I4 (g25413));
ND2X1 gate21257(.O (g26356), .I1 (g16539), .I2 (g25183));
ND2X1 gate21258(.O (g26399), .I1 (g16571), .I2 (g25186));
ND2X1 gate21259(.O (g26440), .I1 (g16595), .I2 (g25190));
ND2X1 gate21260(.O (g26458), .I1 (g25343), .I2 (g65));
ND2X1 gate21261(.O (g26472), .I1 (g16615), .I2 (g25195));
ND2X1 gate21262(.O (g26482), .I1 (g25357), .I2 (g753));
ND2X1 gate21263(.O (g26498), .I1 (g25372), .I2 (g1439));
ND2X1 gate21264(.O (g26513), .I1 (g25389), .I2 (g2133));
ND2X1 gate21265(.O (g26772), .I1 (g26320), .I2 (g3306));
ND2X1 gate21266(.O (g26779), .I1 (g26367), .I2 (g3462));
ND2X1 gate21267(.O (g26785), .I1 (g26410), .I2 (g3618));
ND2X1 gate21268(.O (g26792), .I1 (g26451), .I2 (g3774));
ND2X1 gate21269(.O (I35020), .I1 (g26110), .I2 (g26099));
ND2X1 gate21270(.O (I35021), .I1 (g26110), .I2 (I35020));
ND2X1 gate21271(.O (I35022), .I1 (g26099), .I2 (I35020));
ND2X1 gate21272(.O (g26859), .I1 (I35021), .I2 (I35022));
ND2X1 gate21273(.O (I35034), .I1 (g26087), .I2 (g26154));
ND2X1 gate21274(.O (I35035), .I1 (g26087), .I2 (I35034));
ND2X1 gate21275(.O (I35036), .I1 (g26154), .I2 (I35034));
ND2X1 gate21276(.O (g26865), .I1 (I35035), .I2 (I35036));
ND2X1 gate21277(.O (I35042), .I1 (g26151), .I2 (g26145));
ND2X1 gate21278(.O (I35043), .I1 (g26151), .I2 (I35042));
ND2X1 gate21279(.O (I35044), .I1 (g26145), .I2 (I35042));
ND2X1 gate21280(.O (g26867), .I1 (I35043), .I2 (I35044));
ND2X1 gate21281(.O (I35057), .I1 (g26137), .I2 (g26126));
ND2X1 gate21282(.O (I35058), .I1 (g26137), .I2 (I35057));
ND2X1 gate21283(.O (I35059), .I1 (g26126), .I2 (I35057));
ND2X1 gate21284(.O (g26874), .I1 (I35058), .I2 (I35059));
ND4X1 gate21285(.O (g26892), .I1 (g25699), .I2 (g26283), .I3 (g25569), .I4 (g25631));
ND3X1 gate21286(.O (g26902), .I1 (g25631), .I2 (g26283), .I3 (g25569));
ND4X1 gate21287(.O (g26906), .I1 (g25772), .I2 (g26327), .I3 (g25648), .I4 (g25708));
ND2X1 gate21288(.O (g26911), .I1 (g25569), .I2 (g26283));
ND3X1 gate21289(.O (g26915), .I1 (g25708), .I2 (g26327), .I3 (g25648));
ND4X1 gate21290(.O (g26918), .I1 (g25826), .I2 (g26374), .I3 (g25725), .I4 (g25781));
ND2X1 gate21291(.O (g26925), .I1 (g25648), .I2 (g26327));
ND3X1 gate21292(.O (g26928), .I1 (g25781), .I2 (g26374), .I3 (g25725));
ND4X1 gate21293(.O (g26931), .I1 (g25861), .I2 (g26417), .I3 (g25798), .I4 (g25835));
ND2X1 gate21294(.O (I35123), .I1 (g26107), .I2 (g26096));
ND2X1 gate21295(.O (I35124), .I1 (g26107), .I2 (I35123));
ND2X1 gate21296(.O (I35125), .I1 (g26096), .I2 (I35123));
ND2X1 gate21297(.O (g26934), .I1 (I35124), .I2 (I35125));
ND2X1 gate21298(.O (g26938), .I1 (g25725), .I2 (g26374));
ND3X1 gate21299(.O (g26941), .I1 (g25835), .I2 (g26417), .I3 (g25798));
ND2X1 gate21300(.O (g26947), .I1 (g25798), .I2 (g26417));
ND2X1 gate21301(.O (g27117), .I1 (g26320), .I2 (g6448));
ND2X1 gate21302(.O (g27118), .I1 (g26320), .I2 (g5438));
ND2X1 gate21303(.O (g27119), .I1 (g26367), .I2 (g6713));
ND2X1 gate21304(.O (g27121), .I1 (g26367), .I2 (g5473));
ND2X1 gate21305(.O (g27122), .I1 (g26410), .I2 (g7015));
ND2X1 gate21306(.O (g27124), .I1 (g26410), .I2 (g5512));
ND2X1 gate21307(.O (g27125), .I1 (g26451), .I2 (g7265));
ND2X1 gate21308(.O (g27130), .I1 (g26451), .I2 (g5556));
ND2X1 gate21309(.O (I35701), .I1 (g26867), .I2 (g26874));
ND2X1 gate21310(.O (I35702), .I1 (g26867), .I2 (I35701));
ND2X1 gate21311(.O (I35703), .I1 (g26874), .I2 (I35701));
ND2X1 gate21312(.O (g27379), .I1 (I35702), .I2 (I35703));
ND2X1 gate21313(.O (I35714), .I1 (g26859), .I2 (g26865));
ND2X1 gate21314(.O (I35715), .I1 (g26859), .I2 (I35714));
ND2X1 gate21315(.O (I35716), .I1 (g26865), .I2 (I35714));
ND2X1 gate21316(.O (g27382), .I1 (I35715), .I2 (I35716));
ND2X1 gate21317(.O (g27390), .I1 (g26989), .I2 (g6448));
ND2X1 gate21318(.O (g27395), .I1 (g26989), .I2 (g5438));
ND2X1 gate21319(.O (g27400), .I1 (g27012), .I2 (g6713));
ND2X1 gate21320(.O (g27408), .I1 (g27012), .I2 (g5473));
ND2X1 gate21321(.O (g27413), .I1 (g27038), .I2 (g7015));
ND2X1 gate21322(.O (g27426), .I1 (g27038), .I2 (g5512));
ND2X1 gate21323(.O (g27431), .I1 (g27066), .I2 (g7265));
ND2X1 gate21324(.O (g27447), .I1 (g27066), .I2 (g5556));
ND2X1 gate21325(.O (I35904), .I1 (g27051), .I2 (g14831));
ND2X1 gate21326(.O (I35905), .I1 (g27051), .I2 (I35904));
ND2X1 gate21327(.O (I35906), .I1 (g14831), .I2 (I35904));
ND2X1 gate21328(.O (g27528), .I1 (I35905), .I2 (I35906));
ND2X1 gate21329(.O (I35944), .I1 (g27078), .I2 (g14904));
ND2X1 gate21330(.O (I35945), .I1 (g27078), .I2 (I35944));
ND2X1 gate21331(.O (I35946), .I1 (g14904), .I2 (I35944));
ND2X1 gate21332(.O (g27550), .I1 (I35945), .I2 (I35946));
ND2X1 gate21333(.O (I35974), .I1 (g27094), .I2 (g14985));
ND2X1 gate21334(.O (I35975), .I1 (g27094), .I2 (I35974));
ND2X1 gate21335(.O (I35976), .I1 (g14985), .I2 (I35974));
ND2X1 gate21336(.O (g27566), .I1 (I35975), .I2 (I35976));
ND2X1 gate21337(.O (g27571), .I1 (g26869), .I2 (g56));
ND2X1 gate21338(.O (I35992), .I1 (g27106), .I2 (g15074));
ND2X1 gate21339(.O (I35993), .I1 (g27106), .I2 (I35992));
ND2X1 gate21340(.O (I35994), .I1 (g15074), .I2 (I35992));
ND2X1 gate21341(.O (g27576), .I1 (I35993), .I2 (I35994));
ND2X1 gate21342(.O (g27580), .I1 (g26878), .I2 (g744));
ND2X1 gate21343(.O (g27583), .I1 (g26887), .I2 (g1430));
ND2X1 gate21344(.O (g27587), .I1 (g26897), .I2 (g2124));
ND2X1 gate21345(.O (g27626), .I1 (g26989), .I2 (g3306));
ND2X1 gate21346(.O (g27627), .I1 (g27012), .I2 (g3462));
ND2X1 gate21347(.O (g27628), .I1 (g27038), .I2 (g3618));
ND2X1 gate21348(.O (g27630), .I1 (g27066), .I2 (g3774));
ND2X1 gate21349(.O (g27738), .I1 (g25367), .I2 (g27415));
ND2X1 gate21350(.O (g27743), .I1 (g25384), .I2 (g27436));
ND2X1 gate21351(.O (g27751), .I1 (g25400), .I2 (g27455));
ND2X1 gate21352(.O (g27756), .I1 (g25410), .I2 (g27471));
ND2X1 gate21353(.O (I36256), .I1 (g27527), .I2 (g15859));
ND2X1 gate21354(.O (I36257), .I1 (g27527), .I2 (I36256));
ND2X1 gate21355(.O (I36258), .I1 (g15859), .I2 (I36256));
ND2X1 gate21356(.O (g27801), .I1 (I36257), .I2 (I36258));
ND2X1 gate21357(.O (I36270), .I1 (g27549), .I2 (g15890));
ND2X1 gate21358(.O (I36271), .I1 (g27549), .I2 (I36270));
ND2X1 gate21359(.O (I36272), .I1 (g15890), .I2 (I36270));
ND2X1 gate21360(.O (g27809), .I1 (I36271), .I2 (I36272));
ND2X1 gate21361(.O (I36289), .I1 (g27565), .I2 (g15923));
ND2X1 gate21362(.O (I36290), .I1 (g27565), .I2 (I36289));
ND2X1 gate21363(.O (I36291), .I1 (g15923), .I2 (I36289));
ND2X1 gate21364(.O (g27830), .I1 (I36290), .I2 (I36291));
ND2X1 gate21365(.O (I36300), .I1 (g27382), .I2 (g27379));
ND2X1 gate21366(.O (I36301), .I1 (g27382), .I2 (I36300));
ND2X1 gate21367(.O (I36302), .I1 (g27379), .I2 (I36300));
ND2X1 gate21368(.O (g27838), .I1 (I36301), .I2 (I36302));
ND2X1 gate21369(.O (I36314), .I1 (g27575), .I2 (g15952));
ND2X1 gate21370(.O (I36315), .I1 (g27575), .I2 (I36314));
ND2X1 gate21371(.O (I36316), .I1 (g15952), .I2 (I36314));
ND2X1 gate21372(.O (g27846), .I1 (I36315), .I2 (I36316));
ND2X1 gate21373(.O (I36591), .I1 (g27529), .I2 (g14885));
ND2X1 gate21374(.O (I36592), .I1 (g27529), .I2 (I36591));
ND2X1 gate21375(.O (I36593), .I1 (g14885), .I2 (I36591));
ND2X1 gate21376(.O (g28046), .I1 (I36592), .I2 (I36593));
ND2X1 gate21377(.O (I36666), .I1 (g27551), .I2 (g14966));
ND2X1 gate21378(.O (I36667), .I1 (g27551), .I2 (I36666));
ND2X1 gate21379(.O (I36668), .I1 (g14966), .I2 (I36666));
ND2X1 gate21380(.O (g28075), .I1 (I36667), .I2 (I36668));
ND2X1 gate21381(.O (I36731), .I1 (g27567), .I2 (g15055));
ND2X1 gate21382(.O (I36732), .I1 (g27567), .I2 (I36731));
ND2X1 gate21383(.O (I36733), .I1 (g15055), .I2 (I36731));
ND2X1 gate21384(.O (g28100), .I1 (I36732), .I2 (I36733));
ND2X1 gate21385(.O (I36779), .I1 (g27577), .I2 (g15151));
ND2X1 gate21386(.O (I36780), .I1 (g27577), .I2 (I36779));
ND2X1 gate21387(.O (I36781), .I1 (g15151), .I2 (I36779));
ND2X1 gate21388(.O (g28118), .I1 (I36780), .I2 (I36781));
ND2X1 gate21389(.O (I37295), .I1 (g27827), .I2 (g27814));
ND2X1 gate21390(.O (I37296), .I1 (g27827), .I2 (I37295));
ND2X1 gate21391(.O (I37297), .I1 (g27814), .I2 (I37295));
ND2X1 gate21392(.O (g28384), .I1 (I37296), .I2 (I37297));
ND2X1 gate21393(.O (I37303), .I1 (g27802), .I2 (g27900));
ND2X1 gate21394(.O (I37304), .I1 (g27802), .I2 (I37303));
ND2X1 gate21395(.O (I37305), .I1 (g27900), .I2 (I37303));
ND2X1 gate21396(.O (g28386), .I1 (I37304), .I2 (I37305));
ND2X1 gate21397(.O (I37311), .I1 (g27897), .I2 (g27883));
ND2X1 gate21398(.O (I37312), .I1 (g27897), .I2 (I37311));
ND2X1 gate21399(.O (I37313), .I1 (g27883), .I2 (I37311));
ND2X1 gate21400(.O (g28388), .I1 (I37312), .I2 (I37313));
ND2X1 gate21401(.O (I37322), .I1 (g27865), .I2 (g27855));
ND2X1 gate21402(.O (I37323), .I1 (g27865), .I2 (I37322));
ND2X1 gate21403(.O (I37324), .I1 (g27855), .I2 (I37322));
ND2X1 gate21404(.O (g28391), .I1 (I37323), .I2 (I37324));
ND2X1 gate21405(.O (I37356), .I1 (g27824), .I2 (g27811));
ND2X1 gate21406(.O (I37357), .I1 (g27824), .I2 (I37356));
ND2X1 gate21407(.O (I37358), .I1 (g27811), .I2 (I37356));
ND2X1 gate21408(.O (g28415), .I1 (I37357), .I2 (I37358));
ND2X1 gate21409(.O (I37813), .I1 (g28388), .I2 (g28391));
ND2X1 gate21410(.O (I37814), .I1 (g28388), .I2 (I37813));
ND2X1 gate21411(.O (I37815), .I1 (g28391), .I2 (I37813));
ND2X1 gate21412(.O (g28842), .I1 (I37814), .I2 (I37815));
ND2X1 gate21413(.O (I37822), .I1 (g28384), .I2 (g28386));
ND2X1 gate21414(.O (I37823), .I1 (g28384), .I2 (I37822));
ND2X1 gate21415(.O (I37824), .I1 (g28386), .I2 (I37822));
ND2X1 gate21416(.O (g28845), .I1 (I37823), .I2 (I37824));
ND2X1 gate21417(.O (g28978), .I1 (g9150), .I2 (g28512));
ND2X1 gate21418(.O (g29001), .I1 (g9161), .I2 (g28512));
ND2X1 gate21419(.O (g29008), .I1 (g9174), .I2 (g28540));
ND2X1 gate21420(.O (g29026), .I1 (g9187), .I2 (g28512));
ND2X1 gate21421(.O (g29030), .I1 (g9203), .I2 (g28540));
ND2X1 gate21422(.O (g29038), .I1 (g9216), .I2 (g28567));
ND2X1 gate21423(.O (g29045), .I1 (g9232), .I2 (g28512));
ND2X1 gate21424(.O (g29049), .I1 (g9248), .I2 (g28540));
ND2X1 gate21425(.O (g29053), .I1 (g9264), .I2 (g28567));
ND2X1 gate21426(.O (g29060), .I1 (g9277), .I2 (g28595));
ND2X1 gate21427(.O (g29062), .I1 (g9310), .I2 (g28540));
ND2X1 gate21428(.O (g29068), .I1 (g9326), .I2 (g28567));
ND2X1 gate21429(.O (g29072), .I1 (g9342), .I2 (g28595));
ND2X1 gate21430(.O (g29076), .I1 (g9391), .I2 (g28567));
ND2X1 gate21431(.O (g29080), .I1 (g9407), .I2 (g28595));
ND2X1 gate21432(.O (g29087), .I1 (g9488), .I2 (g28595));
ND2X1 gate21433(.O (g29088), .I1 (g9507), .I2 (g28512));
ND2X1 gate21434(.O (g29096), .I1 (g9649), .I2 (g28540));
ND2X1 gate21435(.O (g29103), .I1 (g9795), .I2 (g28567));
ND2X1 gate21436(.O (g29107), .I1 (g9941), .I2 (g28595));
ND2X1 gate21437(.O (I38378), .I1 (g28845), .I2 (g28842));
ND2X1 gate21438(.O (I38379), .I1 (g28845), .I2 (I38378));
ND2X1 gate21439(.O (I38380), .I1 (g28842), .I2 (I38378));
ND2X1 gate21440(.O (g29265), .I1 (I38379), .I2 (I38380));
ND2X1 gate21441(.O (I38810), .I1 (g29303), .I2 (g15904));
ND2X1 gate21442(.O (I38811), .I1 (g29303), .I2 (I38810));
ND2X1 gate21443(.O (I38812), .I1 (g15904), .I2 (I38810));
ND2X1 gate21444(.O (g29498), .I1 (I38811), .I2 (I38812));
ND2X1 gate21445(.O (I38820), .I1 (g29313), .I2 (g15933));
ND2X1 gate21446(.O (I38821), .I1 (g29313), .I2 (I38820));
ND2X1 gate21447(.O (I38822), .I1 (g15933), .I2 (I38820));
ND2X1 gate21448(.O (g29500), .I1 (I38821), .I2 (I38822));
ND2X1 gate21449(.O (I38831), .I1 (g29324), .I2 (g15962));
ND2X1 gate21450(.O (I38832), .I1 (g29324), .I2 (I38831));
ND2X1 gate21451(.O (I38833), .I1 (g15962), .I2 (I38831));
ND2X1 gate21452(.O (g29503), .I1 (I38832), .I2 (I38833));
ND2X1 gate21453(.O (I38841), .I1 (g29333), .I2 (g15981));
ND2X1 gate21454(.O (I38842), .I1 (g29333), .I2 (I38841));
ND2X1 gate21455(.O (I38843), .I1 (g15981), .I2 (I38841));
ND2X1 gate21456(.O (g29505), .I1 (I38842), .I2 (I38843));
ND2X1 gate21457(.O (I39323), .I1 (g29721), .I2 (g29713));
ND2X1 gate21458(.O (I39324), .I1 (g29721), .I2 (I39323));
ND2X1 gate21459(.O (I39325), .I1 (g29713), .I2 (I39323));
ND2X1 gate21460(.O (g29911), .I1 (I39324), .I2 (I39325));
ND2X1 gate21461(.O (I39331), .I1 (g29705), .I2 (g29751));
ND2X1 gate21462(.O (I39332), .I1 (g29705), .I2 (I39331));
ND2X1 gate21463(.O (I39333), .I1 (g29751), .I2 (I39331));
ND2X1 gate21464(.O (g29913), .I1 (I39332), .I2 (I39333));
ND2X1 gate21465(.O (I39339), .I1 (g29748), .I2 (g29741));
ND2X1 gate21466(.O (I39340), .I1 (g29748), .I2 (I39339));
ND2X1 gate21467(.O (I39341), .I1 (g29741), .I2 (I39339));
ND2X1 gate21468(.O (g29915), .I1 (I39340), .I2 (I39341));
ND2X1 gate21469(.O (I39347), .I1 (g29732), .I2 (g29728));
ND2X1 gate21470(.O (I39348), .I1 (g29732), .I2 (I39347));
ND2X1 gate21471(.O (I39349), .I1 (g29728), .I2 (I39347));
ND2X1 gate21472(.O (g29917), .I1 (I39348), .I2 (I39349));
ND2X1 gate21473(.O (I39359), .I1 (g29766), .I2 (g15880));
ND2X1 gate21474(.O (I39360), .I1 (g29766), .I2 (I39359));
ND2X1 gate21475(.O (I39361), .I1 (g15880), .I2 (I39359));
ND2X1 gate21476(.O (g29923), .I1 (I39360), .I2 (I39361));
ND2X1 gate21477(.O (I39367), .I1 (g29767), .I2 (g15913));
ND2X1 gate21478(.O (I39368), .I1 (g29767), .I2 (I39367));
ND2X1 gate21479(.O (I39369), .I1 (g15913), .I2 (I39367));
ND2X1 gate21480(.O (g29925), .I1 (I39368), .I2 (I39369));
ND2X1 gate21481(.O (I39375), .I1 (g29768), .I2 (g15942));
ND2X1 gate21482(.O (I39376), .I1 (g29768), .I2 (I39375));
ND2X1 gate21483(.O (I39377), .I1 (g15942), .I2 (I39375));
ND2X1 gate21484(.O (g29927), .I1 (I39376), .I2 (I39377));
ND2X1 gate21485(.O (I39384), .I1 (g29718), .I2 (g29710));
ND2X1 gate21486(.O (I39385), .I1 (g29718), .I2 (I39384));
ND2X1 gate21487(.O (I39386), .I1 (g29710), .I2 (I39384));
ND2X1 gate21488(.O (g29930), .I1 (I39385), .I2 (I39386));
ND2X1 gate21489(.O (I39391), .I1 (g29769), .I2 (g15971));
ND2X1 gate21490(.O (I39392), .I1 (g29769), .I2 (I39391));
ND2X1 gate21491(.O (I39393), .I1 (g15971), .I2 (I39391));
ND2X1 gate21492(.O (g29931), .I1 (I39392), .I2 (I39393));
ND2X1 gate21493(.O (I39532), .I1 (g29915), .I2 (g29917));
ND2X1 gate21494(.O (I39533), .I1 (g29915), .I2 (I39532));
ND2X1 gate21495(.O (I39534), .I1 (g29917), .I2 (I39532));
ND2X1 gate21496(.O (g30034), .I1 (I39533), .I2 (I39534));
ND2X1 gate21497(.O (I39539), .I1 (g29911), .I2 (g29913));
ND2X1 gate21498(.O (I39540), .I1 (g29911), .I2 (I39539));
ND2X1 gate21499(.O (I39541), .I1 (g29913), .I2 (I39539));
ND2X1 gate21500(.O (g30035), .I1 (I39540), .I2 (I39541));
ND2X1 gate21501(.O (I39689), .I1 (g30035), .I2 (g30034));
ND2X1 gate21502(.O (I39690), .I1 (g30035), .I2 (I39689));
ND2X1 gate21503(.O (I39691), .I1 (g30034), .I2 (I39689));
ND2X1 gate21504(.O (g30228), .I1 (I39690), .I2 (I39691));
ND2X1 gate21505(.O (I40558), .I1 (g30605), .I2 (g30597));
ND2X1 gate21506(.O (I40559), .I1 (g30605), .I2 (I40558));
ND2X1 gate21507(.O (I40560), .I1 (g30597), .I2 (I40558));
ND2X1 gate21508(.O (g30768), .I1 (I40559), .I2 (I40560));
ND2X1 gate21509(.O (I40571), .I1 (g30588), .I2 (g30632));
ND2X1 gate21510(.O (I40572), .I1 (g30588), .I2 (I40571));
ND2X1 gate21511(.O (I40573), .I1 (g30632), .I2 (I40571));
ND2X1 gate21512(.O (g30771), .I1 (I40572), .I2 (I40573));
ND2X1 gate21513(.O (I40587), .I1 (g30629), .I2 (g30622));
ND2X1 gate21514(.O (I40588), .I1 (g30629), .I2 (I40587));
ND2X1 gate21515(.O (I40589), .I1 (g30622), .I2 (I40587));
ND2X1 gate21516(.O (g30775), .I1 (I40588), .I2 (I40589));
ND2X1 gate21517(.O (I40603), .I1 (g30614), .I2 (g30610));
ND2X1 gate21518(.O (I40604), .I1 (g30614), .I2 (I40603));
ND2X1 gate21519(.O (I40605), .I1 (g30610), .I2 (I40603));
ND2X1 gate21520(.O (g30779), .I1 (I40604), .I2 (I40605));
ND2X1 gate21521(.O (I40627), .I1 (g30602), .I2 (g30594));
ND2X1 gate21522(.O (I40628), .I1 (g30602), .I2 (I40627));
ND2X1 gate21523(.O (I40629), .I1 (g30594), .I2 (I40627));
ND2X1 gate21524(.O (g30791), .I1 (I40628), .I2 (I40629));
ND2X1 gate21525(.O (I41010), .I1 (g30775), .I2 (g30779));
ND2X1 gate21526(.O (I41011), .I1 (g30775), .I2 (I41010));
ND2X1 gate21527(.O (I41012), .I1 (g30779), .I2 (I41010));
ND2X1 gate21528(.O (g30926), .I1 (I41011), .I2 (I41012));
ND2X1 gate21529(.O (I41017), .I1 (g30768), .I2 (g30771));
ND2X1 gate21530(.O (I41018), .I1 (g30768), .I2 (I41017));
ND2X1 gate21531(.O (I41019), .I1 (g30771), .I2 (I41017));
ND2X1 gate21532(.O (g30927), .I1 (I41018), .I2 (I41019));
ND2X1 gate21533(.O (I41064), .I1 (g30927), .I2 (g30926));
ND2X1 gate21534(.O (I41065), .I1 (g30927), .I2 (I41064));
ND2X1 gate21535(.O (I41066), .I1 (g30926), .I2 (I41064));
ND2X1 gate21536(.O (g30952), .I1 (I41065), .I2 (I41066));
NR3X1 gate21537(.O (g7528), .I1 (g3151), .I2 (g3142), .I3 (g3147));
NR2X1 gate21538(.O (g7575), .I1 (g2984), .I2 (g2985));
NR2X1 gate21539(.O (g7795), .I1 (g2992), .I2 (g2991));
NR4X1 gate21540(.O (g8430), .I1 (g3198), .I2 (g8120), .I3 (g3194), .I4 (g3191));
NR3X1 gate21541(.O (g10784), .I1 (g5630), .I2 (g5649), .I3 (g5676));
NR3X1 gate21542(.O (g10789), .I1 (g5650), .I2 (g5677), .I3 (g5709));
NR3X1 gate21543(.O (g10793), .I1 (g5658), .I2 (g5687), .I3 (g5728));
NR3X1 gate21544(.O (g10797), .I1 (g5678), .I2 (g5710), .I3 (g5757));
NR3X1 gate21545(.O (g10801), .I1 (g5688), .I2 (g5729), .I3 (g5767));
NR3X1 gate21546(.O (g10805), .I1 (g5696), .I2 (g5739), .I3 (g5786));
NR3X1 gate21547(.O (g10810), .I1 (g5711), .I2 (g5758), .I3 (g5807));
NR3X1 gate21548(.O (g10814), .I1 (g5730), .I2 (g5768), .I3 (g5816));
NR3X1 gate21549(.O (g10818), .I1 (g5740), .I2 (g5787), .I3 (g5826));
NR3X1 gate21550(.O (g10822), .I1 (g5748), .I2 (g5797), .I3 (g5845));
NR3X1 gate21551(.O (g10831), .I1 (g5769), .I2 (g5817), .I3 (g5863));
NR3X1 gate21552(.O (g10835), .I1 (g5788), .I2 (g5827), .I3 (g5872));
NR3X1 gate21553(.O (g10839), .I1 (g5798), .I2 (g5846), .I3 (g5882));
NR3X1 gate21554(.O (g10851), .I1 (g5828), .I2 (g5873), .I3 (g5910));
NR3X1 gate21555(.O (g10855), .I1 (g5847), .I2 (g5883), .I3 (g5919));
NR3X1 gate21556(.O (g10872), .I1 (g5884), .I2 (g5920), .I3 (g5949));
NR3X1 gate21557(.O (g11600), .I1 (g9049), .I2 (g9064), .I3 (g9078));
NR4X1 gate21558(.O (g11622), .I1 (g8183), .I2 (g11332), .I3 (g7928), .I4 (g11069));
NR3X1 gate21559(.O (g11624), .I1 (g9062), .I2 (g9075), .I3 (g9091));
NR3X1 gate21560(.O (g11627), .I1 (g9063), .I2 (g9077), .I3 (g9093));
NR3X1 gate21561(.O (g11630), .I1 (g9066), .I2 (g9081), .I3 (g9097));
NR4X1 gate21562(.O (g11643), .I1 (g11481), .I2 (g8045), .I3 (g7928), .I4 (g11069));
NR3X1 gate21563(.O (g11644), .I1 (g9076), .I2 (g9092), .I3 (g9102));
NR3X1 gate21564(.O (g11647), .I1 (g9079), .I2 (g9094), .I3 (g9103));
NR3X1 gate21565(.O (g11650), .I1 (g9080), .I2 (g9096), .I3 (g9105));
NR3X1 gate21566(.O (g11653), .I1 (g9083), .I2 (g9100), .I3 (g9109));
NR4X1 gate21567(.O (g11660), .I1 (g8183), .I2 (g8045), .I3 (g7928), .I4 (g11069));
NR3X1 gate21568(.O (g11663), .I1 (g9095), .I2 (g9104), .I3 (g9112));
NR3X1 gate21569(.O (g11666), .I1 (g9098), .I2 (g9106), .I3 (g9113));
NR3X1 gate21570(.O (g11669), .I1 (g9099), .I2 (g9108), .I3 (g9115));
NR3X1 gate21571(.O (g11675), .I1 (g9107), .I2 (g9114), .I3 (g9120));
NR3X1 gate21572(.O (g11678), .I1 (g9110), .I2 (g9116), .I3 (g9121));
NR3X1 gate21573(.O (g11681), .I1 (g9111), .I2 (g9118), .I3 (g9123));
NR3X1 gate21574(.O (g11687), .I1 (g9117), .I2 (g9122), .I3 (g9126));
NR3X1 gate21575(.O (g11690), .I1 (g9119), .I2 (g9124), .I3 (g9127));
NR3X1 gate21576(.O (g11697), .I1 (g9125), .I2 (g9131), .I3 (g9133));
NR3X1 gate21577(.O (g11703), .I1 (g9132), .I2 (g9137), .I3 (g9139));
NR3X1 gate21578(.O (g11711), .I1 (g9138), .I2 (g9143), .I3 (g9145));
NR3X1 gate21579(.O (g11744), .I1 (g9241), .I2 (g9301), .I3 (g9364));
NR3X1 gate21580(.O (g11759), .I1 (g9302), .I2 (g9365), .I3 (g9438));
NR3X1 gate21581(.O (g11760), .I1 (g9319), .I2 (g9382), .I3 (g9461));
NR3X1 gate21582(.O (g11767), .I1 (g9366), .I2 (g9439), .I3 (g9518));
NR3X1 gate21583(.O (g11768), .I1 (g9367), .I2 (g9441), .I3 (g9521));
NR3X1 gate21584(.O (g11772), .I1 (g9383), .I2 (g9462), .I3 (g9580));
NR3X1 gate21585(.O (g11773), .I1 (g9400), .I2 (g9479), .I3 (g9603));
NR3X1 gate21586(.O (g11780), .I1 (g9440), .I2 (g9519), .I3 (g9630));
NR3X1 gate21587(.O (g11781), .I1 (g9442), .I2 (g9522), .I3 (g9633));
NR3X1 gate21588(.O (g11784), .I1 (g9463), .I2 (g9581), .I3 (g9660));
NR3X1 gate21589(.O (g11785), .I1 (g9464), .I2 (g9583), .I3 (g9663));
NR3X1 gate21590(.O (g11789), .I1 (g9480), .I2 (g9604), .I3 (g9722));
NR3X1 gate21591(.O (g11790), .I1 (g9497), .I2 (g9621), .I3 (g9745));
NR3X1 gate21592(.O (g11799), .I1 (g9520), .I2 (g9631), .I3 (g9759));
NR3X1 gate21593(.O (g11800), .I1 (g9523), .I2 (g9634), .I3 (g9762));
NR3X1 gate21594(.O (g11806), .I1 (g9582), .I2 (g9661), .I3 (g9776));
NR3X1 gate21595(.O (g11807), .I1 (g9584), .I2 (g9664), .I3 (g9779));
NR3X1 gate21596(.O (g11810), .I1 (g9605), .I2 (g9723), .I3 (g9806));
NR3X1 gate21597(.O (g11811), .I1 (g9606), .I2 (g9725), .I3 (g9809));
NR3X1 gate21598(.O (g11815), .I1 (g9622), .I2 (g9746), .I3 (g9868));
NR3X1 gate21599(.O (g11822), .I1 (g9632), .I2 (g9760), .I3 (g9888));
NR3X1 gate21600(.O (g11823), .I1 (g9635), .I2 (g9763), .I3 (g9891));
NR3X1 gate21601(.O (g11828), .I1 (g9639), .I2 (g9764), .I3 (g9892));
NR3X1 gate21602(.O (g11830), .I1 (g9647), .I2 (g9773), .I3 (g9901));
NR3X1 gate21603(.O (g11831), .I1 (g9648), .I2 (g9775), .I3 (g9904));
NR3X1 gate21604(.O (g11832), .I1 (g9662), .I2 (g9777), .I3 (g9905));
NR3X1 gate21605(.O (g11833), .I1 (g9665), .I2 (g9780), .I3 (g9908));
NR3X1 gate21606(.O (g11839), .I1 (g9724), .I2 (g9807), .I3 (g9922));
NR3X1 gate21607(.O (g11840), .I1 (g9726), .I2 (g9810), .I3 (g9925));
NR3X1 gate21608(.O (g11843), .I1 (g9747), .I2 (g9869), .I3 (g9952));
NR3X1 gate21609(.O (g11844), .I1 (g9748), .I2 (g9871), .I3 (g9955));
NR3X1 gate21610(.O (g11855), .I1 (g9761), .I2 (g9889), .I3 (g10009));
NR3X1 gate21611(.O (g11860), .I1 (g9765), .I2 (g9893), .I3 (g10012));
NR3X1 gate21612(.O (g11861), .I1 (g9766), .I2 (g9894), .I3 (g10013));
NR3X1 gate21613(.O (g11863), .I1 (g9774), .I2 (g9902), .I3 (g10035));
NR3X1 gate21614(.O (g11864), .I1 (g9778), .I2 (g9906), .I3 (g10042));
NR3X1 gate21615(.O (g11865), .I1 (g9781), .I2 (g9909), .I3 (g10045));
NR3X1 gate21616(.O (g11870), .I1 (g9785), .I2 (g9910), .I3 (g10046));
NR3X1 gate21617(.O (g11872), .I1 (g9793), .I2 (g9919), .I3 (g10055));
NR3X1 gate21618(.O (g11873), .I1 (g9794), .I2 (g9921), .I3 (g10058));
NR3X1 gate21619(.O (g11874), .I1 (g9808), .I2 (g9923), .I3 (g10059));
NR3X1 gate21620(.O (g11875), .I1 (g9811), .I2 (g9926), .I3 (g10062));
NR3X1 gate21621(.O (g11881), .I1 (g9870), .I2 (g9953), .I3 (g10076));
NR3X1 gate21622(.O (g11882), .I1 (g9872), .I2 (g9956), .I3 (g10079));
NR3X1 gate21623(.O (g11889), .I1 (g9887), .I2 (g10007), .I3 (g10101));
NR3X1 gate21624(.O (g11890), .I1 (g9890), .I2 (g10010), .I3 (g10103));
NR3X1 gate21625(.O (g11896), .I1 (g9903), .I2 (g10036), .I3 (g10112));
NR3X1 gate21626(.O (g11897), .I1 (g9907), .I2 (g10043), .I3 (g10118));
NR3X1 gate21627(.O (g11902), .I1 (g9911), .I2 (g10047), .I3 (g10121));
NR3X1 gate21628(.O (g11903), .I1 (g9912), .I2 (g10048), .I3 (g10122));
NR3X1 gate21629(.O (g11905), .I1 (g9920), .I2 (g10056), .I3 (g10144));
NR3X1 gate21630(.O (g11906), .I1 (g9924), .I2 (g10060), .I3 (g10151));
NR3X1 gate21631(.O (g11907), .I1 (g9927), .I2 (g10063), .I3 (g10154));
NR3X1 gate21632(.O (g11912), .I1 (g9931), .I2 (g10064), .I3 (g10155));
NR3X1 gate21633(.O (g11914), .I1 (g9939), .I2 (g10073), .I3 (g10164));
NR3X1 gate21634(.O (g11915), .I1 (g9940), .I2 (g10075), .I3 (g10167));
NR3X1 gate21635(.O (g11916), .I1 (g9954), .I2 (g10077), .I3 (g10168));
NR3X1 gate21636(.O (g11917), .I1 (g9957), .I2 (g10080), .I3 (g10171));
NR3X1 gate21637(.O (g11928), .I1 (g10008), .I2 (g10102), .I3 (g10192));
NR3X1 gate21638(.O (g11934), .I1 (g10011), .I2 (g10104), .I3 (g10193));
NR3X1 gate21639(.O (g11935), .I1 (g10014), .I2 (g10106), .I3 (g10196));
NR3X1 gate21640(.O (g11938), .I1 (g10037), .I2 (g10113), .I3 (g10201));
NR3X1 gate21641(.O (g11939), .I1 (g10041), .I2 (g10116), .I3 (g10206));
NR3X1 gate21642(.O (g11940), .I1 (g10044), .I2 (g10119), .I3 (g10208));
NR3X1 gate21643(.O (g11946), .I1 (g10057), .I2 (g10145), .I3 (g10217));
NR3X1 gate21644(.O (g11947), .I1 (g10061), .I2 (g10152), .I3 (g10223));
NR3X1 gate21645(.O (g11952), .I1 (g10065), .I2 (g10156), .I3 (g10226));
NR3X1 gate21646(.O (g11953), .I1 (g10066), .I2 (g10157), .I3 (g10227));
NR3X1 gate21647(.O (g11955), .I1 (g10074), .I2 (g10165), .I3 (g10249));
NR3X1 gate21648(.O (g11956), .I1 (g10078), .I2 (g10169), .I3 (g10256));
NR3X1 gate21649(.O (g11957), .I1 (g10081), .I2 (g10172), .I3 (g10259));
NR3X1 gate21650(.O (g11962), .I1 (g10085), .I2 (g10173), .I3 (g10260));
NR3X1 gate21651(.O (g11964), .I1 (g10093), .I2 (g10182), .I3 (g10269));
NR3X1 gate21652(.O (g11965), .I1 (g10094), .I2 (g10184), .I3 (g10272));
NR3X1 gate21653(.O (g11974), .I1 (g10105), .I2 (g10194), .I3 (g10279));
NR3X1 gate21654(.O (g11975), .I1 (g10107), .I2 (g10197), .I3 (g10282));
NR3X1 gate21655(.O (g11979), .I1 (g10114), .I2 (g10202), .I3 (g10288));
NR3X1 gate21656(.O (g11980), .I1 (g10115), .I2 (g10204), .I3 (g10291));
NR3X1 gate21657(.O (g11981), .I1 (g10117), .I2 (g10207), .I3 (g10294));
NR3X1 gate21658(.O (g11987), .I1 (g10120), .I2 (g10209), .I3 (g10295));
NR3X1 gate21659(.O (g11988), .I1 (g10123), .I2 (g10211), .I3 (g10298));
NR3X1 gate21660(.O (g11991), .I1 (g10146), .I2 (g10218), .I3 (g10303));
NR3X1 gate21661(.O (g11992), .I1 (g10150), .I2 (g10221), .I3 (g10308));
NR3X1 gate21662(.O (g11993), .I1 (g10153), .I2 (g10224), .I3 (g10310));
NR3X1 gate21663(.O (g11999), .I1 (g10166), .I2 (g10250), .I3 (g10319));
NR3X1 gate21664(.O (g12000), .I1 (g10170), .I2 (g10257), .I3 (g10325));
NR3X1 gate21665(.O (g12005), .I1 (g10174), .I2 (g10261), .I3 (g10328));
NR3X1 gate21666(.O (g12006), .I1 (g10175), .I2 (g10262), .I3 (g10329));
NR3X1 gate21667(.O (g12008), .I1 (g10183), .I2 (g10270), .I3 (g10351));
NR3X1 gate21668(.O (g12026), .I1 (g10195), .I2 (g10280), .I3 (g10360));
NR3X1 gate21669(.O (g12033), .I1 (g10199), .I2 (g10284), .I3 (g10362));
NR3X1 gate21670(.O (g12034), .I1 (g10200), .I2 (g10286), .I3 (g10365));
NR3X1 gate21671(.O (g12035), .I1 (g10203), .I2 (g10289), .I3 (g10367));
NR3X1 gate21672(.O (g12036), .I1 (g10205), .I2 (g10292), .I3 (g10370));
NR3X1 gate21673(.O (g12043), .I1 (g10210), .I2 (g10296), .I3 (g10372));
NR3X1 gate21674(.O (g12044), .I1 (g10212), .I2 (g10299), .I3 (g10375));
NR3X1 gate21675(.O (g12048), .I1 (g10219), .I2 (g10304), .I3 (g10381));
NR3X1 gate21676(.O (g12049), .I1 (g10220), .I2 (g10306), .I3 (g10384));
NR3X1 gate21677(.O (g12050), .I1 (g10222), .I2 (g10309), .I3 (g10387));
NR3X1 gate21678(.O (g12056), .I1 (g10225), .I2 (g10311), .I3 (g10388));
NR3X1 gate21679(.O (g12057), .I1 (g10228), .I2 (g10313), .I3 (g10391));
NR3X1 gate21680(.O (g12060), .I1 (g10251), .I2 (g10320), .I3 (g10396));
NR3X1 gate21681(.O (g12061), .I1 (g10255), .I2 (g10323), .I3 (g10401));
NR3X1 gate21682(.O (g12062), .I1 (g10258), .I2 (g10326), .I3 (g10403));
NR3X1 gate21683(.O (g12068), .I1 (g10271), .I2 (g10352), .I3 (g10412));
NR3X1 gate21684(.O (g12079), .I1 (g10281), .I2 (g10361), .I3 (g10422));
NR3X1 gate21685(.O (g12080), .I1 (g10285), .I2 (g10363), .I3 (g10430));
NR3X1 gate21686(.O (g12081), .I1 (g10287), .I2 (g10366), .I3 (g10433));
NR3X1 gate21687(.O (g12082), .I1 (g10290), .I2 (g10368), .I3 (g10435));
NR3X1 gate21688(.O (g12083), .I1 (g10293), .I2 (g10371), .I3 (g10438));
NR3X1 gate21689(.O (g12090), .I1 (g10297), .I2 (g10373), .I3 (g10439));
NR3X1 gate21690(.O (g12097), .I1 (g10301), .I2 (g10377), .I3 (g10441));
NR3X1 gate21691(.O (g12098), .I1 (g10302), .I2 (g10379), .I3 (g10444));
NR3X1 gate21692(.O (g12099), .I1 (g10305), .I2 (g10382), .I3 (g10446));
NR3X1 gate21693(.O (g12100), .I1 (g10307), .I2 (g10385), .I3 (g10449));
NR3X1 gate21694(.O (g12107), .I1 (g10312), .I2 (g10389), .I3 (g10451));
NR3X1 gate21695(.O (g12108), .I1 (g10314), .I2 (g10392), .I3 (g10454));
NR3X1 gate21696(.O (g12112), .I1 (g10321), .I2 (g10397), .I3 (g10460));
NR3X1 gate21697(.O (g12113), .I1 (g10322), .I2 (g10399), .I3 (g10463));
NR3X1 gate21698(.O (g12114), .I1 (g10324), .I2 (g10402), .I3 (g10466));
NR3X1 gate21699(.O (g12120), .I1 (g10327), .I2 (g10404), .I3 (g10467));
NR3X1 gate21700(.O (g12121), .I1 (g10330), .I2 (g10406), .I3 (g10470));
NR3X1 gate21701(.O (g12124), .I1 (g10353), .I2 (g10413), .I3 (g10475));
NR3X1 gate21702(.O (g12145), .I1 (g10364), .I2 (g10431), .I3 (g10492));
NR3X1 gate21703(.O (g12146), .I1 (g10369), .I2 (g10436), .I3 (g10496));
NR3X1 gate21704(.O (g12151), .I1 (g10374), .I2 (g10440), .I3 (g10498));
NR3X1 gate21705(.O (g12152), .I1 (g10378), .I2 (g10442), .I3 (g10506));
NR3X1 gate21706(.O (g12153), .I1 (g10380), .I2 (g10445), .I3 (g10509));
NR3X1 gate21707(.O (g12154), .I1 (g10383), .I2 (g10447), .I3 (g10511));
NR3X1 gate21708(.O (g12155), .I1 (g10386), .I2 (g10450), .I3 (g10514));
NR3X1 gate21709(.O (g12162), .I1 (g10390), .I2 (g10452), .I3 (g10515));
NR3X1 gate21710(.O (g12169), .I1 (g10394), .I2 (g10456), .I3 (g10517));
NR3X1 gate21711(.O (g12170), .I1 (g10395), .I2 (g10458), .I3 (g10520));
NR3X1 gate21712(.O (g12171), .I1 (g10398), .I2 (g10461), .I3 (g10522));
NR3X1 gate21713(.O (g12172), .I1 (g10400), .I2 (g10464), .I3 (g10525));
NR3X1 gate21714(.O (g12179), .I1 (g10405), .I2 (g10468), .I3 (g10527));
NR3X1 gate21715(.O (g12180), .I1 (g10407), .I2 (g10471), .I3 (g10530));
NR3X1 gate21716(.O (g12184), .I1 (g10414), .I2 (g10476), .I3 (g10536));
NR3X1 gate21717(.O (g12185), .I1 (g10415), .I2 (g10478), .I3 (g10539));
NR3X1 gate21718(.O (g12192), .I1 (g10423), .I2 (g10485), .I3 (g10548));
NR3X1 gate21719(.O (g12193), .I1 (g10432), .I2 (g10493), .I3 (g10555));
NR3X1 gate21720(.O (g12194), .I1 (g10434), .I2 (g10494), .I3 (g10556));
NR3X1 gate21721(.O (g12195), .I1 (g10437), .I2 (g10497), .I3 (g10558));
NR3X1 gate21722(.O (g12207), .I1 (g10443), .I2 (g10507), .I3 (g10566));
NR3X1 gate21723(.O (g12208), .I1 (g10448), .I2 (g10512), .I3 (g10570));
NR3X1 gate21724(.O (g12213), .I1 (g10453), .I2 (g10516), .I3 (g10572));
NR3X1 gate21725(.O (g12214), .I1 (g10457), .I2 (g10518), .I3 (g10580));
NR3X1 gate21726(.O (g12215), .I1 (g10459), .I2 (g10521), .I3 (g10583));
NR3X1 gate21727(.O (g12216), .I1 (g10462), .I2 (g10523), .I3 (g10585));
NR3X1 gate21728(.O (g12217), .I1 (g10465), .I2 (g10526), .I3 (g10588));
NR3X1 gate21729(.O (g12224), .I1 (g10469), .I2 (g10528), .I3 (g10589));
NR3X1 gate21730(.O (g12231), .I1 (g10473), .I2 (g10532), .I3 (g10591));
NR3X1 gate21731(.O (g12232), .I1 (g10474), .I2 (g10534), .I3 (g10594));
NR3X1 gate21732(.O (g12233), .I1 (g10477), .I2 (g10537), .I3 (g10596));
NR3X1 gate21733(.O (g12234), .I1 (g10479), .I2 (g10540), .I3 (g10599));
NR3X1 gate21734(.O (g12245), .I1 (g10495), .I2 (g10557), .I3 (g10604));
NR3X1 gate21735(.O (g12247), .I1 (g10499), .I2 (g10559), .I3 (g10605));
NR3X1 gate21736(.O (g12248), .I1 (g10508), .I2 (g10567), .I3 (g10612));
NR3X1 gate21737(.O (g12249), .I1 (g10510), .I2 (g10568), .I3 (g10613));
NR3X1 gate21738(.O (g12250), .I1 (g10513), .I2 (g10571), .I3 (g10615));
NR3X1 gate21739(.O (g12262), .I1 (g10519), .I2 (g10581), .I3 (g10623));
NR3X1 gate21740(.O (g12263), .I1 (g10524), .I2 (g10586), .I3 (g10627));
NR3X1 gate21741(.O (g12268), .I1 (g10529), .I2 (g10590), .I3 (g10629));
NR3X1 gate21742(.O (g12269), .I1 (g10533), .I2 (g10592), .I3 (g10637));
NR3X1 gate21743(.O (g12270), .I1 (g10535), .I2 (g10595), .I3 (g10640));
NR3X1 gate21744(.O (g12271), .I1 (g10538), .I2 (g10597), .I3 (g10642));
NR3X1 gate21745(.O (g12272), .I1 (g10541), .I2 (g10600), .I3 (g10645));
NR3X1 gate21746(.O (g12288), .I1 (g10569), .I2 (g10614), .I3 (g10651));
NR3X1 gate21747(.O (g12290), .I1 (g10573), .I2 (g10616), .I3 (g10652));
NR3X1 gate21748(.O (g12291), .I1 (g10582), .I2 (g10624), .I3 (g10659));
NR3X1 gate21749(.O (g12292), .I1 (g10584), .I2 (g10625), .I3 (g10660));
NR3X1 gate21750(.O (g12293), .I1 (g10587), .I2 (g10628), .I3 (g10662));
NR3X1 gate21751(.O (g12305), .I1 (g10593), .I2 (g10638), .I3 (g10670));
NR3X1 gate21752(.O (g12306), .I1 (g10598), .I2 (g10643), .I3 (g10674));
NR3X1 gate21753(.O (g12324), .I1 (g10626), .I2 (g10661), .I3 (g10681));
NR3X1 gate21754(.O (g12326), .I1 (g10630), .I2 (g10663), .I3 (g10682));
NR3X1 gate21755(.O (g12327), .I1 (g10639), .I2 (g10671), .I3 (g10689));
NR3X1 gate21756(.O (g12328), .I1 (g10641), .I2 (g10672), .I3 (g10690));
NR3X1 gate21757(.O (g12329), .I1 (g10644), .I2 (g10675), .I3 (g10692));
NR3X1 gate21758(.O (g12339), .I1 (g10650), .I2 (g10678), .I3 (g10704));
NR3X1 gate21759(.O (g12352), .I1 (g10673), .I2 (g10691), .I3 (g10710));
NR3X1 gate21760(.O (g12369), .I1 (g10680), .I2 (g10707), .I3 (g10724));
NR3X1 gate21761(.O (g12388), .I1 (g10709), .I2 (g10727), .I3 (g10745));
NR3X1 gate21762(.O (g12418), .I1 (g10729), .I2 (g10748), .I3 (g10764));
NR2X1 gate21763(.O (g12431), .I1 (g8580), .I2 (g10730));
NR2X1 gate21764(.O (g12436), .I1 (g8587), .I2 (g10749));
NR2X1 gate21765(.O (g12441), .I1 (g8594), .I2 (g10767));
NR2X1 gate21766(.O (g12446), .I1 (g8605), .I2 (g10773));
NR2X1 gate21767(.O (g12451), .I1 (g499), .I2 (g8983));
NR3X1 gate21768(.O (g12457), .I1 (g9009), .I2 (g9033), .I3 (g9048));
NR3X1 gate21769(.O (g12467), .I1 (g9034), .I2 (g9056), .I3 (g9065));
NR3X1 gate21770(.O (g12482), .I1 (g9057), .I2 (g9073), .I3 (g9082));
NR3X1 gate21771(.O (g12487), .I1 (g10108), .I2 (g10198), .I3 (g10283));
NR3X1 gate21772(.O (g12499), .I1 (g9074), .I2 (g9090), .I3 (g9101));
NR3X1 gate21773(.O (g12507), .I1 (g10213), .I2 (g10300), .I3 (g10376));
NR3X1 gate21774(.O (g12524), .I1 (g10315), .I2 (g10393), .I3 (g10455));
NR3X1 gate21775(.O (g12539), .I1 (g10408), .I2 (g10472), .I3 (g10531));
NR3X1 gate21776(.O (g12698), .I1 (g11347), .I2 (g11420), .I3 (g8327));
NR3X1 gate21777(.O (g12747), .I1 (g11421), .I2 (g8328), .I3 (g8385));
NR3X1 gate21778(.O (g12755), .I1 (g11431), .I2 (g8339), .I3 (g8394));
NR2X1 gate21779(.O (g12780), .I1 (g9187), .I2 (g9161));
NR3X1 gate21780(.O (g12781), .I1 (g8329), .I2 (g8386), .I3 (g8431));
NR3X1 gate21781(.O (g12789), .I1 (g8340), .I2 (g8395), .I3 (g8437));
NR3X1 gate21782(.O (g12797), .I1 (g8350), .I2 (g8406), .I3 (g8446));
NR3X1 gate21783(.O (g12814), .I1 (g8387), .I2 (g8432), .I3 (g8463));
NR2X1 gate21784(.O (g12819), .I1 (g9248), .I2 (g9203));
NR3X1 gate21785(.O (g12820), .I1 (g8396), .I2 (g8438), .I3 (g8466));
NR3X1 gate21786(.O (g12828), .I1 (g8407), .I2 (g8447), .I3 (g8472));
NR3X1 gate21787(.O (g12836), .I1 (g8417), .I2 (g8458), .I3 (g8481));
NR3X1 gate21788(.O (g12849), .I1 (g8433), .I2 (g8464), .I3 (g8485));
NR3X1 gate21789(.O (g12852), .I1 (g8439), .I2 (g8467), .I3 (g8488));
NR2X1 gate21790(.O (g12857), .I1 (g9326), .I2 (g9264));
NR3X1 gate21791(.O (g12858), .I1 (g8448), .I2 (g8473), .I3 (g8491));
NR3X1 gate21792(.O (g12866), .I1 (g8459), .I2 (g8482), .I3 (g8497));
NR3X1 gate21793(.O (g12880), .I1 (g8465), .I2 (g8486), .I3 (g8502));
NR2X1 gate21794(.O (g12883), .I1 (g10038), .I2 (g6284));
NR3X1 gate21795(.O (g12890), .I1 (g8468), .I2 (g8489), .I3 (g8505));
NR3X1 gate21796(.O (g12893), .I1 (g8474), .I2 (g8492), .I3 (g8508));
NR2X1 gate21797(.O (g12898), .I1 (g9407), .I2 (g9342));
NR3X1 gate21798(.O (g12899), .I1 (g8483), .I2 (g8498), .I3 (g8511));
NR3X1 gate21799(.O (g12912), .I1 (g8484), .I2 (g8500), .I3 (g8515));
NR3X1 gate21800(.O (g12913), .I1 (g8487), .I2 (g8503), .I3 (g8518));
NR3X1 gate21801(.O (g12920), .I1 (g8490), .I2 (g8506), .I3 (g8521));
NR2X1 gate21802(.O (g12923), .I1 (g10147), .I2 (g6421));
NR3X1 gate21803(.O (g12930), .I1 (g8493), .I2 (g8509), .I3 (g8524));
NR3X1 gate21804(.O (g12933), .I1 (g8499), .I2 (g8512), .I3 (g8527));
NR3X1 gate21805(.O (g12939), .I1 (g8501), .I2 (g8516), .I3 (g8531));
NR3X1 gate21806(.O (g12941), .I1 (g8504), .I2 (g8519), .I3 (g8534));
NR3X1 gate21807(.O (g12942), .I1 (g8507), .I2 (g8522), .I3 (g8537));
NR3X1 gate21808(.O (g12949), .I1 (g8510), .I2 (g8525), .I3 (g8540));
NR2X1 gate21809(.O (g12952), .I1 (g10252), .I2 (g6626));
NR3X1 gate21810(.O (g12959), .I1 (g8513), .I2 (g8528), .I3 (g8543));
NR3X1 gate21811(.O (g12967), .I1 (g8517), .I2 (g8532), .I3 (g8546));
NR3X1 gate21812(.O (g12968), .I1 (g8520), .I2 (g8535), .I3 (g8548));
NR3X1 gate21813(.O (g12970), .I1 (g8523), .I2 (g8538), .I3 (g8551));
NR3X1 gate21814(.O (g12971), .I1 (g8526), .I2 (g8541), .I3 (g8554));
NR3X1 gate21815(.O (g12978), .I1 (g8529), .I2 (g8544), .I3 (g8557));
NR2X1 gate21816(.O (g12981), .I1 (g10354), .I2 (g6890));
NR3X1 gate21817(.O (g12991), .I1 (g8536), .I2 (g8549), .I3 (g8559));
NR3X1 gate21818(.O (g12992), .I1 (g8539), .I2 (g8552), .I3 (g8561));
NR3X1 gate21819(.O (g12994), .I1 (g8542), .I2 (g8555), .I3 (g8564));
NR3X1 gate21820(.O (g12995), .I1 (g8545), .I2 (g8558), .I3 (g8567));
NR3X1 gate21821(.O (g13001), .I1 (g8553), .I2 (g8562), .I3 (g8570));
NR3X1 gate21822(.O (g13002), .I1 (g8556), .I2 (g8565), .I3 (g8572));
NR3X1 gate21823(.O (g13022), .I1 (g8566), .I2 (g8573), .I3 (g8576));
NR4X1 gate21824(.O (g13024), .I1 (g11481), .I2 (g8045), .I3 (g7928), .I4 (g7880));
NR3X1 gate21825(.O (g13111), .I1 (g8601), .I2 (g8612), .I3 (g8621));
NR3X1 gate21826(.O (g13124), .I1 (g8613), .I2 (g8625), .I3 (g8631));
NR3X1 gate21827(.O (g13135), .I1 (g8626), .I2 (g8635), .I3 (g8650));
NR3X1 gate21828(.O (g13143), .I1 (g8636), .I2 (g8654), .I3 (g8666));
NR3X1 gate21829(.O (g13149), .I1 (g8676), .I2 (g8687), .I3 (g8703));
NR3X1 gate21830(.O (g13155), .I1 (g8688), .I2 (g8705), .I3 (g8722));
NR3X1 gate21831(.O (g13160), .I1 (g8704), .I2 (g8717), .I3 (g8751));
NR3X1 gate21832(.O (g13164), .I1 (g8706), .I2 (g8724), .I3 (g8760));
NR3X1 gate21833(.O (g13171), .I1 (g8723), .I2 (g8755), .I3 (g8774));
NR3X1 gate21834(.O (g13175), .I1 (g8725), .I2 (g8762), .I3 (g8783));
NR3X1 gate21835(.O (g13182), .I1 (g8761), .I2 (g8778), .I3 (g8797));
NR3X1 gate21836(.O (g13194), .I1 (g8784), .I2 (g8801), .I3 (g8816));
NR3X1 gate21837(.O (g13228), .I1 (g8841), .I2 (g8861), .I3 (g8892));
NR3X1 gate21838(.O (g13251), .I1 (g8868), .I2 (g8899), .I3 (g8932));
NR3X1 gate21839(.O (g13274), .I1 (g8906), .I2 (g8939), .I3 (g8972));
NR4X1 gate21840(.O (g13286), .I1 (g11481), .I2 (g11332), .I3 (g11190), .I4 (g7880));
NR3X1 gate21841(.O (g13299), .I1 (g8946), .I2 (g8979), .I3 (g9004));
NR4X1 gate21842(.O (g13310), .I1 (g11481), .I2 (g11332), .I3 (g11190), .I4 (g11069));
NR4X1 gate21843(.O (g13313), .I1 (g8183), .I2 (g11332), .I3 (g11190), .I4 (g7880));
NR4X1 gate21844(.O (g13331), .I1 (g8183), .I2 (g11332), .I3 (g11190), .I4 (g11069));
NR4X1 gate21845(.O (g13332), .I1 (g11481), .I2 (g8045), .I3 (g11190), .I4 (g7880));
NR4X1 gate21846(.O (g13353), .I1 (g11481), .I2 (g8045), .I3 (g11190), .I4 (g11069));
NR4X1 gate21847(.O (g13354), .I1 (g8183), .I2 (g8045), .I3 (g11190), .I4 (g7880));
NR4X1 gate21848(.O (g13374), .I1 (g8183), .I2 (g8045), .I3 (g11190), .I4 (g11069));
NR4X1 gate21849(.O (g13375), .I1 (g11481), .I2 (g11332), .I3 (g7928), .I4 (g7880));
NR3X1 gate21850(.O (g13378), .I1 (g9026), .I2 (g9047), .I3 (g9061));
NR4X1 gate21851(.O (g13401), .I1 (g11481), .I2 (g11332), .I3 (g7928), .I4 (g11069));
NR4X1 gate21852(.O (g13404), .I1 (g8183), .I2 (g11332), .I3 (g7928), .I4 (g7880));
NR2X1 gate21853(.O (g15661), .I1 (g11737), .I2 (g7345));
NR2X1 gate21854(.O (g15797), .I1 (g13305), .I2 (g7143));
NR2X1 gate21855(.O (g15873), .I1 (g11617), .I2 (g7562));
NR2X1 gate21856(.O (g15959), .I1 (g2814), .I2 (g13082));
NR2X1 gate21857(.O (g15978), .I1 (g11737), .I2 (g7152));
NR3X1 gate21858(.O (g16020), .I1 (g6200), .I2 (g12457), .I3 (g10952));
NR3X1 gate21859(.O (g16036), .I1 (g6289), .I2 (g12467), .I3 (g10952));
NR3X1 gate21860(.O (g16058), .I1 (g6426), .I2 (g12482), .I3 (g10952));
NR3X1 gate21861(.O (g16082), .I1 (g10952), .I2 (g6140), .I3 (g12487));
NR3X1 gate21862(.O (g16094), .I1 (g6631), .I2 (g12499), .I3 (g10952));
NR3X1 gate21863(.O (g16120), .I1 (g10952), .I2 (g6161), .I3 (g12507));
NR3X1 gate21864(.O (g16171), .I1 (g10952), .I2 (g6188), .I3 (g12524));
NR3X1 gate21865(.O (g16230), .I1 (g10952), .I2 (g6220), .I3 (g12539));
NR2X1 gate21866(.O (g16498), .I1 (g14158), .I2 (g14347));
NR2X1 gate21867(.O (g16520), .I1 (g14273), .I2 (g14459));
NR2X1 gate21868(.O (g16551), .I1 (g14395), .I2 (g14546));
NR3X1 gate21869(.O (g16567), .I1 (g15904), .I2 (g15880), .I3 (g15859));
NR3X1 gate21870(.O (g16570), .I1 (g15904), .I2 (g15880), .I3 (g14630));
NR2X1 gate21871(.O (g16583), .I1 (g14507), .I2 (g14601));
NR3X1 gate21872(.O (g16591), .I1 (g15933), .I2 (g15913), .I3 (g15890));
NR3X1 gate21873(.O (g16594), .I1 (g15933), .I2 (g15913), .I3 (g14650));
NR3X1 gate21874(.O (g16611), .I1 (g15962), .I2 (g15942), .I3 (g15923));
NR3X1 gate21875(.O (g16614), .I1 (g15962), .I2 (g15942), .I3 (g14677));
NR3X1 gate21876(.O (g16629), .I1 (g15981), .I2 (g15971), .I3 (g15952));
NR3X1 gate21877(.O (g16632), .I1 (g15981), .I2 (g15971), .I3 (g14711));
NR3X1 gate21878(.O (g16643), .I1 (g15904), .I2 (g14642), .I3 (g15859));
NR2X1 gate21879(.O (g16654), .I1 (g14690), .I2 (g12477));
NR3X1 gate21880(.O (g16655), .I1 (g15933), .I2 (g14669), .I3 (g15890));
NR2X1 gate21881(.O (g16671), .I1 (g14724), .I2 (g12494));
NR3X1 gate21882(.O (g16672), .I1 (g15962), .I2 (g14703), .I3 (g15923));
NR2X1 gate21883(.O (g16679), .I1 (g14797), .I2 (g14895));
NR2X1 gate21884(.O (g16692), .I1 (g14752), .I2 (g12514));
NR3X1 gate21885(.O (g16693), .I1 (g15981), .I2 (g14737), .I3 (g15952));
NR2X1 gate21886(.O (g16705), .I1 (g14849), .I2 (g14976));
NR2X1 gate21887(.O (g16718), .I1 (g14773), .I2 (g12531));
NR2X1 gate21888(.O (g16736), .I1 (g14922), .I2 (g15065));
NR2X1 gate21889(.O (g16778), .I1 (g15003), .I2 (g15161));
NR2X1 gate21890(.O (g16802), .I1 (g13469), .I2 (g3897));
NR2X1 gate21891(.O (g16803), .I1 (g15593), .I2 (g12908));
NR2X1 gate21892(.O (g16823), .I1 (g5362), .I2 (g13469));
NR2X1 gate21893(.O (g16824), .I1 (g15658), .I2 (g12938));
NR2X1 gate21894(.O (g16829), .I1 (g14956), .I2 (g12564));
NR2X1 gate21895(.O (g16835), .I1 (g15717), .I2 (g12966));
NR2X1 gate21896(.O (g16841), .I1 (g15021), .I2 (g12607));
NR2X1 gate21897(.O (g16844), .I1 (g15754), .I2 (g12989));
NR2X1 gate21898(.O (g16845), .I1 (g15755), .I2 (g12990));
NR2X1 gate21899(.O (g16847), .I1 (g15095), .I2 (g12650));
NR2X1 gate21900(.O (g16851), .I1 (g15781), .I2 (g13000));
NR2X1 gate21901(.O (g16853), .I1 (g15801), .I2 (g13009));
NR2X1 gate21902(.O (g16854), .I1 (g15802), .I2 (g13010));
NR2X1 gate21903(.O (g16857), .I1 (g15817), .I2 (g13023));
NR2X1 gate21904(.O (g16860), .I1 (g15828), .I2 (g13031));
NR2X1 gate21905(.O (g16861), .I1 (g15829), .I2 (g13032));
NR2X1 gate21906(.O (g16866), .I1 (g15840), .I2 (g13042));
NR2X1 gate21907(.O (g16880), .I1 (g15852), .I2 (g13056));
NR3X1 gate21908(.O (g17012), .I1 (g14657), .I2 (g14642), .I3 (g15859));
NR3X1 gate21909(.O (g17025), .I1 (g15904), .I2 (g15880), .I3 (g15859));
NR3X1 gate21910(.O (g17042), .I1 (g14691), .I2 (g14669), .I3 (g15890));
NR3X1 gate21911(.O (g17051), .I1 (g14657), .I2 (g15880), .I3 (g14630));
NR3X1 gate21912(.O (g17059), .I1 (g15933), .I2 (g15913), .I3 (g15890));
NR3X1 gate21913(.O (g17076), .I1 (g14725), .I2 (g14703), .I3 (g15923));
NR3X1 gate21914(.O (g17086), .I1 (g14691), .I2 (g15913), .I3 (g14650));
NR3X1 gate21915(.O (g17094), .I1 (g15962), .I2 (g15942), .I3 (g15923));
NR3X1 gate21916(.O (g17111), .I1 (g14753), .I2 (g14737), .I3 (g15952));
NR3X1 gate21917(.O (g17124), .I1 (g14725), .I2 (g15942), .I3 (g14677));
NR3X1 gate21918(.O (g17132), .I1 (g15981), .I2 (g15971), .I3 (g15952));
NR3X1 gate21919(.O (g17151), .I1 (g14753), .I2 (g15971), .I3 (g14711));
NR2X1 gate21920(.O (g17186), .I1 (g7949), .I2 (g14144));
NR2X1 gate21921(.O (g17197), .I1 (g8000), .I2 (g14259));
NR2X1 gate21922(.O (g17204), .I1 (g8075), .I2 (g14381));
NR2X1 gate21923(.O (g17209), .I1 (g8160), .I2 (g14493));
NR2X1 gate21924(.O (g17213), .I1 (g4326), .I2 (g14442));
NR2X1 gate21925(.O (g17215), .I1 (g15904), .I2 (g14642));
NR2X1 gate21926(.O (g17216), .I1 (g4495), .I2 (g14529));
NR2X1 gate21927(.O (g17218), .I1 (g15933), .I2 (g14669));
NR2X1 gate21928(.O (g17219), .I1 (g4671), .I2 (g14584));
NR2X1 gate21929(.O (g17220), .I1 (g15962), .I2 (g14703));
NR2X1 gate21930(.O (g17221), .I1 (g4848), .I2 (g14618));
NR2X1 gate21931(.O (g17222), .I1 (g15998), .I2 (g16003));
NR2X1 gate21932(.O (g17223), .I1 (g15981), .I2 (g14737));
NR2X1 gate21933(.O (g17224), .I1 (g16004), .I2 (g16009));
NR2X1 gate21934(.O (g17225), .I1 (g16008), .I2 (g16015));
NR2X1 gate21935(.O (g17226), .I1 (g16010), .I2 (g16017));
NR2X1 gate21936(.O (g17228), .I1 (g16016), .I2 (g16029));
NR2X1 gate21937(.O (g17229), .I1 (g16019), .I2 (g16032));
NR2X1 gate21938(.O (g17234), .I1 (g16028), .I2 (g16045));
NR2X1 gate21939(.O (g17235), .I1 (g16030), .I2 (g16047));
NR2X1 gate21940(.O (g17236), .I1 (g16033), .I2 (g16051));
NR2X1 gate21941(.O (g17246), .I1 (g16046), .I2 (g16066));
NR2X1 gate21942(.O (g17247), .I1 (g16050), .I2 (g16070));
NR2X1 gate21943(.O (g17248), .I1 (g16052), .I2 (g16072));
NR2X1 gate21944(.O (g17269), .I1 (g16067), .I2 (g16100));
NR2X1 gate21945(.O (g17270), .I1 (g16071), .I2 (g16104));
NR2X1 gate21946(.O (g17271), .I1 (g16073), .I2 (g16106));
NR2X1 gate21947(.O (g17302), .I1 (g16103), .I2 (g16135));
NR2X1 gate21948(.O (g17303), .I1 (g16105), .I2 (g16137));
NR2X1 gate21949(.O (g17340), .I1 (g16136), .I2 (g16183));
NR2X1 gate21950(.O (g17341), .I1 (g16138), .I2 (g16185));
NR2X1 gate21951(.O (g17383), .I1 (g16184), .I2 (g16238));
NR2X1 gate21952(.O (g17429), .I1 (g16239), .I2 (g16288));
NR2X1 gate21953(.O (g17507), .I1 (g16298), .I2 (g13318));
NR2X1 gate21954(.O (g17896), .I1 (g14352), .I2 (g16020));
NR2X1 gate21955(.O (g18007), .I1 (g14464), .I2 (g16036));
NR2X1 gate21956(.O (g18085), .I1 (g16085), .I2 (g6363));
NR2X1 gate21957(.O (g18124), .I1 (g14551), .I2 (g16058));
NR2X1 gate21958(.O (g18201), .I1 (g16123), .I2 (g6568));
NR2X1 gate21959(.O (g18240), .I1 (g14606), .I2 (g16094));
NR2X1 gate21960(.O (g18308), .I1 (g16174), .I2 (g6832));
NR2X1 gate21961(.O (g18352), .I1 (g16082), .I2 (g14249));
NR2X1 gate21962(.O (g18401), .I1 (g16233), .I2 (g7134));
NR2X1 gate21963(.O (g18430), .I1 (g16020), .I2 (g14352));
NR2X1 gate21964(.O (g18447), .I1 (g16120), .I2 (g14371));
NR2X1 gate21965(.O (g18503), .I1 (g16036), .I2 (g14464));
NR2X1 gate21966(.O (g18520), .I1 (g16171), .I2 (g14483));
NR2X1 gate21967(.O (g18548), .I1 (g14249), .I2 (g16082));
NR2X1 gate21968(.O (g18567), .I1 (g16058), .I2 (g14551));
NR2X1 gate21969(.O (g18584), .I1 (g16230), .I2 (g14570));
NR2X1 gate21970(.O (g18590), .I1 (g16439), .I2 (g7522));
NR2X1 gate21971(.O (g18598), .I1 (g14371), .I2 (g16120));
NR2X1 gate21972(.O (g18617), .I1 (g16094), .I2 (g14606));
NR2X1 gate21973(.O (g18623), .I1 (g15902), .I2 (g2814));
NR2X1 gate21974(.O (g18626), .I1 (g16463), .I2 (g7549));
NR2X1 gate21975(.O (g18630), .I1 (g14483), .I2 (g16171));
NR2X1 gate21976(.O (g18639), .I1 (g14570), .I2 (g16230));
NR2X1 gate21977(.O (g18669), .I1 (g13623), .I2 (g13634));
NR2X1 gate21978(.O (g18678), .I1 (g13625), .I2 (g11771));
NR2X1 gate21979(.O (g18707), .I1 (g13636), .I2 (g11788));
NR2X1 gate21980(.O (g18719), .I1 (g13643), .I2 (g13656));
NR2X1 gate21981(.O (g18726), .I1 (g13645), .I2 (g11805));
NR2X1 gate21982(.O (g18743), .I1 (g13648), .I2 (g11814));
NR2X1 gate21983(.O (g18754), .I1 (g13655), .I2 (g11816));
NR2X1 gate21984(.O (g18755), .I1 (g13871), .I2 (g12274));
NR2X1 gate21985(.O (g18763), .I1 (g13671), .I2 (g11838));
NR2X1 gate21986(.O (g18780), .I1 (g13674), .I2 (g11847));
NR2X1 gate21987(.O (g18781), .I1 (g13675), .I2 (g11851));
NR2X1 gate21988(.O (g18782), .I1 (g13676), .I2 (g13705));
NR2X1 gate21989(.O (g18794), .I1 (g13701), .I2 (g11880));
NR2X1 gate21990(.O (g18803), .I1 (g13704), .I2 (g11885));
NR2X1 gate21991(.O (g18804), .I1 (g13905), .I2 (g12331));
NR2X1 gate21992(.O (g18820), .I1 (g13738), .I2 (g11922));
NR2X1 gate21993(.O (g18821), .I1 (g13740), .I2 (g11926));
NR2X1 gate21994(.O (g18835), .I1 (g13788), .I2 (g11966));
NR2X1 gate21995(.O (g18836), .I1 (g13789), .I2 (g11967));
NR2X1 gate21996(.O (g18837), .I1 (g13998), .I2 (g12376));
NR2X1 gate21997(.O (g18852), .I1 (g13815), .I2 (g12012));
NR2X1 gate21998(.O (g18866), .I1 (g13834), .I2 (g12069));
NR2X1 gate21999(.O (g18867), .I1 (g13835), .I2 (g12070));
NR2X1 gate22000(.O (g18868), .I1 (g14143), .I2 (g12419));
NR2X1 gate22001(.O (g18883), .I1 (g13846), .I2 (g12128));
NR2X1 gate22002(.O (g18885), .I1 (g13847), .I2 (g12129));
NR2X1 gate22003(.O (g18906), .I1 (g13855), .I2 (g12186));
NR2X1 gate22004(.O (g18907), .I1 (g14336), .I2 (g12429));
NR2X1 gate22005(.O (g18942), .I1 (g13870), .I2 (g12273));
NR2X1 gate22006(.O (g18957), .I1 (g13884), .I2 (g12307));
NR2X1 gate22007(.O (g18968), .I1 (g13904), .I2 (g12330));
NR2X1 gate22008(.O (g18975), .I1 (g13944), .I2 (g12353));
NR2X1 gate22009(.O (g19144), .I1 (g17268), .I2 (g14884));
NR2X1 gate22010(.O (g19149), .I1 (g17339), .I2 (g15020));
NR2X1 gate22011(.O (g19153), .I1 (g17381), .I2 (g15093));
NR2X1 gate22012(.O (g19154), .I1 (g17382), .I2 (g15094));
NR2X1 gate22013(.O (g19157), .I1 (g17428), .I2 (g15171));
NR2X1 gate22014(.O (g19160), .I1 (g17446), .I2 (g15178));
NR2X1 gate22015(.O (g19162), .I1 (g17485), .I2 (g15243));
NR2X1 gate22016(.O (g19163), .I1 (g17486), .I2 (g15244));
NR2X1 gate22017(.O (g19165), .I1 (g17526), .I2 (g15264));
NR2X1 gate22018(.O (g19167), .I1 (g17556), .I2 (g15320));
NR2X1 gate22019(.O (g19171), .I1 (g17616), .I2 (g15356));
NR2X1 gate22020(.O (g19172), .I1 (g17635), .I2 (g15388));
NR2X1 gate22021(.O (g19173), .I1 (g17636), .I2 (g15389));
NR2X1 gate22022(.O (g19177), .I1 (g17713), .I2 (g15442));
NR2X1 gate22023(.O (g19178), .I1 (g17718), .I2 (g15452));
NR2X1 gate22024(.O (g19179), .I1 (g17719), .I2 (g15453));
NR2X1 gate22025(.O (g19184), .I1 (g17798), .I2 (g15520));
NR2X1 gate22026(.O (g19219), .I1 (g18165), .I2 (g15753));
NR2X1 gate22027(.O (g20008), .I1 (g18977), .I2 (g7338));
NR2X1 gate22028(.O (g20054), .I1 (g19001), .I2 (g16867));
NR2X1 gate22029(.O (g20095), .I1 (g16507), .I2 (g16895));
NR2X1 gate22030(.O (g20120), .I1 (g16529), .I2 (g16924));
NR2X1 gate22031(.O (g20150), .I1 (g16560), .I2 (g16954));
NR2X1 gate22032(.O (g20153), .I1 (g16536), .I2 (g7583));
NR2X1 gate22033(.O (g20299), .I1 (g16665), .I2 (g16884));
NR2X1 gate22034(.O (g20310), .I1 (g16850), .I2 (g13654));
NR2X1 gate22035(.O (g20314), .I1 (g13646), .I2 (g16855));
NR2X1 gate22036(.O (g20318), .I1 (g16686), .I2 (g16913));
NR2X1 gate22037(.O (g20333), .I1 (g13672), .I2 (g16859));
NR2X1 gate22038(.O (g20337), .I1 (g16712), .I2 (g16943));
NR2X1 gate22039(.O (g20343), .I1 (g16856), .I2 (g13703));
NR2X1 gate22040(.O (g20353), .I1 (g13702), .I2 (g16864));
NR2X1 gate22041(.O (g20357), .I1 (g16743), .I2 (g16974));
NR2X1 gate22042(.O (g20375), .I1 (g13739), .I2 (g16879));
NR2X1 gate22043(.O (g20376), .I1 (g16865), .I2 (g13787));
NR2X1 gate22044(.O (g20417), .I1 (g16907), .I2 (g13833));
NR2X1 gate22045(.O (g20682), .I1 (g19160), .I2 (g10024));
NR2X1 gate22046(.O (g20717), .I1 (g19165), .I2 (g10133));
NR2X1 gate22047(.O (g20752), .I1 (g19171), .I2 (g10238));
NR2X1 gate22048(.O (g20789), .I1 (g19177), .I2 (g10340));
NR2X1 gate22049(.O (g20841), .I1 (g14767), .I2 (g19552));
NR2X1 gate22050(.O (g20874), .I1 (g17301), .I2 (g19594));
NR2X1 gate22051(.O (g20875), .I1 (g19584), .I2 (g17352));
NR2X1 gate22052(.O (g20876), .I1 (g19585), .I2 (g17353));
NR2X1 gate22053(.O (g20877), .I1 (g3919), .I2 (g19830));
NR2X1 gate22054(.O (g20878), .I1 (g19600), .I2 (g17395));
NR2X1 gate22055(.O (g20879), .I1 (g19601), .I2 (g17396));
NR2X1 gate22056(.O (g20880), .I1 (g19602), .I2 (g17397));
NR2X1 gate22057(.O (g20881), .I1 (g19603), .I2 (g17398));
NR2X1 gate22058(.O (g20882), .I1 (g19614), .I2 (g17408));
NR2X1 gate22059(.O (g20883), .I1 (g19615), .I2 (g17409));
NR2X1 gate22060(.O (g20884), .I1 (g5394), .I2 (g19830));
NR2X1 gate22061(.O (g20891), .I1 (g19626), .I2 (g17447));
NR2X1 gate22062(.O (g20892), .I1 (g19627), .I2 (g17448));
NR2X1 gate22063(.O (g20893), .I1 (g19628), .I2 (g17449));
NR2X1 gate22064(.O (g20894), .I1 (g19629), .I2 (g17450));
NR2X1 gate22065(.O (g20895), .I1 (g19633), .I2 (g17461));
NR2X1 gate22066(.O (g20896), .I1 (g19634), .I2 (g17462));
NR2X1 gate22067(.O (g20897), .I1 (g19635), .I2 (g17463));
NR2X1 gate22068(.O (g20898), .I1 (g19636), .I2 (g17464));
NR2X1 gate22069(.O (g20899), .I1 (g19647), .I2 (g17474));
NR2X1 gate22070(.O (g20900), .I1 (g19648), .I2 (g17475));
NR2X1 gate22071(.O (g20901), .I1 (g19660), .I2 (g17508));
NR2X1 gate22072(.O (g20902), .I1 (g19661), .I2 (g17509));
NR2X1 gate22073(.O (g20903), .I1 (g19662), .I2 (g17510));
NR2X1 gate22074(.O (g20910), .I1 (g19666), .I2 (g17527));
NR2X1 gate22075(.O (g20911), .I1 (g19667), .I2 (g17528));
NR2X1 gate22076(.O (g20912), .I1 (g19668), .I2 (g17529));
NR2X1 gate22077(.O (g20913), .I1 (g19669), .I2 (g17530));
NR2X1 gate22078(.O (g20914), .I1 (g19673), .I2 (g17541));
NR2X1 gate22079(.O (g20915), .I1 (g19674), .I2 (g17542));
NR2X1 gate22080(.O (g20916), .I1 (g19675), .I2 (g17543));
NR2X1 gate22081(.O (g20917), .I1 (g19676), .I2 (g17544));
NR2X1 gate22082(.O (g20918), .I1 (g19687), .I2 (g17554));
NR2X1 gate22083(.O (g20919), .I1 (g19688), .I2 (g17555));
NR2X1 gate22084(.O (g20920), .I1 (g19691), .I2 (g19726));
NR2X1 gate22085(.O (g20921), .I1 (g19697), .I2 (g17576));
NR2X1 gate22086(.O (g20922), .I1 (g19698), .I2 (g17577));
NR2X1 gate22087(.O (g20923), .I1 (g19699), .I2 (g17578));
NR2X1 gate22088(.O (g20924), .I1 (g19700), .I2 (g15257));
NR2X1 gate22089(.O (g20925), .I1 (g19708), .I2 (g17598));
NR2X1 gate22090(.O (g20926), .I1 (g19709), .I2 (g17599));
NR2X1 gate22091(.O (g20927), .I1 (g19710), .I2 (g17600));
NR2X1 gate22092(.O (g20934), .I1 (g19714), .I2 (g17617));
NR2X1 gate22093(.O (g20935), .I1 (g19715), .I2 (g17618));
NR2X1 gate22094(.O (g20936), .I1 (g19716), .I2 (g17619));
NR2X1 gate22095(.O (g20937), .I1 (g19717), .I2 (g17620));
NR2X1 gate22096(.O (g20938), .I1 (g19721), .I2 (g17631));
NR2X1 gate22097(.O (g20939), .I1 (g19722), .I2 (g17632));
NR2X1 gate22098(.O (g20940), .I1 (g19723), .I2 (g17633));
NR2X1 gate22099(.O (g20941), .I1 (g19724), .I2 (g17634));
NR2X1 gate22100(.O (g20944), .I1 (g19731), .I2 (g17652));
NR2X1 gate22101(.O (g20945), .I1 (g19732), .I2 (g17653));
NR2X1 gate22102(.O (g20946), .I1 (g19733), .I2 (g17654));
NR2X1 gate22103(.O (g20947), .I1 (g19734), .I2 (g15335));
NR2X1 gate22104(.O (g20948), .I1 (g19735), .I2 (g15336));
NR2X1 gate22105(.O (g20949), .I1 (g19741), .I2 (g17673));
NR2X1 gate22106(.O (g20950), .I1 (g19742), .I2 (g17674));
NR2X1 gate22107(.O (g20951), .I1 (g19743), .I2 (g17675));
NR2X1 gate22108(.O (g20952), .I1 (g19744), .I2 (g15349));
NR2X1 gate22109(.O (g20953), .I1 (g19752), .I2 (g17695));
NR2X1 gate22110(.O (g20954), .I1 (g19753), .I2 (g17696));
NR2X1 gate22111(.O (g20955), .I1 (g19754), .I2 (g17697));
NR2X1 gate22112(.O (g20962), .I1 (g19758), .I2 (g17714));
NR2X1 gate22113(.O (g20963), .I1 (g19759), .I2 (g17715));
NR2X1 gate22114(.O (g20964), .I1 (g19760), .I2 (g17716));
NR2X1 gate22115(.O (g20965), .I1 (g19761), .I2 (g17717));
NR2X1 gate22116(.O (g20966), .I1 (g19765), .I2 (g17734));
NR2X1 gate22117(.O (g20967), .I1 (g19766), .I2 (g17735));
NR2X1 gate22118(.O (g20968), .I1 (g19767), .I2 (g17736));
NR2X1 gate22119(.O (g20969), .I1 (g19768), .I2 (g15402));
NR2X1 gate22120(.O (g20970), .I1 (g19769), .I2 (g15403));
NR2X1 gate22121(.O (g20972), .I1 (g19774), .I2 (g17752));
NR2X1 gate22122(.O (g20973), .I1 (g19775), .I2 (g17753));
NR2X1 gate22123(.O (g20974), .I1 (g19776), .I2 (g17754));
NR2X1 gate22124(.O (g20975), .I1 (g19777), .I2 (g15421));
NR2X1 gate22125(.O (g20976), .I1 (g19778), .I2 (g15422));
NR2X1 gate22126(.O (g20977), .I1 (g19784), .I2 (g17773));
NR2X1 gate22127(.O (g20978), .I1 (g19785), .I2 (g17774));
NR2X1 gate22128(.O (g20979), .I1 (g19786), .I2 (g17775));
NR2X1 gate22129(.O (g20980), .I1 (g19787), .I2 (g15435));
NR2X1 gate22130(.O (g20981), .I1 (g19795), .I2 (g17795));
NR2X1 gate22131(.O (g20982), .I1 (g19796), .I2 (g17796));
NR2X1 gate22132(.O (g20983), .I1 (g19797), .I2 (g17797));
NR2X1 gate22133(.O (g20989), .I1 (g19802), .I2 (g17812));
NR2X1 gate22134(.O (g20990), .I1 (g19803), .I2 (g17813));
NR2X1 gate22135(.O (g20991), .I1 (g19804), .I2 (g17814));
NR2X1 gate22136(.O (g20992), .I1 (g19805), .I2 (g15470));
NR2X1 gate22137(.O (g20993), .I1 (g19807), .I2 (g17835));
NR2X1 gate22138(.O (g20994), .I1 (g19808), .I2 (g17836));
NR2X1 gate22139(.O (g20995), .I1 (g19809), .I2 (g17837));
NR2X1 gate22140(.O (g20996), .I1 (g19810), .I2 (g15486));
NR2X1 gate22141(.O (g20997), .I1 (g19811), .I2 (g15487));
NR2X1 gate22142(.O (g20999), .I1 (g19816), .I2 (g17853));
NR2X1 gate22143(.O (g21000), .I1 (g19817), .I2 (g17854));
NR2X1 gate22144(.O (g21001), .I1 (g19818), .I2 (g17855));
NR2X1 gate22145(.O (g21002), .I1 (g19819), .I2 (g15505));
NR2X1 gate22146(.O (g21003), .I1 (g19820), .I2 (g15506));
NR2X1 gate22147(.O (g21004), .I1 (g19826), .I2 (g17874));
NR2X1 gate22148(.O (g21005), .I1 (g19827), .I2 (g17875));
NR2X1 gate22149(.O (g21006), .I1 (g19828), .I2 (g17876));
NR2X1 gate22150(.O (g21007), .I1 (g19829), .I2 (g15519));
NR2X1 gate22151(.O (g21008), .I1 (g19836), .I2 (g17877));
NR2X1 gate22152(.O (g21009), .I1 (g19839), .I2 (g17900));
NR2X1 gate22153(.O (g21010), .I1 (g19840), .I2 (g17901));
NR2X1 gate22154(.O (g21011), .I1 (g19841), .I2 (g17902));
NR2X1 gate22155(.O (g21015), .I1 (g19846), .I2 (g17924));
NR2X1 gate22156(.O (g21016), .I1 (g19847), .I2 (g17925));
NR2X1 gate22157(.O (g21017), .I1 (g19848), .I2 (g17926));
NR2X1 gate22158(.O (g21018), .I1 (g19849), .I2 (g15556));
NR2X1 gate22159(.O (g21019), .I1 (g19851), .I2 (g17947));
NR2X1 gate22160(.O (g21020), .I1 (g19852), .I2 (g17948));
NR2X1 gate22161(.O (g21021), .I1 (g19853), .I2 (g17949));
NR2X1 gate22162(.O (g21022), .I1 (g19854), .I2 (g15572));
NR2X1 gate22163(.O (g21023), .I1 (g19855), .I2 (g15573));
NR2X1 gate22164(.O (g21025), .I1 (g19860), .I2 (g17965));
NR2X1 gate22165(.O (g21026), .I1 (g19861), .I2 (g17966));
NR2X1 gate22166(.O (g21027), .I1 (g19862), .I2 (g17967));
NR2X1 gate22167(.O (g21028), .I1 (g19863), .I2 (g15591));
NR2X1 gate22168(.O (g21029), .I1 (g19864), .I2 (g15592));
NR2X1 gate22169(.O (g21031), .I1 (g19869), .I2 (g17989));
NR2X1 gate22170(.O (g21032), .I1 (g19870), .I2 (g17990));
NR2X1 gate22171(.O (g21033), .I1 (g19872), .I2 (g18011));
NR2X1 gate22172(.O (g21034), .I1 (g19873), .I2 (g18012));
NR2X1 gate22173(.O (g21035), .I1 (g19874), .I2 (g18013));
NR2X1 gate22174(.O (g21039), .I1 (g19879), .I2 (g18035));
NR2X1 gate22175(.O (g21040), .I1 (g19880), .I2 (g18036));
NR2X1 gate22176(.O (g21041), .I1 (g19881), .I2 (g18037));
NR2X1 gate22177(.O (g21042), .I1 (g19882), .I2 (g15634));
NR2X1 gate22178(.O (g21043), .I1 (g19884), .I2 (g18058));
NR2X1 gate22179(.O (g21044), .I1 (g19885), .I2 (g18059));
NR2X1 gate22180(.O (g21045), .I1 (g19886), .I2 (g18060));
NR2X1 gate22181(.O (g21046), .I1 (g19887), .I2 (g15650));
NR2X1 gate22182(.O (g21047), .I1 (g19888), .I2 (g15651));
NR2X1 gate22183(.O (g21048), .I1 (g19889), .I2 (g18062));
NR2X1 gate22184(.O (g21051), .I1 (g19895), .I2 (g18088));
NR2X1 gate22185(.O (g21052), .I1 (g19900), .I2 (g18106));
NR2X1 gate22186(.O (g21053), .I1 (g19901), .I2 (g18107));
NR2X1 gate22187(.O (g21054), .I1 (g19903), .I2 (g18128));
NR2X1 gate22188(.O (g21055), .I1 (g19904), .I2 (g18129));
NR2X1 gate22189(.O (g21056), .I1 (g19905), .I2 (g18130));
NR2X1 gate22190(.O (g21060), .I1 (g19910), .I2 (g18152));
NR2X1 gate22191(.O (g21061), .I1 (g19911), .I2 (g18153));
NR2X1 gate22192(.O (g21062), .I1 (g19912), .I2 (g18154));
NR2X1 gate22193(.O (g21063), .I1 (g19913), .I2 (g15710));
NR2X1 gate22194(.O (g21065), .I1 (g19914), .I2 (g18169));
NR2X1 gate22195(.O (g21070), .I1 (g19920), .I2 (g18204));
NR2X1 gate22196(.O (g21071), .I1 (g19925), .I2 (g18222));
NR2X1 gate22197(.O (g21072), .I1 (g19926), .I2 (g18223));
NR2X1 gate22198(.O (g21073), .I1 (g19928), .I2 (g18244));
NR2X1 gate22199(.O (g21074), .I1 (g19929), .I2 (g18245));
NR2X1 gate22200(.O (g21075), .I1 (g19930), .I2 (g18246));
NR2X1 gate22201(.O (g21080), .I1 (g19935), .I2 (g18311));
NR2X1 gate22202(.O (g21081), .I1 (g19940), .I2 (g18329));
NR2X1 gate22203(.O (g21082), .I1 (g19941), .I2 (g18330));
NR2X1 gate22204(.O (g21083), .I1 (g19943), .I2 (g18333));
NR2X1 gate22205(.O (g21084), .I1 (g20011), .I2 (g20048));
NR2X1 gate22206(.O (g21094), .I1 (g19952), .I2 (g18404));
NR3X1 gate22207(.O (g21095), .I1 (g20012), .I2 (g20049), .I3 (g20084));
NR3X1 gate22208(.O (g21096), .I1 (g20013), .I2 (g20051), .I3 (g20087));
NR3X1 gate22209(.O (g21104), .I1 (g20050), .I2 (g20085), .I3 (g20106));
NR3X1 gate22210(.O (g21105), .I1 (g20052), .I2 (g20088), .I3 (g20109));
NR3X1 gate22211(.O (g21106), .I1 (g20053), .I2 (g20090), .I3 (g20112));
NR3X1 gate22212(.O (g21116), .I1 (g20086), .I2 (g20107), .I3 (g20131));
NR3X1 gate22213(.O (g21117), .I1 (g20089), .I2 (g20110), .I3 (g20133));
NR3X1 gate22214(.O (g21118), .I1 (g20091), .I2 (g20113), .I3 (g20136));
NR3X1 gate22215(.O (g21119), .I1 (g20092), .I2 (g20115), .I3 (g20139));
NR3X1 gate22216(.O (g21133), .I1 (g20108), .I2 (g20132), .I3 (g20156));
NR3X1 gate22217(.O (g21134), .I1 (g20111), .I2 (g20134), .I3 (g20157));
NR3X1 gate22218(.O (g21135), .I1 (g20114), .I2 (g20137), .I3 (g20160));
NR3X1 gate22219(.O (g21147), .I1 (g20135), .I2 (g20158), .I3 (g20188));
NR3X1 gate22220(.O (g21148), .I1 (g20138), .I2 (g20161), .I3 (g20190));
NR2X1 gate22221(.O (g21149), .I1 (g20015), .I2 (g19981));
NR2X1 gate22222(.O (g21167), .I1 (g20159), .I2 (g20189));
NR3X1 gate22223(.O (g21168), .I1 (g20162), .I2 (g20191), .I3 (g20220));
NR2X1 gate22224(.O (g21169), .I1 (g20057), .I2 (g20019));
NR2X1 gate22225(.O (g21183), .I1 (g20192), .I2 (g20221));
NR2X1 gate22226(.O (g21189), .I1 (g20098), .I2 (g20061));
NR2X1 gate22227(.O (g21204), .I1 (g20123), .I2 (g20102));
NR2X1 gate22228(.O (g21211), .I1 (g19240), .I2 (g19230));
NR2X1 gate22229(.O (g21219), .I1 (g19253), .I2 (g19243));
NR3X1 gate22230(.O (g21227), .I1 (g18414), .I2 (g18485), .I3 (g20295));
NR2X1 gate22231(.O (g21228), .I1 (g19388), .I2 (g17118));
NR2X1 gate22232(.O (g21230), .I1 (g19266), .I2 (g19256));
NR2X1 gate22233(.O (g21233), .I1 (g19418), .I2 (g17145));
NR2X1 gate22234(.O (g21235), .I1 (g19281), .I2 (g19269));
NR2X1 gate22235(.O (g21238), .I1 (g19954), .I2 (g5890));
NR2X1 gate22236(.O (g21242), .I1 (g19455), .I2 (g17168));
NR2X1 gate22237(.O (g21246), .I1 (g19984), .I2 (g5929));
NR2X1 gate22238(.O (g21250), .I1 (g19482), .I2 (g17183));
NR2X1 gate22239(.O (g21255), .I1 (g20022), .I2 (g5963));
NR2X1 gate22240(.O (g21263), .I1 (g20064), .I2 (g5992));
NR2X1 gate22241(.O (g21316), .I1 (g20460), .I2 (g16111));
NR2X1 gate22242(.O (g21331), .I1 (g20472), .I2 (g16153));
NR2X1 gate22243(.O (g21346), .I1 (g20480), .I2 (g13247));
NR2X1 gate22244(.O (g21364), .I1 (g20486), .I2 (g13266));
NR2X1 gate22245(.O (g21385), .I1 (g20492), .I2 (g13289));
NR2X1 gate22246(.O (g21407), .I1 (g20499), .I2 (g13316));
NR2X1 gate22247(.O (g21432), .I1 (g20502), .I2 (g13335));
NR2X1 gate22248(.O (g21435), .I1 (g20503), .I2 (g16385));
NR2X1 gate22249(.O (g21467), .I1 (g20506), .I2 (g13355));
NR2X1 gate22250(.O (g21470), .I1 (g20512), .I2 (g16417));
NR2X1 gate22251(.O (g21502), .I1 (g20525), .I2 (g16445));
NR2X1 gate22252(.O (g21615), .I1 (g16567), .I2 (g19957));
NR3X1 gate22253(.O (g21618), .I1 (g20016), .I2 (g14079), .I3 (g14165));
NR2X1 gate22254(.O (g21636), .I1 (g20473), .I2 (g6513));
NR2X1 gate22255(.O (g21643), .I1 (g16591), .I2 (g19987));
NR3X1 gate22256(.O (g21646), .I1 (g20058), .I2 (g14194), .I3 (g14280));
NR2X1 gate22257(.O (g21665), .I1 (g20507), .I2 (g18352));
NR2X1 gate22258(.O (g21667), .I1 (g20481), .I2 (g6777));
NR2X1 gate22259(.O (g21674), .I1 (g16611), .I2 (g20025));
NR3X1 gate22260(.O (g21677), .I1 (g20099), .I2 (g14309), .I3 (g14402));
NR2X1 gate22261(.O (g21694), .I1 (g20526), .I2 (g18447));
NR2X1 gate22262(.O (g21696), .I1 (g20487), .I2 (g7079));
NR2X1 gate22263(.O (g21703), .I1 (g16629), .I2 (g20067));
NR3X1 gate22264(.O (g21706), .I1 (g20124), .I2 (g14431), .I3 (g14514));
NR2X1 gate22265(.O (g21711), .I1 (g19830), .I2 (g15780));
NR2X1 gate22266(.O (g21730), .I1 (g20545), .I2 (g18520));
NR2X1 gate22267(.O (g21732), .I1 (g20493), .I2 (g7329));
NR3X1 gate22268(.O (g21738), .I1 (g19444), .I2 (g17893), .I3 (g14079));
NR2X1 gate22269(.O (g21739), .I1 (g20507), .I2 (g18430));
NR2X1 gate22270(.O (g21756), .I1 (g19070), .I2 (g18584));
NR3X1 gate22271(.O (g21762), .I1 (g19471), .I2 (g18004), .I3 (g14194));
NR2X1 gate22272(.O (g21763), .I1 (g20526), .I2 (g18503));
NR3X1 gate22273(.O (g21778), .I1 (g19494), .I2 (g18121), .I3 (g14309));
NR2X1 gate22274(.O (g21779), .I1 (g20545), .I2 (g18567));
NR3X1 gate22275(.O (g21793), .I1 (g19515), .I2 (g18237), .I3 (g14431));
NR2X1 gate22276(.O (g21794), .I1 (g19070), .I2 (g18617));
NR2X1 gate22277(.O (g21796), .I1 (g19830), .I2 (g13004));
NR2X1 gate22278(.O (g21842), .I1 (g13609), .I2 (g19150));
NR2X1 gate22279(.O (g21843), .I1 (g13619), .I2 (g19155));
NR2X1 gate22280(.O (g21845), .I1 (g13631), .I2 (g19161));
NR2X1 gate22281(.O (g21847), .I1 (g13642), .I2 (g19166));
NR2X1 gate22282(.O (g21851), .I1 (g19252), .I2 (g8842));
NR2X1 gate22283(.O (g21878), .I1 (g16964), .I2 (g19228));
NR2X1 gate22284(.O (g21880), .I1 (g13854), .I2 (g19236));
NR2X1 gate22285(.O (g21882), .I1 (g13862), .I2 (g19248));
NR2X1 gate22286(.O (g21884), .I1 (g19260), .I2 (g19284));
NR2X1 gate22287(.O (g21887), .I1 (g13519), .I2 (g19289));
NR2X1 gate22288(.O (g21889), .I1 (g19285), .I2 (g19316));
NR2X1 gate22289(.O (g21890), .I1 (g13530), .I2 (g19307));
NR2X1 gate22290(.O (g21893), .I1 (g13541), .I2 (g19328));
NR2X1 gate22291(.O (g21894), .I1 (g19317), .I2 (g19356));
NR2X1 gate22292(.O (g21901), .I1 (g13552), .I2 (g19355));
NR2X1 gate22293(.O (g21968), .I1 (g21234), .I2 (g19476));
NR2X1 gate22294(.O (g21969), .I1 (g20895), .I2 (g10133));
NR2X1 gate22295(.O (g21970), .I1 (g17182), .I2 (g21226));
NR2X1 gate22296(.O (g21971), .I1 (g21243), .I2 (g19499));
NR2X1 gate22297(.O (g21972), .I1 (g20914), .I2 (g10238));
NR2X1 gate22298(.O (g21973), .I1 (g21251), .I2 (g19520));
NR2X1 gate22299(.O (g21974), .I1 (g20938), .I2 (g10340));
NR2X1 gate22300(.O (g21975), .I1 (g21245), .I2 (g21259));
NR3X1 gate22301(.O (g21980), .I1 (g21252), .I2 (g19531), .I3 (g19540));
NR2X1 gate22302(.O (g21981), .I1 (g21254), .I2 (g21267));
NR3X1 gate22303(.O (g21987), .I1 (g21260), .I2 (g19541), .I3 (g19544));
NR2X1 gate22304(.O (g21988), .I1 (g21262), .I2 (g21276));
NR3X1 gate22305(.O (g22000), .I1 (g21268), .I2 (g19545), .I3 (g19547));
NR2X1 gate22306(.O (g22001), .I1 (g21270), .I2 (g21283));
NR3X1 gate22307(.O (g22013), .I1 (g21277), .I2 (g19548), .I3 (g19551));
NR2X1 gate22308(.O (g22025), .I1 (g21284), .I2 (g19549));
NR2X1 gate22309(.O (g22026), .I1 (g21083), .I2 (g18407));
NR2X1 gate22310(.O (g22027), .I1 (g21290), .I2 (g19553));
NR2X1 gate22311(.O (g22028), .I1 (g21291), .I2 (g19554));
NR2X1 gate22312(.O (g22029), .I1 (g21292), .I2 (g19555));
NR2X1 gate22313(.O (g22030), .I1 (g21298), .I2 (g19557));
NR2X1 gate22314(.O (g22031), .I1 (g21299), .I2 (g19558));
NR2X1 gate22315(.O (g22032), .I1 (g21300), .I2 (g19559));
NR2X1 gate22316(.O (g22033), .I1 (g21301), .I2 (g19560));
NR2X1 gate22317(.O (g22034), .I1 (g21302), .I2 (g19561));
NR2X1 gate22318(.O (g22035), .I1 (g21303), .I2 (g19562));
NR2X1 gate22319(.O (g22037), .I1 (g21304), .I2 (g19564));
NR2X1 gate22320(.O (g22038), .I1 (g21305), .I2 (g19565));
NR2X1 gate22321(.O (g22039), .I1 (g21306), .I2 (g19566));
NR2X1 gate22322(.O (g22040), .I1 (g21307), .I2 (g19567));
NR2X1 gate22323(.O (g22041), .I1 (g21308), .I2 (g19568));
NR2X1 gate22324(.O (g22042), .I1 (g21309), .I2 (g19569));
NR2X1 gate22325(.O (g22043), .I1 (g21310), .I2 (g19570));
NR2X1 gate22326(.O (g22044), .I1 (g21311), .I2 (g19571));
NR2X1 gate22327(.O (g22045), .I1 (g21312), .I2 (g19572));
NR2X1 gate22328(.O (g22047), .I1 (g21313), .I2 (g19574));
NR2X1 gate22329(.O (g22048), .I1 (g21314), .I2 (g19575));
NR2X1 gate22330(.O (g22049), .I1 (g21315), .I2 (g19576));
NR2X1 gate22331(.O (g22054), .I1 (g21319), .I2 (g19586));
NR2X1 gate22332(.O (g22055), .I1 (g21320), .I2 (g19587));
NR2X1 gate22333(.O (g22056), .I1 (g21321), .I2 (g19588));
NR2X1 gate22334(.O (g22057), .I1 (g21322), .I2 (g19589));
NR2X1 gate22335(.O (g22058), .I1 (g21323), .I2 (g19590));
NR2X1 gate22336(.O (g22059), .I1 (g21324), .I2 (g19591));
NR2X1 gate22337(.O (g22060), .I1 (g21325), .I2 (g19592));
NR2X1 gate22338(.O (g22061), .I1 (g21326), .I2 (g19593));
NR2X1 gate22339(.O (g22063), .I1 (g21328), .I2 (g19597));
NR2X1 gate22340(.O (g22064), .I1 (g21329), .I2 (g19598));
NR2X1 gate22341(.O (g22065), .I1 (g21330), .I2 (g19599));
NR2X1 gate22342(.O (g22066), .I1 (g21334), .I2 (g19604));
NR2X1 gate22343(.O (g22067), .I1 (g21335), .I2 (g19605));
NR2X1 gate22344(.O (g22068), .I1 (g21336), .I2 (g19606));
NR2X1 gate22345(.O (g22073), .I1 (g21337), .I2 (g19616));
NR2X1 gate22346(.O (g22074), .I1 (g21338), .I2 (g19617));
NR2X1 gate22347(.O (g22075), .I1 (g21339), .I2 (g19618));
NR2X1 gate22348(.O (g22076), .I1 (g21340), .I2 (g19619));
NR2X1 gate22349(.O (g22077), .I1 (g21341), .I2 (g19620));
NR2X1 gate22350(.O (g22078), .I1 (g21342), .I2 (g19621));
NR2X1 gate22351(.O (g22079), .I1 (g21343), .I2 (g19623));
NR2X1 gate22352(.O (g22080), .I1 (g21344), .I2 (g19624));
NR2X1 gate22353(.O (g22081), .I1 (g21345), .I2 (g19625));
NR2X1 gate22354(.O (g22087), .I1 (g21349), .I2 (g19630));
NR2X1 gate22355(.O (g22088), .I1 (g21350), .I2 (g19631));
NR2X1 gate22356(.O (g22089), .I1 (g21351), .I2 (g19632));
NR2X1 gate22357(.O (g22090), .I1 (g21352), .I2 (g19637));
NR2X1 gate22358(.O (g22091), .I1 (g21353), .I2 (g19638));
NR2X1 gate22359(.O (g22092), .I1 (g21354), .I2 (g19639));
NR2X1 gate22360(.O (g22097), .I1 (g21355), .I2 (g19649));
NR2X1 gate22361(.O (g22098), .I1 (g21356), .I2 (g19650));
NR2X1 gate22362(.O (g22099), .I1 (g21357), .I2 (g19651));
NR2X1 gate22363(.O (g22100), .I1 (g21360), .I2 (g19653));
NR2X1 gate22364(.O (g22101), .I1 (g21361), .I2 (g19654));
NR2X1 gate22365(.O (g22102), .I1 (g21362), .I2 (g19655));
NR2X1 gate22366(.O (g22103), .I1 (g21363), .I2 (g19656));
NR2X1 gate22367(.O (g22104), .I1 (g21367), .I2 (g19663));
NR2X1 gate22368(.O (g22105), .I1 (g21368), .I2 (g19664));
NR2X1 gate22369(.O (g22106), .I1 (g21369), .I2 (g19665));
NR2X1 gate22370(.O (g22112), .I1 (g21370), .I2 (g19670));
NR2X1 gate22371(.O (g22113), .I1 (g21371), .I2 (g19671));
NR2X1 gate22372(.O (g22114), .I1 (g21372), .I2 (g19672));
NR2X1 gate22373(.O (g22115), .I1 (g21373), .I2 (g19677));
NR2X1 gate22374(.O (g22116), .I1 (g21374), .I2 (g19678));
NR2X1 gate22375(.O (g22117), .I1 (g21375), .I2 (g19679));
NR2X1 gate22376(.O (g22122), .I1 (g21378), .I2 (g19692));
NR2X1 gate22377(.O (g22123), .I1 (g21379), .I2 (g19693));
NR2X1 gate22378(.O (g22124), .I1 (g21380), .I2 (g19694));
NR2X1 gate22379(.O (g22125), .I1 (g21381), .I2 (g19695));
NR2X1 gate22380(.O (g22126), .I1 (g21389), .I2 (g19701));
NR2X1 gate22381(.O (g22127), .I1 (g21390), .I2 (g19702));
NR2X1 gate22382(.O (g22128), .I1 (g21391), .I2 (g19703));
NR2X1 gate22383(.O (g22129), .I1 (g21392), .I2 (g19704));
NR2X1 gate22384(.O (g22130), .I1 (g21393), .I2 (g19711));
NR2X1 gate22385(.O (g22131), .I1 (g21394), .I2 (g19712));
NR2X1 gate22386(.O (g22132), .I1 (g21395), .I2 (g19713));
NR2X1 gate22387(.O (g22138), .I1 (g21396), .I2 (g19718));
NR2X1 gate22388(.O (g22139), .I1 (g21397), .I2 (g19719));
NR2X1 gate22389(.O (g22140), .I1 (g21398), .I2 (g19720));
NR2X1 gate22390(.O (g22141), .I1 (g21401), .I2 (g19727));
NR2X1 gate22391(.O (g22142), .I1 (g21402), .I2 (g19728));
NR2X1 gate22392(.O (g22143), .I1 (g21403), .I2 (g19729));
NR2X1 gate22393(.O (g22144), .I1 (g21410), .I2 (g19730));
NR2X1 gate22394(.O (g22145), .I1 (g21411), .I2 (g19736));
NR2X1 gate22395(.O (g22146), .I1 (g21412), .I2 (g19737));
NR2X1 gate22396(.O (g22147), .I1 (g21413), .I2 (g19738));
NR2X1 gate22397(.O (g22148), .I1 (g21414), .I2 (g19739));
NR2X1 gate22398(.O (g22149), .I1 (g21419), .I2 (g19745));
NR2X1 gate22399(.O (g22150), .I1 (g21420), .I2 (g19746));
NR2X1 gate22400(.O (g22151), .I1 (g21421), .I2 (g19747));
NR2X1 gate22401(.O (g22152), .I1 (g21422), .I2 (g19748));
NR2X1 gate22402(.O (g22153), .I1 (g21423), .I2 (g19755));
NR2X1 gate22403(.O (g22154), .I1 (g21424), .I2 (g19756));
NR2X1 gate22404(.O (g22155), .I1 (g21425), .I2 (g19757));
NR2X1 gate22405(.O (g22161), .I1 (g21428), .I2 (g19764));
NR2X1 gate22406(.O (g22162), .I1 (g21438), .I2 (g19770));
NR2X1 gate22407(.O (g22163), .I1 (g21439), .I2 (g19771));
NR2X1 gate22408(.O (g22164), .I1 (g21440), .I2 (g19772));
NR2X1 gate22409(.O (g22165), .I1 (g21444), .I2 (g19773));
NR2X1 gate22410(.O (g22166), .I1 (g21445), .I2 (g19779));
NR2X1 gate22411(.O (g22167), .I1 (g21446), .I2 (g19780));
NR2X1 gate22412(.O (g22168), .I1 (g21447), .I2 (g19781));
NR2X1 gate22413(.O (g22169), .I1 (g21448), .I2 (g19782));
NR2X1 gate22414(.O (g22170), .I1 (g21453), .I2 (g19788));
NR2X1 gate22415(.O (g22171), .I1 (g21454), .I2 (g19789));
NR2X1 gate22416(.O (g22172), .I1 (g21455), .I2 (g19790));
NR2X1 gate22417(.O (g22173), .I1 (g21456), .I2 (g19791));
NR2X1 gate22418(.O (g22174), .I1 (g19868), .I2 (g21593));
NR2X1 gate22419(.O (g22177), .I1 (g21476), .I2 (g19806));
NR2X1 gate22420(.O (g22178), .I1 (g21480), .I2 (g19812));
NR2X1 gate22421(.O (g22179), .I1 (g21481), .I2 (g19813));
NR2X1 gate22422(.O (g22180), .I1 (g21482), .I2 (g19814));
NR2X1 gate22423(.O (g22181), .I1 (g21486), .I2 (g19815));
NR2X1 gate22424(.O (g22182), .I1 (g21487), .I2 (g19821));
NR2X1 gate22425(.O (g22183), .I1 (g21488), .I2 (g19822));
NR2X1 gate22426(.O (g22184), .I1 (g21489), .I2 (g19823));
NR2X1 gate22427(.O (g22185), .I1 (g21490), .I2 (g19824));
NR2X1 gate22428(.O (g22186), .I1 (g21497), .I2 (g19837));
NR2X1 gate22429(.O (g22189), .I1 (g19899), .I2 (g21622));
NR2X1 gate22430(.O (g22191), .I1 (g21517), .I2 (g19850));
NR2X1 gate22431(.O (g22192), .I1 (g21521), .I2 (g19856));
NR2X1 gate22432(.O (g22193), .I1 (g21522), .I2 (g19857));
NR2X1 gate22433(.O (g22194), .I1 (g21523), .I2 (g19858));
NR2X1 gate22434(.O (g22195), .I1 (g21527), .I2 (g19859));
NR2X1 gate22435(.O (g22198), .I1 (g19924), .I2 (g21650));
NR2X1 gate22436(.O (g22200), .I1 (g21553), .I2 (g19883));
NR2X1 gate22437(.O (g22204), .I1 (g19939), .I2 (g21681));
NR2X1 gate22438(.O (g22210), .I1 (g21610), .I2 (g19932));
NR2X1 gate22439(.O (g22216), .I1 (g21635), .I2 (g19944));
NR2X1 gate22440(.O (g22218), .I1 (g21639), .I2 (g19949));
NR2X1 gate22441(.O (g22227), .I1 (g21658), .I2 (g19953));
NR2X1 gate22442(.O (g22231), .I1 (g21666), .I2 (g19971));
NR2X1 gate22443(.O (g22234), .I1 (g21670), .I2 (g19976));
NR2X1 gate22444(.O (g22242), .I1 (g21687), .I2 (g19983));
NR2X1 gate22445(.O (g22247), .I1 (g21695), .I2 (g20001));
NR2X1 gate22446(.O (g22249), .I1 (g21699), .I2 (g20006));
NR2X1 gate22447(.O (g22263), .I1 (g21723), .I2 (g20021));
NR2X1 gate22448(.O (g22267), .I1 (g21731), .I2 (g20039));
NR2X1 gate22449(.O (g22269), .I1 (g21735), .I2 (g20044));
NR2X1 gate22450(.O (g22280), .I1 (g21749), .I2 (g20063));
NR2X1 gate22451(.O (g22284), .I1 (g21757), .I2 (g20081));
NR2X1 gate22452(.O (g22288), .I1 (g20144), .I2 (g21805));
NR2X1 gate22453(.O (g22299), .I1 (g21773), .I2 (g20104));
NR2X1 gate22454(.O (g22308), .I1 (g20182), .I2 (g21812));
NR2X1 gate22455(.O (g22336), .I1 (g20216), .I2 (g21818));
NR2X1 gate22456(.O (g22361), .I1 (g20246), .I2 (g21822));
NR2X1 gate22457(.O (g22454), .I1 (g17012), .I2 (g21891));
NR2X1 gate22458(.O (g22493), .I1 (g17042), .I2 (g21899));
NR2X1 gate22459(.O (g22536), .I1 (g17076), .I2 (g21911));
NR2X1 gate22460(.O (g22576), .I1 (g17111), .I2 (g21925));
NR2X1 gate22461(.O (g22578), .I1 (g21892), .I2 (g18982));
NR2X1 gate22462(.O (g22615), .I1 (g21900), .I2 (g18990));
NR2X1 gate22463(.O (g22651), .I1 (g21912), .I2 (g18997));
NR2X1 gate22464(.O (g22687), .I1 (g21926), .I2 (g19010));
NR2X1 gate22465(.O (g22755), .I1 (g21271), .I2 (g20842));
NR2X1 gate22466(.O (g22784), .I1 (g16075), .I2 (g20885));
NR2X1 gate22467(.O (g22789), .I1 (g21278), .I2 (g20850));
NR3X1 gate22468(.O (g22810), .I1 (g16075), .I2 (g20842), .I3 (g21271));
NR2X1 gate22469(.O (g22826), .I1 (g16113), .I2 (g20904));
NR2X1 gate22470(.O (g22831), .I1 (g21285), .I2 (g20858));
NR3X1 gate22471(.O (g22851), .I1 (g16113), .I2 (g20850), .I3 (g21278));
NR2X1 gate22472(.O (g22865), .I1 (g16164), .I2 (g20928));
NR2X1 gate22473(.O (g22870), .I1 (g21293), .I2 (g20866));
NR3X1 gate22474(.O (g22886), .I1 (g16164), .I2 (g20858), .I3 (g21285));
NR2X1 gate22475(.O (g22900), .I1 (g16223), .I2 (g20956));
NR3X1 gate22476(.O (g22921), .I1 (g16223), .I2 (g20866), .I3 (g21293));
NR2X1 gate22477(.O (g22935), .I1 (g21903), .I2 (g7466));
NR2X1 gate22478(.O (g22953), .I1 (g20700), .I2 (g7595));
NR2X1 gate22479(.O (g22985), .I1 (g21618), .I2 (g21049));
NR2X1 gate22480(.O (g22987), .I1 (g21646), .I2 (g21068));
NR2X1 gate22481(.O (g22990), .I1 (g21677), .I2 (g21078));
NR2X1 gate22482(.O (g22997), .I1 (g21706), .I2 (g21092));
NR2X1 gate22483(.O (g22999), .I1 (g21085), .I2 (g19241));
NR2X1 gate22484(.O (g23000), .I1 (g16909), .I2 (g21067));
NR2X1 gate22485(.O (g23009), .I1 (g21738), .I2 (g21107));
NR2X1 gate22486(.O (g23013), .I1 (g21097), .I2 (g19254));
NR2X1 gate22487(.O (g23014), .I1 (g16939), .I2 (g21077));
NR2X1 gate22488(.O (g23022), .I1 (g16968), .I2 (g21086));
NR3X1 gate22489(.O (g23023), .I1 (g14256), .I2 (g14175), .I3 (g21123));
NR2X1 gate22490(.O (g23025), .I1 (g21762), .I2 (g21124));
NR2X1 gate22491(.O (g23029), .I1 (g21111), .I2 (g19267));
NR2X1 gate22492(.O (g23030), .I1 (g16970), .I2 (g21091));
NR2X1 gate22493(.O (g23039), .I1 (g16989), .I2 (g21098));
NR3X1 gate22494(.O (g23040), .I1 (g14378), .I2 (g14290), .I3 (g21142));
NR2X1 gate22495(.O (g23042), .I1 (g21778), .I2 (g21143));
NR2X1 gate22496(.O (g23046), .I1 (g21128), .I2 (g19282));
NR2X1 gate22497(.O (g23047), .I1 (g16991), .I2 (g21103));
NR2X1 gate22498(.O (g23051), .I1 (g21121), .I2 (g21153));
NR2X1 gate22499(.O (g23058), .I1 (g16999), .I2 (g21112));
NR3X1 gate22500(.O (g23059), .I1 (g14490), .I2 (g14412), .I3 (g21162));
NR2X1 gate22501(.O (g23061), .I1 (g21793), .I2 (g21163));
NR3X1 gate22502(.O (g23066), .I1 (g21138), .I2 (g19303), .I3 (g19320));
NR2X1 gate22503(.O (g23067), .I1 (g17015), .I2 (g21122));
NR2X1 gate22504(.O (g23070), .I1 (g21140), .I2 (g21173));
NR2X1 gate22505(.O (g23076), .I1 (g17023), .I2 (g21129));
NR3X1 gate22506(.O (g23077), .I1 (g14577), .I2 (g14524), .I3 (g21182));
NR3X1 gate22507(.O (g23080), .I1 (g21158), .I2 (g19324), .I3 (g19347));
NR2X1 gate22508(.O (g23081), .I1 (g17045), .I2 (g21141));
NR2X1 gate22509(.O (g23083), .I1 (g21160), .I2 (g21193));
NR2X1 gate22510(.O (g23092), .I1 (g17055), .I2 (g21154));
NR2X1 gate22511(.O (g23093), .I1 (g17056), .I2 (g21155));
NR3X1 gate22512(.O (g23096), .I1 (g21178), .I2 (g19351), .I3 (g19381));
NR2X1 gate22513(.O (g23097), .I1 (g17079), .I2 (g21161));
NR2X1 gate22514(.O (g23099), .I1 (g21180), .I2 (g21208));
NR2X1 gate22515(.O (g23110), .I1 (g17090), .I2 (g21174));
NR2X1 gate22516(.O (g23111), .I1 (g17091), .I2 (g21175));
NR3X1 gate22517(.O (g23113), .I1 (g21198), .I2 (g19385), .I3 (g19413));
NR2X1 gate22518(.O (g23114), .I1 (g17114), .I2 (g21181));
NR2X1 gate22519(.O (g23117), .I1 (g17117), .I2 (g21188));
NR2X1 gate22520(.O (g23123), .I1 (g17128), .I2 (g21194));
NR2X1 gate22521(.O (g23124), .I1 (g17129), .I2 (g21195));
NR2X1 gate22522(.O (g23126), .I1 (g17144), .I2 (g21203));
NR2X1 gate22523(.O (g23132), .I1 (g17155), .I2 (g21209));
NR2X1 gate22524(.O (g23133), .I1 (g17156), .I2 (g21210));
NR2X1 gate22525(.O (g23135), .I1 (g21229), .I2 (g19449));
NR2X1 gate22526(.O (g23136), .I1 (g20878), .I2 (g10024));
NR2X1 gate22527(.O (g23137), .I1 (g17167), .I2 (g21218));
NR2X1 gate22528(.O (g23324), .I1 (g22144), .I2 (g10024));
NR2X1 gate22529(.O (g23329), .I1 (g22165), .I2 (g10133));
NR2X1 gate22530(.O (g23330), .I1 (g22186), .I2 (g22777));
NR2X1 gate22531(.O (g23339), .I1 (g22181), .I2 (g10238));
NR2X1 gate22532(.O (g23348), .I1 (g22195), .I2 (g10340));
NR2X1 gate22533(.O (g23357), .I1 (g22210), .I2 (g20127));
NR2X1 gate22534(.O (g23358), .I1 (g22227), .I2 (g18407));
NR2X1 gate22535(.O (g23359), .I1 (g22216), .I2 (g22907));
NR2X1 gate22536(.O (g23385), .I1 (g17393), .I2 (g22517));
NR2X1 gate22537(.O (g23386), .I1 (g22483), .I2 (g21388));
NR2X1 gate22538(.O (g23392), .I1 (g17460), .I2 (g22557));
NR2X1 gate22539(.O (g23393), .I1 (g22526), .I2 (g21418));
NR2X1 gate22540(.O (g23399), .I1 (g17506), .I2 (g22581));
NR2X1 gate22541(.O (g23400), .I1 (g17540), .I2 (g22597));
NR2X1 gate22542(.O (g23401), .I1 (g22566), .I2 (g21452));
NR2X1 gate22543(.O (g23406), .I1 (g17597), .I2 (g22618));
NR2X1 gate22544(.O (g23407), .I1 (g17630), .I2 (g22634));
NR2X1 gate22545(.O (g23408), .I1 (g22606), .I2 (g21494));
NR2X1 gate22546(.O (g23413), .I1 (g17694), .I2 (g22654));
NR2X1 gate22547(.O (g23418), .I1 (g17794), .I2 (g22690));
NR2X1 gate22548(.O (g23427), .I1 (g22699), .I2 (g21589));
NR2X1 gate22549(.O (g23433), .I1 (g22726), .I2 (g21611));
NR2X1 gate22550(.O (g23461), .I1 (g22841), .I2 (g21707));
NR2X1 gate22551(.O (g23477), .I1 (g22906), .I2 (g21758));
NR2X1 gate22552(.O (g23497), .I1 (g22876), .I2 (g5606));
NR2X1 gate22553(.O (g23513), .I1 (g22911), .I2 (g5631));
NR2X1 gate22554(.O (g23528), .I1 (g22936), .I2 (g5659));
NR2X1 gate22555(.O (g23539), .I1 (g22942), .I2 (g5697));
NR2X1 gate22556(.O (g23545), .I1 (g22984), .I2 (g20285));
NR3X1 gate22557(.O (g23823), .I1 (g23009), .I2 (g18490), .I3 (g4456));
NR3X1 gate22558(.O (g23858), .I1 (g23025), .I2 (g18554), .I3 (g4632));
NR3X1 gate22559(.O (g23892), .I1 (g23042), .I2 (g18604), .I3 (g4809));
NR3X1 gate22560(.O (g23913), .I1 (g23061), .I2 (g18636), .I3 (g4985));
NR2X1 gate22561(.O (g23922), .I1 (g4456), .I2 (g22985));
NR3X1 gate22562(.O (g23945), .I1 (g4456), .I2 (g13565), .I3 (g23009));
NR2X1 gate22563(.O (g23950), .I1 (g22992), .I2 (g6707));
NR2X1 gate22564(.O (g23954), .I1 (g4632), .I2 (g22987));
NR3X1 gate22565(.O (g23974), .I1 (g4632), .I2 (g13573), .I3 (g23025));
NR2X1 gate22566(.O (g23979), .I1 (g23003), .I2 (g7009));
NR2X1 gate22567(.O (g23983), .I1 (g4809), .I2 (g22990));
NR3X1 gate22568(.O (g24004), .I1 (g4809), .I2 (g13582), .I3 (g23042));
NR2X1 gate22569(.O (g24009), .I1 (g23017), .I2 (g7259));
NR2X1 gate22570(.O (g24013), .I1 (g4985), .I2 (g22997));
NR3X1 gate22571(.O (g24038), .I1 (g4985), .I2 (g13602), .I3 (g23061));
NR2X1 gate22572(.O (g24043), .I1 (g23033), .I2 (g7455));
NR2X1 gate22573(.O (g24059), .I1 (g21990), .I2 (g20809));
NR2X1 gate22574(.O (g24072), .I1 (g22004), .I2 (g20826));
NR2X1 gate22575(.O (g24083), .I1 (g22015), .I2 (g20836));
NR2X1 gate22576(.O (g24092), .I1 (g22020), .I2 (g20840));
NR2X1 gate22577(.O (g24174), .I1 (g16894), .I2 (g22206));
NR2X1 gate22578(.O (g24178), .I1 (g16908), .I2 (g22211));
NR2X1 gate22579(.O (g24179), .I1 (g16923), .I2 (g22214));
NR2X1 gate22580(.O (g24181), .I1 (g16938), .I2 (g22220));
NR2X1 gate22581(.O (g24182), .I1 (g16953), .I2 (g22223));
NR2X1 gate22582(.O (g24206), .I1 (g16966), .I2 (g22228));
NR2X1 gate22583(.O (g24207), .I1 (g16967), .I2 (g22229));
NR2X1 gate22584(.O (g24208), .I1 (g16969), .I2 (g22235));
NR2X1 gate22585(.O (g24209), .I1 (g16984), .I2 (g22238));
NR2X1 gate22586(.O (g24212), .I1 (g16987), .I2 (g22244));
NR2X1 gate22587(.O (g24213), .I1 (g16988), .I2 (g22245));
NR2X1 gate22588(.O (g24214), .I1 (g16990), .I2 (g22250));
NR2X1 gate22589(.O (g24215), .I1 (g16993), .I2 (g22254));
NR2X1 gate22590(.O (g24216), .I1 (g16994), .I2 (g22255));
NR2X1 gate22591(.O (g24218), .I1 (g16997), .I2 (g22264));
NR2X1 gate22592(.O (g24219), .I1 (g16998), .I2 (g22265));
NR2X1 gate22593(.O (g24222), .I1 (g17017), .I2 (g22272));
NR2X1 gate22594(.O (g24223), .I1 (g17018), .I2 (g22273));
NR2X1 gate22595(.O (g24225), .I1 (g17021), .I2 (g22281));
NR2X1 gate22596(.O (g24226), .I1 (g17022), .I2 (g22282));
NR2X1 gate22597(.O (g24227), .I1 (g22270), .I2 (g21137));
NR2X1 gate22598(.O (g24228), .I1 (g17028), .I2 (g22285));
NR2X1 gate22599(.O (g24230), .I1 (g17047), .I2 (g22291));
NR2X1 gate22600(.O (g24231), .I1 (g17048), .I2 (g22292));
NR2X1 gate22601(.O (g24232), .I1 (g22637), .I2 (g22665));
NR2X1 gate22602(.O (g24234), .I1 (g22289), .I2 (g21157));
NR2X1 gate22603(.O (g24235), .I1 (g17062), .I2 (g22305));
NR2X1 gate22604(.O (g24237), .I1 (g17081), .I2 (g22311));
NR2X1 gate22605(.O (g24238), .I1 (g17082), .I2 (g22312));
NR2X1 gate22606(.O (g24242), .I1 (g22309), .I2 (g21177));
NR2X1 gate22607(.O (g24243), .I1 (g17097), .I2 (g22333));
NR2X1 gate22608(.O (g24249), .I1 (g22337), .I2 (g21197));
NR2X1 gate22609(.O (g24250), .I1 (g17135), .I2 (g22358));
NR2X1 gate22610(.O (g24426), .I1 (g23386), .I2 (g10024));
NR2X1 gate22611(.O (g24428), .I1 (g23544), .I2 (g22398));
NR2X1 gate22612(.O (g24430), .I1 (g23393), .I2 (g10133));
NR2X1 gate22613(.O (g24434), .I1 (g23401), .I2 (g10238));
NR2X1 gate22614(.O (g24438), .I1 (g23408), .I2 (g10340));
NR2X1 gate22615(.O (g24445), .I1 (g23427), .I2 (g22777));
NR2X1 gate22616(.O (g24446), .I1 (g23433), .I2 (g22907));
NR2X1 gate22617(.O (g24473), .I1 (g23461), .I2 (g18407));
NR2X1 gate22618(.O (g24476), .I1 (g23477), .I2 (g20127));
NR2X1 gate22619(.O (g24479), .I1 (g23593), .I2 (g22516));
NR2X1 gate22620(.O (g24480), .I1 (g23617), .I2 (g23659));
NR2X1 gate22621(.O (g24481), .I1 (g23618), .I2 (g19696));
NR2X1 gate22622(.O (g24485), .I1 (g23625), .I2 (g22556));
NR2X1 gate22623(.O (g24486), .I1 (g23643), .I2 (g22577));
NR2X1 gate22624(.O (g24487), .I1 (g23666), .I2 (g23709));
NR2X1 gate22625(.O (g24488), .I1 (g23667), .I2 (g19740));
NR2X1 gate22626(.O (g24489), .I1 (g23674), .I2 (g22596));
NR2X1 gate22627(.O (g24490), .I1 (g23686), .I2 (g22607));
NR2X1 gate22628(.O (g24491), .I1 (g15247), .I2 (g23735));
NR2X1 gate22629(.O (g24492), .I1 (g23689), .I2 (g22610));
NR2X1 gate22630(.O (g24493), .I1 (g23693), .I2 (g22614));
NR2X1 gate22631(.O (g24494), .I1 (g23716), .I2 (g23763));
NR2X1 gate22632(.O (g24495), .I1 (g23717), .I2 (g19783));
NR2X1 gate22633(.O (g24496), .I1 (g23724), .I2 (g22633));
NR2X1 gate22634(.O (g24497), .I1 (g23734), .I2 (g22638));
NR2X1 gate22635(.O (g24498), .I1 (g15324), .I2 (g23777));
NR2X1 gate22636(.O (g24499), .I1 (g15325), .I2 (g23778));
NR2X1 gate22637(.O (g24500), .I1 (g23740), .I2 (g22643));
NR2X1 gate22638(.O (g24501), .I1 (g15339), .I2 (g23790));
NR2X1 gate22639(.O (g24502), .I1 (g23743), .I2 (g22646));
NR2X1 gate22640(.O (g24503), .I1 (g23747), .I2 (g22650));
NR2X1 gate22641(.O (g24504), .I1 (g23770), .I2 (g23818));
NR2X1 gate22642(.O (g24505), .I1 (g23771), .I2 (g19825));
NR2X1 gate22643(.O (g24506), .I1 (g23776), .I2 (g22667));
NR2X1 gate22644(.O (g24507), .I1 (g15391), .I2 (g23824));
NR2X1 gate22645(.O (g24508), .I1 (g15392), .I2 (g23825));
NR2X1 gate22646(.O (g24509), .I1 (g23789), .I2 (g22674));
NR2X1 gate22647(.O (g24510), .I1 (g15410), .I2 (g23830));
NR2X1 gate22648(.O (g24511), .I1 (g15411), .I2 (g23831));
NR2X1 gate22649(.O (g24512), .I1 (g23795), .I2 (g22679));
NR2X1 gate22650(.O (g24513), .I1 (g15425), .I2 (g23843));
NR2X1 gate22651(.O (g24514), .I1 (g23798), .I2 (g22682));
NR2X1 gate22652(.O (g24515), .I1 (g23802), .I2 (g22686));
NR2X1 gate22653(.O (g24516), .I1 (g23820), .I2 (g22700));
NR2X1 gate22654(.O (g24517), .I1 (g23822), .I2 (g22701));
NR2X1 gate22655(.O (g24519), .I1 (g15459), .I2 (g23855));
NR2X1 gate22656(.O (g24520), .I1 (g23829), .I2 (g22707));
NR2X1 gate22657(.O (g24521), .I1 (g15475), .I2 (g23859));
NR2X1 gate22658(.O (g24522), .I1 (g15476), .I2 (g23860));
NR2X1 gate22659(.O (g24523), .I1 (g23842), .I2 (g22714));
NR2X1 gate22660(.O (g24524), .I1 (g15494), .I2 (g23865));
NR2X1 gate22661(.O (g24525), .I1 (g15495), .I2 (g23866));
NR2X1 gate22662(.O (g24526), .I1 (g23848), .I2 (g22719));
NR2X1 gate22663(.O (g24527), .I1 (g15509), .I2 (g23878));
NR2X1 gate22664(.O (g24528), .I1 (g23851), .I2 (g22722));
NR2X1 gate22665(.O (g24530), .I1 (g23857), .I2 (g22732));
NR2X1 gate22666(.O (g24532), .I1 (g15545), .I2 (g23889));
NR2X1 gate22667(.O (g24533), .I1 (g23864), .I2 (g22738));
NR2X1 gate22668(.O (g24534), .I1 (g15561), .I2 (g23893));
NR2X1 gate22669(.O (g24535), .I1 (g15562), .I2 (g23894));
NR2X1 gate22670(.O (g24536), .I1 (g23877), .I2 (g22745));
NR2X1 gate22671(.O (g24537), .I1 (g15580), .I2 (g23899));
NR2X1 gate22672(.O (g24538), .I1 (g15581), .I2 (g23900));
NR2X1 gate22673(.O (g24543), .I1 (g23891), .I2 (g22764));
NR2X1 gate22674(.O (g24545), .I1 (g15623), .I2 (g23910));
NR2X1 gate22675(.O (g24546), .I1 (g23898), .I2 (g22770));
NR2X1 gate22676(.O (g24547), .I1 (g15639), .I2 (g23914));
NR2X1 gate22677(.O (g24548), .I1 (g15640), .I2 (g23915));
NR2X1 gate22678(.O (g24555), .I1 (g23912), .I2 (g22798));
NR2X1 gate22679(.O (g24557), .I1 (g15699), .I2 (g23942));
NR2X1 gate22680(.O (g24558), .I1 (g23917), .I2 (g22804));
NR2X1 gate22681(.O (g24566), .I1 (g23944), .I2 (g22842));
NR2X1 gate22682(.O (g24575), .I1 (g23972), .I2 (g22874));
NR2X1 gate22683(.O (g24606), .I1 (g24183), .I2 (g537));
NR2X1 gate22684(.O (g24613), .I1 (g23592), .I2 (g22515));
NR2X1 gate22685(.O (g24622), .I1 (g23616), .I2 (g22546));
NR2X1 gate22686(.O (g24623), .I1 (g24183), .I2 (g529));
NR2X1 gate22687(.O (g24624), .I1 (g23624), .I2 (g22555));
NR2X1 gate22688(.O (g24636), .I1 (g24183), .I2 (g530));
NR2X1 gate22689(.O (g24637), .I1 (g23665), .I2 (g22587));
NR2X1 gate22690(.O (g24638), .I1 (g23673), .I2 (g22595));
NR2X1 gate22691(.O (g24652), .I1 (g24183), .I2 (g531));
NR2X1 gate22692(.O (g24656), .I1 (g23715), .I2 (g22624));
NR2X1 gate22693(.O (g24657), .I1 (g23723), .I2 (g22632));
NR2X1 gate22694(.O (g24663), .I1 (g24183), .I2 (g532));
NR2X1 gate22695(.O (g24675), .I1 (g23769), .I2 (g22660));
NR2X1 gate22696(.O (g24681), .I1 (g24183), .I2 (g533));
NR2X1 gate22697(.O (g24682), .I1 (g23688), .I2 (g24183));
NR2X1 gate22698(.O (g24694), .I1 (g24183), .I2 (g534));
NR2X1 gate22699(.O (g24708), .I1 (g23854), .I2 (g22727));
NR2X1 gate22700(.O (g24711), .I1 (g24183), .I2 (g536));
NR2X1 gate22701(.O (g24717), .I1 (g23886), .I2 (g22754));
NR2X1 gate22702(.O (g24720), .I1 (g23888), .I2 (g22759));
NR2X1 gate22703(.O (g24728), .I1 (g23907), .I2 (g22788));
NR2X1 gate22704(.O (g24731), .I1 (g23909), .I2 (g22793));
NR2X1 gate22705(.O (g24736), .I1 (g23939), .I2 (g22830));
NR2X1 gate22706(.O (g24739), .I1 (g23941), .I2 (g22835));
NR2X1 gate22707(.O (g24742), .I1 (g23971), .I2 (g22869));
NR2X1 gate22708(.O (g24756), .I1 (g16089), .I2 (g24211));
NR2X1 gate22709(.O (g24770), .I1 (g16119), .I2 (g24217));
NR2X1 gate22710(.O (g24782), .I1 (g16160), .I2 (g24221));
NR2X1 gate22711(.O (g24783), .I1 (g16161), .I2 (g24224));
NR2X1 gate22712(.O (g24800), .I1 (g16211), .I2 (g24229));
NR2X1 gate22713(.O (g24819), .I1 (g16262), .I2 (g24236));
NR2X1 gate22714(.O (g24836), .I1 (g16309), .I2 (g24241));
NR2X1 gate22715(.O (g24845), .I1 (g16350), .I2 (g24246));
NR2X1 gate22716(.O (g24847), .I1 (g16356), .I2 (g24247));
NR2X1 gate22717(.O (g24859), .I1 (g16390), .I2 (g24253));
NR2X1 gate22718(.O (g24871), .I1 (g16422), .I2 (g24256));
NR2X1 gate22719(.O (g25027), .I1 (g24227), .I2 (g17001));
NR2X1 gate22720(.O (g25042), .I1 (g24234), .I2 (g17031));
NR2X1 gate22721(.O (g25056), .I1 (g24242), .I2 (g17065));
NR2X1 gate22722(.O (g25067), .I1 (g24249), .I2 (g17100));
NR2X1 gate22723(.O (g25075), .I1 (g13880), .I2 (g23483));
NR2X1 gate22724(.O (g25076), .I1 (g23409), .I2 (g22187));
NR2X1 gate22725(.O (g25077), .I1 (g23414), .I2 (g22196));
NR2X1 gate22726(.O (g25078), .I1 (g23419), .I2 (g22201));
NR2X1 gate22727(.O (g25081), .I1 (g23423), .I2 (g22202));
NR2X1 gate22728(.O (g25082), .I1 (g23428), .I2 (g22207));
NR2X1 gate22729(.O (g25085), .I1 (g23432), .I2 (g22208));
NR2X1 gate22730(.O (g25091), .I1 (g23434), .I2 (g22215));
NR2X1 gate22731(.O (g25099), .I1 (g23440), .I2 (g22224));
NR2X1 gate22732(.O (g25125), .I1 (g23510), .I2 (g22340));
NR2X1 gate22733(.O (g25127), .I1 (g23525), .I2 (g22363));
NR2X1 gate22734(.O (g25129), .I1 (g23536), .I2 (g22383));
NR2X1 gate22735(.O (g25185), .I1 (g24492), .I2 (g10024));
NR2X1 gate22736(.O (g25189), .I1 (g24502), .I2 (g10133));
NR2X1 gate22737(.O (g25191), .I1 (g24516), .I2 (g22777));
NR2X1 gate22738(.O (g25194), .I1 (g24514), .I2 (g10238));
NR2X1 gate22739(.O (g25197), .I1 (g24528), .I2 (g10340));
NR2X1 gate22740(.O (g25199), .I1 (g24558), .I2 (g20127));
NR2X1 gate22741(.O (g25201), .I1 (g24575), .I2 (g18407));
NR2X1 gate22742(.O (g25202), .I1 (g24566), .I2 (g22907));
NR2X1 gate22743(.O (g25204), .I1 (g24745), .I2 (g23547));
NR2X1 gate22744(.O (g25206), .I1 (g24746), .I2 (g23550));
NR2X1 gate22745(.O (g25207), .I1 (g24747), .I2 (g23551));
NR2X1 gate22746(.O (g25208), .I1 (g24748), .I2 (g23552));
NR2X1 gate22747(.O (g25209), .I1 (g24749), .I2 (g23554));
NR2X1 gate22748(.O (g25211), .I1 (g24750), .I2 (g23558));
NR2X1 gate22749(.O (g25212), .I1 (g24751), .I2 (g23559));
NR2X1 gate22750(.O (g25213), .I1 (g24752), .I2 (g23560));
NR2X1 gate22751(.O (g25214), .I1 (g24754), .I2 (g23563));
NR2X1 gate22752(.O (g25215), .I1 (g24755), .I2 (g23564));
NR2X1 gate22753(.O (g25216), .I1 (g24757), .I2 (g23565));
NR2X1 gate22754(.O (g25217), .I1 (g24758), .I2 (g23567));
NR2X1 gate22755(.O (g25218), .I1 (g24760), .I2 (g23571));
NR2X1 gate22756(.O (g25219), .I1 (g24761), .I2 (g23572));
NR2X1 gate22757(.O (g25220), .I1 (g24762), .I2 (g23573));
NR2X1 gate22758(.O (g25221), .I1 (g24767), .I2 (g23577));
NR2X1 gate22759(.O (g25222), .I1 (g24768), .I2 (g23578));
NR2X1 gate22760(.O (g25223), .I1 (g24769), .I2 (g23579));
NR2X1 gate22761(.O (g25224), .I1 (g24772), .I2 (g23582));
NR2X1 gate22762(.O (g25225), .I1 (g24773), .I2 (g23583));
NR2X1 gate22763(.O (g25226), .I1 (g24774), .I2 (g23584));
NR2X1 gate22764(.O (g25227), .I1 (g24775), .I2 (g23586));
NR2X1 gate22765(.O (g25228), .I1 (g24776), .I2 (g23590));
NR2X1 gate22766(.O (g25229), .I1 (g24777), .I2 (g23591));
NR2X1 gate22767(.O (g25230), .I1 (g24779), .I2 (g23598));
NR2X1 gate22768(.O (g25231), .I1 (g24780), .I2 (g23599));
NR2X1 gate22769(.O (g25232), .I1 (g24781), .I2 (g23600));
NR2X1 gate22770(.O (g25233), .I1 (g24788), .I2 (g23604));
NR2X1 gate22771(.O (g25234), .I1 (g24789), .I2 (g23605));
NR2X1 gate22772(.O (g25235), .I1 (g24790), .I2 (g23606));
NR2X1 gate22773(.O (g25236), .I1 (g24792), .I2 (g23609));
NR2X1 gate22774(.O (g25237), .I1 (g24793), .I2 (g23610));
NR2X1 gate22775(.O (g25238), .I1 (g24794), .I2 (g23611));
NR2X1 gate22776(.O (g25239), .I1 (g24796), .I2 (g23615));
NR2X1 gate22777(.O (g25240), .I1 (g24798), .I2 (g23622));
NR2X1 gate22778(.O (g25241), .I1 (g24799), .I2 (g23623));
NR2X1 gate22779(.O (g25242), .I1 (g24802), .I2 (g23630));
NR2X1 gate22780(.O (g25243), .I1 (g24803), .I2 (g23631));
NR2X1 gate22781(.O (g25244), .I1 (g24804), .I2 (g23632));
NR2X1 gate22782(.O (g25245), .I1 (g24809), .I2 (g23636));
NR2X1 gate22783(.O (g25246), .I1 (g24810), .I2 (g23637));
NR2X1 gate22784(.O (g25247), .I1 (g24811), .I2 (g23638));
NR2X1 gate22785(.O (g25248), .I1 (g24818), .I2 (g23664));
NR2X1 gate22786(.O (g25249), .I1 (g24821), .I2 (g23671));
NR2X1 gate22787(.O (g25250), .I1 (g24822), .I2 (g23672));
NR2X1 gate22788(.O (g25251), .I1 (g24824), .I2 (g23679));
NR2X1 gate22789(.O (g25252), .I1 (g24825), .I2 (g23680));
NR2X1 gate22790(.O (g25253), .I1 (g24826), .I2 (g23681));
NR2X1 gate22791(.O (g25254), .I1 (g24831), .I2 (g23687));
NR2X1 gate22792(.O (g25255), .I1 (g24838), .I2 (g23714));
NR2X1 gate22793(.O (g25256), .I1 (g24840), .I2 (g23721));
NR2X1 gate22794(.O (g25257), .I1 (g24841), .I2 (g23722));
NR2X1 gate22795(.O (g25258), .I1 (g24846), .I2 (g23741));
NR2X1 gate22796(.O (g25259), .I1 (g24853), .I2 (g23768));
NR2X1 gate22797(.O (g25260), .I1 (g24858), .I2 (g17737));
NR2X1 gate22798(.O (g25261), .I1 (g24861), .I2 (g23796));
NR2X1 gate22799(.O (g25262), .I1 (g24869), .I2 (g17824));
NR2X1 gate22800(.O (g25263), .I1 (g24874), .I2 (g17838));
NR2X1 gate22801(.O (g25264), .I1 (g24876), .I2 (g23849));
NR2X1 gate22802(.O (g25265), .I1 (g24878), .I2 (g23852));
NR2X1 gate22803(.O (g25266), .I1 (g24881), .I2 (g17912));
NR2X1 gate22804(.O (g25267), .I1 (g24884), .I2 (g17936));
NR2X1 gate22805(.O (g25268), .I1 (g24888), .I2 (g17950));
NR2X1 gate22806(.O (g25270), .I1 (g24898), .I2 (g18023));
NR2X1 gate22807(.O (g25271), .I1 (g24901), .I2 (g18047));
NR2X1 gate22808(.O (g25272), .I1 (g24905), .I2 (g18061));
NR2X1 gate22809(.O (g25273), .I1 (g24907), .I2 (g23904));
NR2X1 gate22810(.O (g25279), .I1 (g24921), .I2 (g18140));
NR2X1 gate22811(.O (g25280), .I1 (g24924), .I2 (g18164));
NR2X1 gate22812(.O (g25288), .I1 (g24938), .I2 (g18256));
NR2X1 gate22813(.O (g25311), .I1 (g24964), .I2 (g24029));
NR2X1 gate22814(.O (g25343), .I1 (g24975), .I2 (g5623));
NR2X1 gate22815(.O (g25357), .I1 (g24986), .I2 (g5651));
NR2X1 gate22816(.O (g25372), .I1 (g24997), .I2 (g5689));
NR2X1 gate22817(.O (g25389), .I1 (g25005), .I2 (g5741));
NR2X1 gate22818(.O (g25418), .I1 (g24482), .I2 (g22319));
NR2X1 gate22819(.O (g25426), .I1 (g24183), .I2 (g24616));
NR2X1 gate22820(.O (g25429), .I1 (g24482), .I2 (g22319));
NR2X1 gate22821(.O (g25450), .I1 (g16018), .I2 (g25086));
NR2X1 gate22822(.O (g25451), .I1 (g16048), .I2 (g25102));
NR2X1 gate22823(.O (g25452), .I1 (g16101), .I2 (g25117));
NR2X1 gate22824(.O (g25523), .I1 (g20842), .I2 (g24429));
NR2X1 gate22825(.O (g25539), .I1 (g25088), .I2 (g6157));
NR2X1 gate22826(.O (g25569), .I1 (g24708), .I2 (g24490));
NR2X1 gate22827(.O (g25589), .I1 (g20850), .I2 (g24433));
NR2X1 gate22828(.O (g25605), .I1 (g25096), .I2 (g6184));
NR2X1 gate22829(.O (g25631), .I1 (g24717), .I2 (g24497));
NR2X1 gate22830(.O (g25648), .I1 (g24720), .I2 (g24500));
NR2X1 gate22831(.O (g25668), .I1 (g20858), .I2 (g24437));
NR2X1 gate22832(.O (g25684), .I1 (g25106), .I2 (g6216));
NR2X1 gate22833(.O (g25699), .I1 (g24613), .I2 (g24506));
NR2X1 gate22834(.O (g25708), .I1 (g24728), .I2 (g24509));
NR2X1 gate22835(.O (g25725), .I1 (g24731), .I2 (g24512));
NR2X1 gate22836(.O (g25745), .I1 (g20866), .I2 (g24440));
NR2X1 gate22837(.O (g25761), .I1 (g25112), .I2 (g6305));
NR2X1 gate22838(.O (g25764), .I1 (g25076), .I2 (g21615));
NR2X1 gate22839(.O (g25772), .I1 (g24624), .I2 (g24520));
NR2X1 gate22840(.O (g25781), .I1 (g24736), .I2 (g24523));
NR2X1 gate22841(.O (g25798), .I1 (g24739), .I2 (g24526));
NR2X1 gate22842(.O (g25818), .I1 (g25077), .I2 (g21643));
NR2X1 gate22843(.O (g25826), .I1 (g24638), .I2 (g24533));
NR2X1 gate22844(.O (g25835), .I1 (g24742), .I2 (g24536));
NR3X1 gate22845(.O (g25852), .I1 (g4456), .I2 (g14831), .I3 (g25078));
NR2X1 gate22846(.O (g25853), .I1 (g25081), .I2 (g21674));
NR2X1 gate22847(.O (g25861), .I1 (g24657), .I2 (g24546));
NR4X1 gate22848(.O (g25870), .I1 (g4456), .I2 (g25078), .I3 (g18429), .I4 (g16075));
NR3X1 gate22849(.O (g25873), .I1 (g4632), .I2 (g14904), .I3 (g25082));
NR2X1 gate22850(.O (g25874), .I1 (g25085), .I2 (g21703));
NR4X1 gate22851(.O (g25882), .I1 (g4632), .I2 (g25082), .I3 (g18502), .I4 (g16113));
NR3X1 gate22852(.O (g25885), .I1 (g4809), .I2 (g14985), .I3 (g25091));
NR4X1 gate22853(.O (g25887), .I1 (g4809), .I2 (g25091), .I3 (g18566), .I4 (g16164));
NR3X1 gate22854(.O (g25890), .I1 (g4985), .I2 (g15074), .I3 (g25099));
NR4X1 gate22855(.O (g25892), .I1 (g4985), .I2 (g25099), .I3 (g18616), .I4 (g16223));
NR2X1 gate22856(.O (g25932), .I1 (g25125), .I2 (g17001));
NR2X1 gate22857(.O (g25935), .I1 (g25127), .I2 (g17031));
NR2X1 gate22858(.O (g25938), .I1 (g25129), .I2 (g17065));
NR2X1 gate22859(.O (g25940), .I1 (g24428), .I2 (g17100));
NR2X1 gate22860(.O (g25941), .I1 (g24529), .I2 (g24540));
NR2X1 gate22861(.O (g25943), .I1 (g24541), .I2 (g24550));
NR2X1 gate22862(.O (g25944), .I1 (g24542), .I2 (g24552));
NR2X1 gate22863(.O (g25946), .I1 (g24553), .I2 (g24561));
NR2X1 gate22864(.O (g25947), .I1 (g24554), .I2 (g24563));
NR2X1 gate22865(.O (g25948), .I1 (g24564), .I2 (g24571));
NR2X1 gate22866(.O (g25949), .I1 (g24565), .I2 (g24573));
NR2X1 gate22867(.O (g25950), .I1 (g24574), .I2 (g24580));
NR2X1 gate22868(.O (g25962), .I1 (g24591), .I2 (g23496));
NR2X1 gate22869(.O (g25967), .I1 (g24596), .I2 (g23512));
NR2X1 gate22870(.O (g25974), .I1 (g24604), .I2 (g23527));
NR2X1 gate22871(.O (g25979), .I1 (g24611), .I2 (g23538));
NR2X1 gate22872(.O (g26025), .I1 (g25392), .I2 (g17193));
NR2X1 gate22873(.O (g26031), .I1 (g25273), .I2 (g22777));
NR2X1 gate22874(.O (g26037), .I1 (g25311), .I2 (g18407));
NR2X1 gate22875(.O (g26041), .I1 (g25475), .I2 (g24855));
NR2X1 gate22876(.O (g26042), .I1 (g25505), .I2 (g24867));
NR2X1 gate22877(.O (g26043), .I1 (g25506), .I2 (g24870));
NR2X1 gate22878(.O (g26044), .I1 (g25552), .I2 (g24882));
NR2X1 gate22879(.O (g26045), .I1 (g25553), .I2 (g24885));
NR2X1 gate22880(.O (g26046), .I1 (g25618), .I2 (g24899));
NR2X1 gate22881(.O (g26047), .I1 (g25619), .I2 (g24902));
NR2X1 gate22882(.O (g26048), .I1 (g25628), .I2 (g24906));
NR2X1 gate22883(.O (g26049), .I1 (g25629), .I2 (g24908));
NR2X1 gate22884(.O (g26050), .I1 (g25697), .I2 (g24922));
NR2X1 gate22885(.O (g26055), .I1 (g25881), .I2 (g24974));
NR2X1 gate22886(.O (g26081), .I1 (g25470), .I2 (g25482));
NR2X1 gate22887(.O (g26083), .I1 (g25426), .I2 (g22319));
NR2X1 gate22888(.O (g26084), .I1 (g25487), .I2 (g25513));
NR3X1 gate22889(.O (g26087), .I1 (g6068), .I2 (g24183), .I3 (g25319));
NR2X1 gate22890(.O (g26090), .I1 (g25518), .I2 (g25560));
NR3X1 gate22891(.O (g26096), .I1 (g6068), .I2 (g24183), .I3 (g25394));
NR3X1 gate22892(.O (g26099), .I1 (g6068), .I2 (g24183), .I3 (g25313));
NR2X1 gate22893(.O (g26103), .I1 (g25565), .I2 (g25626));
NR3X1 gate22894(.O (g26107), .I1 (g6068), .I2 (g24183), .I3 (g25383));
NR3X1 gate22895(.O (g26110), .I1 (g6068), .I2 (g24183), .I3 (g25305));
NR2X1 gate22896(.O (g26113), .I1 (g25426), .I2 (g22319));
NR3X1 gate22897(.O (g26126), .I1 (g6068), .I2 (g24183), .I3 (g25368));
NR3X1 gate22898(.O (g26137), .I1 (g6068), .I2 (g24183), .I3 (g25355));
NR2X1 gate22899(.O (g26140), .I1 (g24183), .I2 (g25430));
NR3X1 gate22900(.O (g26145), .I1 (g6068), .I2 (g24183), .I3 (g25347));
NR3X1 gate22901(.O (g26151), .I1 (g6068), .I2 (g24183), .I3 (g25335));
NR3X1 gate22902(.O (g26154), .I1 (g6068), .I2 (g24183), .I3 (g25329));
NR2X1 gate22903(.O (g26160), .I1 (g25951), .I2 (g16162));
NR2X1 gate22904(.O (g26168), .I1 (g25953), .I2 (g16212));
NR2X1 gate22905(.O (g26183), .I1 (g25957), .I2 (g13270));
NR2X1 gate22906(.O (g26199), .I1 (g25961), .I2 (g13291));
NR2X1 gate22907(.O (g26217), .I1 (g25963), .I2 (g13320));
NR2X1 gate22908(.O (g26240), .I1 (g25968), .I2 (g13340));
NR2X1 gate22909(.O (g26265), .I1 (g25972), .I2 (g13360));
NR2X1 gate22910(.O (g26272), .I1 (g25973), .I2 (g16423));
NR2X1 gate22911(.O (g26283), .I1 (g25954), .I2 (g24486));
NR2X1 gate22912(.O (g26295), .I1 (g25977), .I2 (g13385));
NR2X1 gate22913(.O (g26304), .I1 (g25978), .I2 (g16451));
NR2X1 gate22914(.O (g26327), .I1 (g25958), .I2 (g24493));
NR2X1 gate22915(.O (g26336), .I1 (g25981), .I2 (g13481));
NR2X1 gate22916(.O (g26374), .I1 (g25964), .I2 (g24503));
NR2X1 gate22917(.O (g26417), .I1 (g25969), .I2 (g24515));
NR2X1 gate22918(.O (g26529), .I1 (g25962), .I2 (g17001));
NR2X1 gate22919(.O (g26530), .I1 (g25967), .I2 (g17031));
NR2X1 gate22920(.O (g26531), .I1 (g25974), .I2 (g17065));
NR2X1 gate22921(.O (g26532), .I1 (g25979), .I2 (g17100));
NR2X1 gate22922(.O (g26534), .I1 (g25321), .I2 (g8869));
NR2X1 gate22923(.O (g26541), .I1 (g13755), .I2 (g25269));
NR2X1 gate22924(.O (g26545), .I1 (g13790), .I2 (g25277));
NR2X1 gate22925(.O (g26547), .I1 (g13796), .I2 (g25278));
NR2X1 gate22926(.O (g26553), .I1 (g13816), .I2 (g25282));
NR2X1 gate22927(.O (g26557), .I1 (g13818), .I2 (g25286));
NR2X1 gate22928(.O (g26559), .I1 (g13824), .I2 (g25287));
NR2X1 gate22929(.O (g26560), .I1 (g25281), .I2 (g24559));
NR2X1 gate22930(.O (g26569), .I1 (g13837), .I2 (g25290));
NR2X1 gate22931(.O (g26573), .I1 (g13839), .I2 (g25294));
NR2X1 gate22932(.O (g26575), .I1 (g13845), .I2 (g25295));
NR2X1 gate22933(.O (g26583), .I1 (g25289), .I2 (g24569));
NR2X1 gate22934(.O (g26592), .I1 (g13851), .I2 (g25300));
NR2X1 gate22935(.O (g26596), .I1 (g13853), .I2 (g25304));
NR2X1 gate22936(.O (g26607), .I1 (g25299), .I2 (g24578));
NR2X1 gate22937(.O (g26616), .I1 (g13860), .I2 (g25310));
NR2X1 gate22938(.O (g26630), .I1 (g25309), .I2 (g24585));
NR2X1 gate22939(.O (g26655), .I1 (g25328), .I2 (g17084));
NR2X1 gate22940(.O (g26659), .I1 (g25334), .I2 (g17116));
NR2X1 gate22941(.O (g26660), .I1 (g25208), .I2 (g10024));
NR2X1 gate22942(.O (g26661), .I1 (g25337), .I2 (g17122));
NR2X1 gate22943(.O (g26664), .I1 (g25346), .I2 (g17138));
NR2X1 gate22944(.O (g26665), .I1 (g25348), .I2 (g17143));
NR2X1 gate22945(.O (g26666), .I1 (g25216), .I2 (g10133));
NR2X1 gate22946(.O (g26667), .I1 (g25351), .I2 (g17149));
NR2X1 gate22947(.O (g26669), .I1 (g25360), .I2 (g17161));
NR2X1 gate22948(.O (g26670), .I1 (g25362), .I2 (g17166));
NR2X1 gate22949(.O (g26671), .I1 (g25226), .I2 (g10238));
NR2X1 gate22950(.O (g26672), .I1 (g25365), .I2 (g17172));
NR2X1 gate22951(.O (g26675), .I1 (g25375), .I2 (g17176));
NR2X1 gate22952(.O (g26676), .I1 (g25377), .I2 (g17181));
NR2X1 gate22953(.O (g26677), .I1 (g25238), .I2 (g10340));
NR2X1 gate22954(.O (g26776), .I1 (g26042), .I2 (g10024));
NR2X1 gate22955(.O (g26781), .I1 (g26044), .I2 (g10133));
NR2X1 gate22956(.O (g26786), .I1 (g26049), .I2 (g22777));
NR2X1 gate22957(.O (g26789), .I1 (g26046), .I2 (g10238));
NR2X1 gate22958(.O (g26795), .I1 (g26050), .I2 (g10340));
NR2X1 gate22959(.O (g26798), .I1 (g26055), .I2 (g18407));
NR2X1 gate22960(.O (g26799), .I1 (g26158), .I2 (g25453));
NR2X1 gate22961(.O (g26800), .I1 (g26163), .I2 (g25457));
NR2X1 gate22962(.O (g26801), .I1 (g26171), .I2 (g25461));
NR2X1 gate22963(.O (g26802), .I1 (g26188), .I2 (g25466));
NR2X1 gate22964(.O (g26803), .I1 (g15105), .I2 (g26213));
NR2X1 gate22965(.O (g26804), .I1 (g15172), .I2 (g26235));
NR2X1 gate22966(.O (g26805), .I1 (g15173), .I2 (g26236));
NR2X1 gate22967(.O (g26806), .I1 (g15197), .I2 (g26244));
NR2X1 gate22968(.O (g26807), .I1 (g15245), .I2 (g26261));
NR2X1 gate22969(.O (g26808), .I1 (g15246), .I2 (g26262));
NR2X1 gate22970(.O (g26809), .I1 (g15258), .I2 (g26270));
NR2X1 gate22971(.O (g26810), .I1 (g15259), .I2 (g26271));
NR2X1 gate22972(.O (g26811), .I1 (g15283), .I2 (g26279));
NR2X1 gate22973(.O (g26812), .I1 (g15321), .I2 (g26291));
NR2X1 gate22974(.O (g26813), .I1 (g15337), .I2 (g26302));
NR2X1 gate22975(.O (g26814), .I1 (g15338), .I2 (g26303));
NR2X1 gate22976(.O (g26815), .I1 (g15350), .I2 (g26311));
NR2X1 gate22977(.O (g26816), .I1 (g15351), .I2 (g26312));
NR2X1 gate22978(.O (g26817), .I1 (g15375), .I2 (g26317));
NR2X1 gate22979(.O (g26818), .I1 (g15407), .I2 (g26335));
NR2X1 gate22980(.O (g26820), .I1 (g15423), .I2 (g26346));
NR2X1 gate22981(.O (g26821), .I1 (g15424), .I2 (g26347));
NR2X1 gate22982(.O (g26822), .I1 (g15436), .I2 (g26352));
NR2X1 gate22983(.O (g26823), .I1 (g15437), .I2 (g26353));
NR2X1 gate22984(.O (g26824), .I1 (g15491), .I2 (g26382));
NR2X1 gate22985(.O (g26825), .I1 (g15507), .I2 (g26390));
NR2X1 gate22986(.O (g26826), .I1 (g15508), .I2 (g26391));
NR2X1 gate22987(.O (g26827), .I1 (g15577), .I2 (g26425));
NR2X1 gate22988(.O (g26869), .I1 (g26458), .I2 (g5642));
NR2X1 gate22989(.O (g26873), .I1 (g25483), .I2 (g26260));
NR2X1 gate22990(.O (g26877), .I1 (g26140), .I2 (g22319));
NR2X1 gate22991(.O (g26878), .I1 (g26482), .I2 (g5680));
NR2X1 gate22992(.O (g26882), .I1 (g25514), .I2 (g26301));
NR2X1 gate22993(.O (g26885), .I1 (g26140), .I2 (g22319));
NR2X1 gate22994(.O (g26887), .I1 (g26498), .I2 (g5732));
NR2X1 gate22995(.O (g26891), .I1 (g25561), .I2 (g26345));
NR2X1 gate22996(.O (g26897), .I1 (g26513), .I2 (g5790));
NR2X1 gate22997(.O (g26901), .I1 (g25627), .I2 (g26389));
NR2X1 gate22998(.O (g26905), .I1 (g26096), .I2 (g22319));
NR2X1 gate22999(.O (g26914), .I1 (g26107), .I2 (g22319));
NR2X1 gate23000(.O (g26988), .I1 (g24893), .I2 (g26023));
NR2X1 gate23001(.O (g26989), .I1 (g26663), .I2 (g21913));
NR2X1 gate23002(.O (g27011), .I1 (g24916), .I2 (g26026));
NR2X1 gate23003(.O (g27012), .I1 (g26668), .I2 (g21931));
NR2X1 gate23004(.O (g27037), .I1 (g24933), .I2 (g26028));
NR2X1 gate23005(.O (g27038), .I1 (g26674), .I2 (g20640));
NR2X1 gate23006(.O (g27051), .I1 (g4456), .I2 (g26081));
NR2X1 gate23007(.O (g27065), .I1 (g24945), .I2 (g26029));
NR2X1 gate23008(.O (g27066), .I1 (g26024), .I2 (g20665));
NR2X1 gate23009(.O (g27078), .I1 (g4632), .I2 (g26084));
NR2X1 gate23010(.O (g27094), .I1 (g4809), .I2 (g26090));
NR2X1 gate23011(.O (g27106), .I1 (g4985), .I2 (g26103));
NR2X1 gate23012(.O (g27120), .I1 (g26560), .I2 (g17001));
NR2X1 gate23013(.O (g27123), .I1 (g26583), .I2 (g17031));
NR2X1 gate23014(.O (g27129), .I1 (g26607), .I2 (g17065));
NR2X1 gate23015(.O (g27131), .I1 (g26630), .I2 (g17100));
NR2X1 gate23016(.O (g27144), .I1 (g23451), .I2 (g26052));
NR2X1 gate23017(.O (g27147), .I1 (g23458), .I2 (g26054));
NR2X1 gate23018(.O (g27149), .I1 (g23462), .I2 (g26060));
NR2X1 gate23019(.O (g27152), .I1 (g23467), .I2 (g26062));
NR2X1 gate23020(.O (g27157), .I1 (g23471), .I2 (g26067));
NR2X1 gate23021(.O (g27160), .I1 (g23476), .I2 (g26069));
NR2X1 gate23022(.O (g27165), .I1 (g23484), .I2 (g26074));
NR2X1 gate23023(.O (g27174), .I1 (g23494), .I2 (g26080));
NR2X1 gate23024(.O (g27175), .I1 (g26075), .I2 (g25342));
NR2X1 gate23025(.O (g27179), .I1 (g26082), .I2 (g25356));
NR2X1 gate23026(.O (g27184), .I1 (g26085), .I2 (g25371));
NR2X1 gate23027(.O (g27188), .I1 (g26091), .I2 (g25388));
NR2X1 gate23028(.O (g27243), .I1 (g26802), .I2 (g10340));
NR2X1 gate23029(.O (g27250), .I1 (g26955), .I2 (g26166));
NR2X1 gate23030(.O (g27251), .I1 (g26958), .I2 (g26186));
NR2X1 gate23031(.O (g27252), .I1 (g26963), .I2 (g26207));
NR2X1 gate23032(.O (g27253), .I1 (g26965), .I2 (g26212));
NR2X1 gate23033(.O (g27254), .I1 (g26968), .I2 (g26231));
NR2X1 gate23034(.O (g27255), .I1 (g26969), .I2 (g26233));
NR2X1 gate23035(.O (g27256), .I1 (g26970), .I2 (g26234));
NR2X1 gate23036(.O (g27257), .I1 (g26971), .I2 (g26243));
NR2X1 gate23037(.O (g27258), .I1 (g26977), .I2 (g26257));
NR2X1 gate23038(.O (g27259), .I1 (g26978), .I2 (g26258));
NR2X1 gate23039(.O (g27260), .I1 (g26979), .I2 (g26259));
NR2X1 gate23040(.O (g27261), .I1 (g26980), .I2 (g26263));
NR2X1 gate23041(.O (g27262), .I1 (g26981), .I2 (g26268));
NR2X1 gate23042(.O (g27263), .I1 (g26982), .I2 (g26269));
NR2X1 gate23043(.O (g27264), .I1 (g26984), .I2 (g26278));
NR2X1 gate23044(.O (g27265), .I1 (g26993), .I2 (g26288));
NR2X1 gate23045(.O (g27266), .I1 (g26994), .I2 (g26289));
NR2X1 gate23046(.O (g27267), .I1 (g26995), .I2 (g26290));
NR2X1 gate23047(.O (g27268), .I1 (g26996), .I2 (g26292));
NR2X1 gate23048(.O (g27269), .I1 (g26997), .I2 (g26293));
NR2X1 gate23049(.O (g27270), .I1 (g26998), .I2 (g26298));
NR2X1 gate23050(.O (g27271), .I1 (g26999), .I2 (g26299));
NR2X1 gate23051(.O (g27272), .I1 (g27000), .I2 (g26300));
NR2X1 gate23052(.O (g27273), .I1 (g27001), .I2 (g26307));
NR2X1 gate23053(.O (g27274), .I1 (g27002), .I2 (g26309));
NR2X1 gate23054(.O (g27275), .I1 (g27003), .I2 (g26310));
NR2X1 gate23055(.O (g27276), .I1 (g27004), .I2 (g26316));
NR2X1 gate23056(.O (g27277), .I1 (g27005), .I2 (g26318));
NR2X1 gate23057(.O (g27278), .I1 (g27006), .I2 (g26319));
NR2X1 gate23058(.O (g27279), .I1 (g27007), .I2 (g26324));
NR2X1 gate23059(.O (g27280), .I1 (g27008), .I2 (g26325));
NR2X1 gate23060(.O (g27281), .I1 (g27009), .I2 (g26326));
NR2X1 gate23061(.O (g27282), .I1 (g27016), .I2 (g26332));
NR2X1 gate23062(.O (g27283), .I1 (g27017), .I2 (g26333));
NR2X1 gate23063(.O (g27284), .I1 (g27018), .I2 (g26334));
NR2X1 gate23064(.O (g27285), .I1 (g27019), .I2 (g26339));
NR2X1 gate23065(.O (g27286), .I1 (g27020), .I2 (g26340));
NR2X1 gate23066(.O (g27287), .I1 (g27021), .I2 (g26342));
NR2X1 gate23067(.O (g27288), .I1 (g27022), .I2 (g26343));
NR2X1 gate23068(.O (g27289), .I1 (g27023), .I2 (g26344));
NR2X1 gate23069(.O (g27290), .I1 (g27024), .I2 (g26348));
NR2X1 gate23070(.O (g27291), .I1 (g27025), .I2 (g26350));
NR2X1 gate23071(.O (g27292), .I1 (g27026), .I2 (g26351));
NR2X1 gate23072(.O (g27293), .I1 (g27027), .I2 (g26357));
NR2X1 gate23073(.O (g27294), .I1 (g27028), .I2 (g26361));
NR2X1 gate23074(.O (g27295), .I1 (g27029), .I2 (g26362));
NR2X1 gate23075(.O (g27296), .I1 (g27030), .I2 (g26363));
NR2X1 gate23076(.O (g27297), .I1 (g27031), .I2 (g26365));
NR2X1 gate23077(.O (g27298), .I1 (g27032), .I2 (g26366));
NR2X1 gate23078(.O (g27299), .I1 (g27033), .I2 (g26371));
NR2X1 gate23079(.O (g27300), .I1 (g27034), .I2 (g26372));
NR2X1 gate23080(.O (g27301), .I1 (g27035), .I2 (g26373));
NR2X1 gate23081(.O (g27302), .I1 (g27042), .I2 (g26379));
NR2X1 gate23082(.O (g27303), .I1 (g27043), .I2 (g26380));
NR2X1 gate23083(.O (g27304), .I1 (g27044), .I2 (g26381));
NR2X1 gate23084(.O (g27305), .I1 (g27045), .I2 (g26383));
NR2X1 gate23085(.O (g27306), .I1 (g27046), .I2 (g26384));
NR2X1 gate23086(.O (g27307), .I1 (g27047), .I2 (g26386));
NR2X1 gate23087(.O (g27308), .I1 (g27048), .I2 (g26387));
NR2X1 gate23088(.O (g27309), .I1 (g27049), .I2 (g26388));
NR2X1 gate23089(.O (g27310), .I1 (g27050), .I2 (g26392));
NR2X1 gate23090(.O (g27311), .I1 (g27053), .I2 (g26396));
NR2X1 gate23091(.O (g27312), .I1 (g27054), .I2 (g26397));
NR2X1 gate23092(.O (g27313), .I1 (g27055), .I2 (g26400));
NR2X1 gate23093(.O (g27314), .I1 (g27056), .I2 (g26404));
NR2X1 gate23094(.O (g27315), .I1 (g27057), .I2 (g26405));
NR2X1 gate23095(.O (g27316), .I1 (g27058), .I2 (g26406));
NR2X1 gate23096(.O (g27317), .I1 (g27059), .I2 (g26408));
NR2X1 gate23097(.O (g27318), .I1 (g27060), .I2 (g26409));
NR2X1 gate23098(.O (g27319), .I1 (g27061), .I2 (g26414));
NR2X1 gate23099(.O (g27320), .I1 (g27062), .I2 (g26415));
NR2X1 gate23100(.O (g27321), .I1 (g27063), .I2 (g26416));
NR2X1 gate23101(.O (g27322), .I1 (g27070), .I2 (g26422));
NR2X1 gate23102(.O (g27323), .I1 (g27071), .I2 (g26423));
NR2X1 gate23103(.O (g27324), .I1 (g27072), .I2 (g26424));
NR2X1 gate23104(.O (g27325), .I1 (g27073), .I2 (g26426));
NR2X1 gate23105(.O (g27326), .I1 (g27074), .I2 (g26427));
NR2X1 gate23106(.O (g27327), .I1 (g27077), .I2 (g26432));
NR2X1 gate23107(.O (g27328), .I1 (g27080), .I2 (g26437));
NR2X1 gate23108(.O (g27329), .I1 (g27081), .I2 (g26438));
NR2X1 gate23109(.O (g27330), .I1 (g27082), .I2 (g26441));
NR2X1 gate23110(.O (g27331), .I1 (g27083), .I2 (g26445));
NR2X1 gate23111(.O (g27332), .I1 (g27084), .I2 (g26446));
NR2X1 gate23112(.O (g27333), .I1 (g27085), .I2 (g26447));
NR2X1 gate23113(.O (g27334), .I1 (g27086), .I2 (g26449));
NR2X1 gate23114(.O (g27335), .I1 (g27087), .I2 (g26450));
NR2X1 gate23115(.O (g27336), .I1 (g27088), .I2 (g26455));
NR2X1 gate23116(.O (g27337), .I1 (g27089), .I2 (g26456));
NR2X1 gate23117(.O (g27338), .I1 (g27090), .I2 (g26457));
NR2X1 gate23118(.O (g27339), .I1 (g27093), .I2 (g26464));
NR2X1 gate23119(.O (g27340), .I1 (g27096), .I2 (g26469));
NR2X1 gate23120(.O (g27341), .I1 (g27097), .I2 (g26470));
NR2X1 gate23121(.O (g27342), .I1 (g27098), .I2 (g26473));
NR2X1 gate23122(.O (g27343), .I1 (g27099), .I2 (g26477));
NR2X1 gate23123(.O (g27344), .I1 (g27100), .I2 (g26478));
NR2X1 gate23124(.O (g27345), .I1 (g27101), .I2 (g26479));
NR2X1 gate23125(.O (g27346), .I1 (g27105), .I2 (g26488));
NR2X1 gate23126(.O (g27347), .I1 (g27108), .I2 (g26493));
NR2X1 gate23127(.O (g27348), .I1 (g27109), .I2 (g26494));
NR2X1 gate23128(.O (g27354), .I1 (g27112), .I2 (g26504));
NR2X1 gate23129(.O (g27414), .I1 (g26770), .I2 (g25187));
NR3X1 gate23130(.O (g27415), .I1 (g23104), .I2 (g27181), .I3 (g25128));
NR2X1 gate23131(.O (g27435), .I1 (g26777), .I2 (g25193));
NR3X1 gate23132(.O (g27436), .I1 (g23118), .I2 (g27187), .I3 (g24427));
NR2X1 gate23133(.O (g27450), .I1 (g26902), .I2 (g24613));
NR2X1 gate23134(.O (g27454), .I1 (g26783), .I2 (g25196));
NR3X1 gate23135(.O (g27455), .I1 (g23127), .I2 (g26758), .I3 (g24431));
NR2X1 gate23136(.O (g27462), .I1 (g26892), .I2 (g24622));
NR2X1 gate23137(.O (g27464), .I1 (g27178), .I2 (g25975));
NR2X1 gate23138(.O (g27466), .I1 (g26915), .I2 (g24624));
NR2X1 gate23139(.O (g27470), .I1 (g26790), .I2 (g25198));
NR3X1 gate23140(.O (g27471), .I1 (g23138), .I2 (g26764), .I3 (g24435));
NR2X1 gate23141(.O (g27478), .I1 (g26754), .I2 (g24432));
NR2X1 gate23142(.O (g27481), .I1 (g27182), .I2 (g25980));
NR2X1 gate23143(.O (g27482), .I1 (g26906), .I2 (g24637));
NR2X1 gate23144(.O (g27485), .I1 (g26928), .I2 (g24638));
NR3X1 gate23145(.O (g27492), .I1 (g24958), .I2 (g24633), .I3 (g26771));
NR2X1 gate23146(.O (g27496), .I1 (g27185), .I2 (g25178));
NR2X1 gate23147(.O (g27501), .I1 (g26763), .I2 (g24436));
NR2X1 gate23148(.O (g27504), .I1 (g26918), .I2 (g24656));
NR2X1 gate23149(.O (g27507), .I1 (g26941), .I2 (g24657));
NR3X1 gate23150(.O (g27513), .I1 (g24969), .I2 (g24653), .I3 (g26778));
NR2X1 gate23151(.O (g27521), .I1 (g26766), .I2 (g24439));
NR2X1 gate23152(.O (g27524), .I1 (g26931), .I2 (g24675));
NR2X1 gate23153(.O (g27527), .I1 (g26759), .I2 (g19087));
NR2X1 gate23154(.O (g27529), .I1 (g4456), .I2 (g26873));
NR2X1 gate23155(.O (g27531), .I1 (g26760), .I2 (g25181));
NR2X1 gate23156(.O (g27532), .I1 (g26761), .I2 (g25182));
NR3X1 gate23157(.O (g27538), .I1 (g24982), .I2 (g24672), .I3 (g26784));
NR2X1 gate23158(.O (g27546), .I1 (g26769), .I2 (g24441));
NR2X1 gate23159(.O (g27549), .I1 (g26765), .I2 (g19093));
NR2X1 gate23160(.O (g27551), .I1 (g4632), .I2 (g26882));
NR3X1 gate23161(.O (g27558), .I1 (g24993), .I2 (g24691), .I3 (g26791));
NR2X1 gate23162(.O (g27563), .I1 (g26922), .I2 (g24708));
NR2X1 gate23163(.O (g27564), .I1 (g26767), .I2 (g25184));
NR2X1 gate23164(.O (g27565), .I1 (g26768), .I2 (g19100));
NR2X1 gate23165(.O (g27567), .I1 (g4809), .I2 (g26891));
NR2X1 gate23166(.O (g27572), .I1 (g26911), .I2 (g24717));
NR2X1 gate23167(.O (g27573), .I1 (g26773), .I2 (g25188));
NR2X1 gate23168(.O (g27574), .I1 (g26935), .I2 (g24720));
NR2X1 gate23169(.O (g27575), .I1 (g26774), .I2 (g19107));
NR2X1 gate23170(.O (g27577), .I1 (g4985), .I2 (g26901));
NR2X1 gate23171(.O (g27579), .I1 (g26775), .I2 (g25192));
NR2X1 gate23172(.O (g27581), .I1 (g26925), .I2 (g24728));
NR2X1 gate23173(.O (g27582), .I1 (g26944), .I2 (g24731));
NR2X1 gate23174(.O (g27584), .I1 (g26938), .I2 (g24736));
NR2X1 gate23175(.O (g27585), .I1 (g26950), .I2 (g24739));
NR2X1 gate23176(.O (g27588), .I1 (g26947), .I2 (g24742));
NR2X1 gate23177(.O (g27594), .I1 (g27175), .I2 (g17001));
NR2X1 gate23178(.O (g27603), .I1 (g27179), .I2 (g17031));
NR2X1 gate23179(.O (g27612), .I1 (g27184), .I2 (g17065));
NR2X1 gate23180(.O (g27621), .I1 (g27188), .I2 (g17100));
NR2X1 gate23181(.O (g27629), .I1 (g26829), .I2 (g26051));
NR2X1 gate23182(.O (g27631), .I1 (g26833), .I2 (g26053));
NR2X1 gate23183(.O (g27655), .I1 (g26842), .I2 (g26061));
NR2X1 gate23184(.O (g27658), .I1 (g26851), .I2 (g26068));
NR2X1 gate23185(.O (g27672), .I1 (g26799), .I2 (g10024));
NR2X1 gate23186(.O (g27678), .I1 (g26800), .I2 (g10133));
NR2X1 gate23187(.O (g27682), .I1 (g26801), .I2 (g10238));
NR2X1 gate23188(.O (g27718), .I1 (g27251), .I2 (g10133));
NR2X1 gate23189(.O (g27722), .I1 (g27252), .I2 (g10238));
NR2X1 gate23190(.O (g27724), .I1 (g27254), .I2 (g10340));
NR2X1 gate23191(.O (g27735), .I1 (g27394), .I2 (g26961));
NR2X1 gate23192(.O (g27736), .I1 (g27396), .I2 (g26962));
NR2X1 gate23193(.O (g27741), .I1 (g27407), .I2 (g26966));
NR2X1 gate23194(.O (g27742), .I1 (g27409), .I2 (g26967));
NR2X1 gate23195(.O (g27746), .I1 (g27425), .I2 (g26972));
NR2X1 gate23196(.O (g27747), .I1 (g27427), .I2 (g26973));
NR2X1 gate23197(.O (g27754), .I1 (g27446), .I2 (g26985));
NR2X1 gate23198(.O (g27755), .I1 (g27448), .I2 (g26986));
NR2X1 gate23199(.O (g27759), .I1 (g27495), .I2 (g27052));
NR2X1 gate23200(.O (g27760), .I1 (g27509), .I2 (g27076));
NR2X1 gate23201(.O (g27761), .I1 (g27516), .I2 (g27079));
NR2X1 gate23202(.O (g27762), .I1 (g27530), .I2 (g27091));
NR2X1 gate23203(.O (g27763), .I1 (g27534), .I2 (g27092));
NR2X1 gate23204(.O (g27764), .I1 (g27541), .I2 (g27095));
NR2X1 gate23205(.O (g27765), .I1 (g27552), .I2 (g27103));
NR2X1 gate23206(.O (g27766), .I1 (g27554), .I2 (g27104));
NR2X1 gate23207(.O (g27767), .I1 (g27561), .I2 (g27107));
NR2X1 gate23208(.O (g27768), .I1 (g27568), .I2 (g27110));
NR2X1 gate23209(.O (g27769), .I1 (g27570), .I2 (g27111));
NR2X1 gate23210(.O (g27771), .I1 (g27578), .I2 (g27115));
NR2X1 gate23211(.O (g27798), .I1 (g27632), .I2 (g1223));
NR3X1 gate23212(.O (g27802), .I1 (g6087), .I2 (g27632), .I3 (g25330));
NR2X1 gate23213(.O (g27810), .I1 (g27632), .I2 (g1215));
NR3X1 gate23214(.O (g27811), .I1 (g6087), .I2 (g27632), .I3 (g25404));
NR3X1 gate23215(.O (g27814), .I1 (g6087), .I2 (g27632), .I3 (g25322));
NR2X1 gate23216(.O (g27823), .I1 (g27632), .I2 (g1216));
NR3X1 gate23217(.O (g27824), .I1 (g6087), .I2 (g27632), .I3 (g25399));
NR3X1 gate23218(.O (g27827), .I1 (g6087), .I2 (g27632), .I3 (g25314));
NR2X1 gate23219(.O (g27834), .I1 (g27478), .I2 (g14630));
NR2X1 gate23220(.O (g27842), .I1 (g27632), .I2 (g1217));
NR2X1 gate23221(.O (g27850), .I1 (g27501), .I2 (g14650));
NR2X1 gate23222(.O (g27854), .I1 (g27632), .I2 (g1218));
NR3X1 gate23223(.O (g27855), .I1 (g6087), .I2 (g27632), .I3 (g25385));
NR2X1 gate23224(.O (g27864), .I1 (g27632), .I2 (g1219));
NR3X1 gate23225(.O (g27865), .I1 (g6087), .I2 (g27632), .I3 (g25370));
NR2X1 gate23226(.O (g27868), .I1 (g23742), .I2 (g27632));
NR2X1 gate23227(.O (g27869), .I1 (g27632), .I2 (g25437));
NR2X1 gate23228(.O (g27875), .I1 (g27521), .I2 (g14677));
NR2X1 gate23229(.O (g27882), .I1 (g27632), .I2 (g1220));
NR3X1 gate23230(.O (g27883), .I1 (g6087), .I2 (g27632), .I3 (g25361));
NR2X1 gate23231(.O (g27886), .I1 (g27632), .I2 (g24627));
NR2X1 gate23232(.O (g27892), .I1 (g27546), .I2 (g14711));
NR2X1 gate23233(.O (g27896), .I1 (g27632), .I2 (g1222));
NR3X1 gate23234(.O (g27897), .I1 (g6087), .I2 (g27632), .I3 (g25349));
NR3X1 gate23235(.O (g27900), .I1 (g6087), .I2 (g27632), .I3 (g25338));
NR2X1 gate23236(.O (g27906), .I1 (g16127), .I2 (g27656));
NR2X1 gate23237(.O (g27911), .I1 (g16170), .I2 (g27657));
NR2X1 gate23238(.O (g27916), .I1 (g16219), .I2 (g27659));
NR2X1 gate23239(.O (g27917), .I1 (g16220), .I2 (g27660));
NR2X1 gate23240(.O (g27925), .I1 (g16276), .I2 (g27661));
NR2X1 gate23241(.O (g27937), .I1 (g16321), .I2 (g27666));
NR2X1 gate23242(.O (g27950), .I1 (g16367), .I2 (g27673));
NR2X1 gate23243(.O (g27962), .I1 (g16394), .I2 (g27679));
NR2X1 gate23244(.O (g27964), .I1 (g16400), .I2 (g27680));
NR2X1 gate23245(.O (g27980), .I1 (g16428), .I2 (g27681));
NR2X1 gate23246(.O (g27997), .I1 (g16456), .I2 (g27242));
NR2X1 gate23247(.O (g28002), .I1 (g26032), .I2 (g27246));
NR2X1 gate23248(.O (g28029), .I1 (g26033), .I2 (g27247));
NR2X1 gate23249(.O (g28059), .I1 (g26034), .I2 (g27248));
NR2X1 gate23250(.O (g28088), .I1 (g26036), .I2 (g27249));
NR2X1 gate23251(.O (g28145), .I1 (g27629), .I2 (g17001));
NR2X1 gate23252(.O (g28146), .I1 (g27631), .I2 (g17031));
NR2X1 gate23253(.O (g28147), .I1 (g27655), .I2 (g17065));
NR2X1 gate23254(.O (g28148), .I1 (g27658), .I2 (g17100));
NR2X1 gate23255(.O (g28157), .I1 (g13902), .I2 (g27370));
NR2X1 gate23256(.O (g28185), .I1 (g27356), .I2 (g26845));
NR2X1 gate23257(.O (g28189), .I1 (g27359), .I2 (g26853));
NR2X1 gate23258(.O (g28191), .I1 (g27365), .I2 (g26860));
NR2X1 gate23259(.O (g28192), .I1 (g27372), .I2 (g26866));
NR2X1 gate23260(.O (g28199), .I1 (g27250), .I2 (g10024));
NR2X1 gate23261(.O (g28321), .I1 (g27742), .I2 (g10133));
NR2X1 gate23262(.O (g28325), .I1 (g27747), .I2 (g10238));
NR2X1 gate23263(.O (g28328), .I1 (g27755), .I2 (g10340));
NR2X1 gate23264(.O (g28342), .I1 (g15460), .I2 (g28008));
NR2X1 gate23265(.O (g28344), .I1 (g15526), .I2 (g28027));
NR2X1 gate23266(.O (g28345), .I1 (g15527), .I2 (g28028));
NR2X1 gate23267(.O (g28346), .I1 (g15546), .I2 (g28035));
NR2X1 gate23268(.O (g28348), .I1 (g15594), .I2 (g28050));
NR2X1 gate23269(.O (g28349), .I1 (g15595), .I2 (g28051));
NR2X1 gate23270(.O (g28350), .I1 (g15604), .I2 (g28057));
NR2X1 gate23271(.O (g28351), .I1 (g15605), .I2 (g28058));
NR2X1 gate23272(.O (g28352), .I1 (g15624), .I2 (g28065));
NR2X1 gate23273(.O (g28353), .I1 (g15666), .I2 (g28073));
NR2X1 gate23274(.O (g28354), .I1 (g15670), .I2 (g28079));
NR2X1 gate23275(.O (g28355), .I1 (g15671), .I2 (g28080));
NR2X1 gate23276(.O (g28356), .I1 (g15680), .I2 (g28086));
NR2X1 gate23277(.O (g28357), .I1 (g15681), .I2 (g28087));
NR2X1 gate23278(.O (g28358), .I1 (g15700), .I2 (g28094));
NR2X1 gate23279(.O (g28360), .I1 (g15725), .I2 (g28098));
NR2X1 gate23280(.O (g28361), .I1 (g15729), .I2 (g28104));
NR2X1 gate23281(.O (g28362), .I1 (g15730), .I2 (g28105));
NR2X1 gate23282(.O (g28363), .I1 (g15739), .I2 (g28111));
NR2X1 gate23283(.O (g28364), .I1 (g15740), .I2 (g28112));
NR2X1 gate23284(.O (g28366), .I1 (g15765), .I2 (g28116));
NR2X1 gate23285(.O (g28367), .I1 (g15769), .I2 (g28122));
NR2X1 gate23286(.O (g28368), .I1 (g15770), .I2 (g28123));
NR2X1 gate23287(.O (g28371), .I1 (g15793), .I2 (g28127));
NR2X1 gate23288(.O (g28392), .I1 (g27886), .I2 (g22344));
NR2X1 gate23289(.O (g28394), .I1 (g27869), .I2 (g22344));
NR2X1 gate23290(.O (g28397), .I1 (g27869), .I2 (g22344));
NR2X1 gate23291(.O (g28400), .I1 (g27886), .I2 (g22344));
NR2X1 gate23292(.O (g28403), .I1 (g27811), .I2 (g22344));
NR2X1 gate23293(.O (g28406), .I1 (g27824), .I2 (g22344));
NR2X1 gate23294(.O (g28409), .I1 (g24676), .I2 (g27801));
NR2X1 gate23295(.O (g28410), .I1 (g27748), .I2 (g22344));
NR2X1 gate23296(.O (g28413), .I1 (g24695), .I2 (g27809));
NR2X1 gate23297(.O (g28414), .I1 (g27748), .I2 (g22344));
NR2X1 gate23298(.O (g28417), .I1 (g24712), .I2 (g27830));
NR2X1 gate23299(.O (g28418), .I1 (g24723), .I2 (g27846));
NR2X1 gate23300(.O (g28420), .I1 (g16031), .I2 (g28171));
NR2X1 gate23301(.O (g28421), .I1 (g16068), .I2 (g28176));
NR2X1 gate23302(.O (g28425), .I1 (g16133), .I2 (g28188));
NR2X1 gate23303(.O (g28449), .I1 (g27727), .I2 (g26780));
NR2X1 gate23304(.O (g28461), .I1 (g27729), .I2 (g26787));
NR2X1 gate23305(.O (g28470), .I1 (g27671), .I2 (g28193));
NR2X1 gate23306(.O (g28473), .I1 (g27730), .I2 (g26794));
NR2X1 gate23307(.O (g28482), .I1 (g27731), .I2 (g26797));
NR2X1 gate23308(.O (g28488), .I1 (g26755), .I2 (g27719));
NR2X1 gate23309(.O (g28489), .I1 (g26756), .I2 (g27720));
NR2X1 gate23310(.O (g28490), .I1 (g27240), .I2 (g27721));
NR2X1 gate23311(.O (g28495), .I1 (g27244), .I2 (g27723));
NR2X1 gate23312(.O (g28499), .I1 (g26027), .I2 (g27725));
NR2X1 gate23313(.O (g28523), .I1 (g26035), .I2 (g27732));
NR2X1 gate23314(.O (g28525), .I1 (g27245), .I2 (g27726));
NR2X1 gate23315(.O (g28528), .I1 (g26030), .I2 (g27728));
NR2X1 gate23316(.O (g28551), .I1 (g26038), .I2 (g27733));
NR2X1 gate23317(.O (g28578), .I1 (g26039), .I2 (g27734));
NR2X1 gate23318(.O (g28606), .I1 (g26040), .I2 (g27737));
NR2X1 gate23319(.O (g28634), .I1 (g28185), .I2 (g17001));
NR2X1 gate23320(.O (g28635), .I1 (g28189), .I2 (g17031));
NR2X1 gate23321(.O (g28636), .I1 (g28191), .I2 (g17065));
NR2X1 gate23322(.O (g28637), .I1 (g28192), .I2 (g17100));
NR2X1 gate23323(.O (g28654), .I1 (g27770), .I2 (g27355));
NR2X1 gate23324(.O (g28656), .I1 (g27772), .I2 (g27358));
NR2X1 gate23325(.O (g28658), .I1 (g27773), .I2 (g27364));
NR2X1 gate23326(.O (g28661), .I1 (g27775), .I2 (g27371));
NR2X1 gate23327(.O (g28668), .I1 (g27736), .I2 (g10024));
NR2X1 gate23328(.O (g28728), .I1 (g28422), .I2 (g27904));
NR2X1 gate23329(.O (g28731), .I1 (g28423), .I2 (g27908));
NR2X1 gate23330(.O (g28732), .I1 (g14894), .I2 (g28426));
NR2X1 gate23331(.O (g28733), .I1 (g28424), .I2 (g27909));
NR2X1 gate23332(.O (g28735), .I1 (g14957), .I2 (g28430));
NR2X1 gate23333(.O (g28736), .I1 (g28427), .I2 (g27913));
NR2X1 gate23334(.O (g28737), .I1 (g28428), .I2 (g27914));
NR2X1 gate23335(.O (g28738), .I1 (g14975), .I2 (g28433));
NR2X1 gate23336(.O (g28739), .I1 (g28429), .I2 (g27915));
NR2X1 gate23337(.O (g28744), .I1 (g15030), .I2 (g28439));
NR2X1 gate23338(.O (g28745), .I1 (g28431), .I2 (g27922));
NR2X1 gate23339(.O (g28746), .I1 (g15046), .I2 (g28441));
NR2X1 gate23340(.O (g28747), .I1 (g28434), .I2 (g27923));
NR2X1 gate23341(.O (g28748), .I1 (g28435), .I2 (g27924));
NR2X1 gate23342(.O (g28749), .I1 (g15064), .I2 (g28444));
NR2X1 gate23343(.O (g28750), .I1 (g28436), .I2 (g27926));
NR2X1 gate23344(.O (g28754), .I1 (g28440), .I2 (g27931));
NR2X1 gate23345(.O (g28758), .I1 (g15126), .I2 (g28451));
NR2X1 gate23346(.O (g28759), .I1 (g28442), .I2 (g27935));
NR2X1 gate23347(.O (g28760), .I1 (g15142), .I2 (g28453));
NR2X1 gate23348(.O (g28761), .I1 (g28445), .I2 (g27936));
NR2X1 gate23349(.O (g28762), .I1 (g28446), .I2 (g27938));
NR2X1 gate23350(.O (g28763), .I1 (g15160), .I2 (g28456));
NR2X1 gate23351(.O (g28767), .I1 (g28452), .I2 (g27945));
NR2X1 gate23352(.O (g28771), .I1 (g15218), .I2 (g28463));
NR2X1 gate23353(.O (g28772), .I1 (g28454), .I2 (g27949));
NR2X1 gate23354(.O (g28773), .I1 (g15234), .I2 (g28465));
NR2X1 gate23355(.O (g28774), .I1 (g28457), .I2 (g27951));
NR2X1 gate23356(.O (g28778), .I1 (g28464), .I2 (g27963));
NR2X1 gate23357(.O (g28782), .I1 (g15304), .I2 (g28475));
NR2X1 gate23358(.O (g28783), .I1 (g28466), .I2 (g27968));
NR2X1 gate23359(.O (g28784), .I1 (g28468), .I2 (g27970));
NR2X1 gate23360(.O (g28788), .I1 (g28476), .I2 (g27984));
NR2X1 gate23361(.O (g28789), .I1 (g28477), .I2 (g27985));
NR2X1 gate23362(.O (g28790), .I1 (g28478), .I2 (g27991));
NR2X1 gate23363(.O (g28794), .I1 (g28484), .I2 (g28009));
NR2X1 gate23364(.O (g28795), .I1 (g28485), .I2 (g28015));
NR2X1 gate23365(.O (g28802), .I1 (g28492), .I2 (g28036));
NR2X1 gate23366(.O (g28803), .I1 (g28493), .I2 (g28042));
NR2X1 gate23367(.O (g28813), .I1 (g28497), .I2 (g28066));
NR2X1 gate23368(.O (g28874), .I1 (g28657), .I2 (g16221));
NR2X1 gate23369(.O (g28886), .I1 (g28659), .I2 (g16277));
NR2X1 gate23370(.O (g28903), .I1 (g28660), .I2 (g13295));
NR2X1 gate23371(.O (g28920), .I1 (g28662), .I2 (g13322));
NR2X1 gate23372(.O (g28941), .I1 (g28663), .I2 (g13343));
NR3X1 gate23373(.O (g28954), .I1 (g26673), .I2 (g27241), .I3 (g28323));
NR2X1 gate23374(.O (g28963), .I1 (g28664), .I2 (g13365));
NR2X1 gate23375(.O (g28982), .I1 (g28665), .I2 (g28670));
NR2X1 gate23376(.O (g28987), .I1 (g28666), .I2 (g13390));
NR2X1 gate23377(.O (g28990), .I1 (g28667), .I2 (g16457));
NR2X1 gate23378(.O (g29009), .I1 (g28669), .I2 (g28320));
NR2X1 gate23379(.O (g29013), .I1 (g28671), .I2 (g11607));
NR2X1 gate23380(.O (g29016), .I1 (g28672), .I2 (g13487));
NR2X1 gate23381(.O (g29031), .I1 (g28319), .I2 (g28324));
NR2X1 gate23382(.O (g29039), .I1 (g28322), .I2 (g13500));
NR2X1 gate23383(.O (g29063), .I1 (g28326), .I2 (g28329));
NR2X1 gate23384(.O (g29064), .I1 (g28327), .I2 (g28330));
NR2X1 gate23385(.O (g29083), .I1 (g28331), .I2 (g28333));
NR2X1 gate23386(.O (g29090), .I1 (g28332), .I2 (g28334));
NR2X1 gate23387(.O (g29097), .I1 (g28335), .I2 (g28336));
NR2X1 gate23388(.O (g29109), .I1 (g28654), .I2 (g17001));
NR2X1 gate23389(.O (g29110), .I1 (g28656), .I2 (g17031));
NR2X1 gate23390(.O (g29111), .I1 (g28658), .I2 (g17065));
NR2X1 gate23391(.O (g29112), .I1 (g28661), .I2 (g17100));
NR2X1 gate23392(.O (g29113), .I1 (g28381), .I2 (g8907));
NR2X1 gate23393(.O (g29126), .I1 (g28373), .I2 (g27774));
NR2X1 gate23394(.O (g29127), .I1 (g28376), .I2 (g27779));
NR2X1 gate23395(.O (g29128), .I1 (g28380), .I2 (g27783));
NR2X1 gate23396(.O (g29129), .I1 (g28385), .I2 (g27790));
NR2X1 gate23397(.O (g29167), .I1 (g28841), .I2 (g28396));
NR2X1 gate23398(.O (g29169), .I1 (g28843), .I2 (g28398));
NR2X1 gate23399(.O (g29170), .I1 (g28844), .I2 (g28399));
NR2X1 gate23400(.O (g29172), .I1 (g28846), .I2 (g28401));
NR2X1 gate23401(.O (g29173), .I1 (g28847), .I2 (g28402));
NR2X1 gate23402(.O (g29178), .I1 (g28848), .I2 (g28404));
NR2X1 gate23403(.O (g29179), .I1 (g28849), .I2 (g28405));
NR2X1 gate23404(.O (g29181), .I1 (g28850), .I2 (g28407));
NR2X1 gate23405(.O (g29182), .I1 (g28851), .I2 (g28408));
NR2X1 gate23406(.O (g29184), .I1 (g28852), .I2 (g28411));
NR2X1 gate23407(.O (g29185), .I1 (g28853), .I2 (g28412));
NR2X1 gate23408(.O (g29187), .I1 (g28854), .I2 (g28416));
NR2X1 gate23409(.O (g29194), .I1 (g14958), .I2 (g28881));
NR2X1 gate23410(.O (g29195), .I1 (g28880), .I2 (g28438));
NR2X1 gate23411(.O (g29197), .I1 (g15031), .I2 (g28893));
NR2X1 gate23412(.O (g29198), .I1 (g15047), .I2 (g28898));
NR2X1 gate23413(.O (g29199), .I1 (g28892), .I2 (g28448));
NR2X1 gate23414(.O (g29201), .I1 (g15104), .I2 (g28910));
NR2X1 gate23415(.O (g29202), .I1 (g28897), .I2 (g28450));
NR2X1 gate23416(.O (g29204), .I1 (g15127), .I2 (g28915));
NR2X1 gate23417(.O (g29205), .I1 (g15143), .I2 (g28923));
NR2X1 gate23418(.O (g29206), .I1 (g28909), .I2 (g28459));
NR2X1 gate23419(.O (g29207), .I1 (g28914), .I2 (g28460));
NR2X1 gate23420(.O (g29209), .I1 (g15196), .I2 (g28936));
NR2X1 gate23421(.O (g29210), .I1 (g28919), .I2 (g28462));
NR2X1 gate23422(.O (g29212), .I1 (g15219), .I2 (g28944));
NR2X1 gate23423(.O (g29213), .I1 (g15235), .I2 (g28949));
NR2X1 gate23424(.O (g29214), .I1 (g28931), .I2 (g28469));
NR2X1 gate23425(.O (g29215), .I1 (g28935), .I2 (g28471));
NR2X1 gate23426(.O (g29216), .I1 (g28940), .I2 (g28472));
NR2X1 gate23427(.O (g29218), .I1 (g15282), .I2 (g28966));
NR2X1 gate23428(.O (g29219), .I1 (g28948), .I2 (g28474));
NR2X1 gate23429(.O (g29221), .I1 (g15305), .I2 (g28971));
NR2X1 gate23430(.O (g29222), .I1 (g28958), .I2 (g28479));
NR2X1 gate23431(.O (g29223), .I1 (g28962), .I2 (g28480));
NR2X1 gate23432(.O (g29224), .I1 (g28970), .I2 (g28481));
NR2X1 gate23433(.O (g29226), .I1 (g15374), .I2 (g28997));
NR2X1 gate23434(.O (g29227), .I1 (g28986), .I2 (g28486));
NR2X1 gate23435(.O (g29228), .I1 (g28996), .I2 (g28487));
NR2X1 gate23436(.O (g29231), .I1 (g29022), .I2 (g28494));
NR2X1 gate23437(.O (g29303), .I1 (g28716), .I2 (g19112));
NR2X1 gate23438(.O (g29313), .I1 (g28717), .I2 (g19117));
NR2X1 gate23439(.O (g29324), .I1 (g28718), .I2 (g19124));
NR2X1 gate23440(.O (g29333), .I1 (g28719), .I2 (g19131));
NR2X1 gate23441(.O (g29340), .I1 (g28337), .I2 (g28722));
NR2X1 gate23442(.O (g29343), .I1 (g28338), .I2 (g28724));
NR2X1 gate23443(.O (g29345), .I1 (g28339), .I2 (g28726));
NR2X1 gate23444(.O (g29347), .I1 (g28340), .I2 (g28729));
NR2X1 gate23445(.O (g29353), .I1 (g29126), .I2 (g17001));
NR2X1 gate23446(.O (g29354), .I1 (g29127), .I2 (g17031));
NR2X1 gate23447(.O (g29355), .I1 (g29128), .I2 (g17065));
NR2X1 gate23448(.O (g29357), .I1 (g29129), .I2 (g17100));
NR2X1 gate23449(.O (g29399), .I1 (g28834), .I2 (g28378));
NR2X1 gate23450(.O (g29403), .I1 (g28836), .I2 (g28383));
NR2X1 gate23451(.O (g29406), .I1 (g28838), .I2 (g28387));
NR2X1 gate23452(.O (g29409), .I1 (g28840), .I2 (g28389));
NR2X1 gate23453(.O (g29552), .I1 (g29130), .I2 (g29411));
NR2X1 gate23454(.O (g29569), .I1 (g28708), .I2 (g29174));
NR2X1 gate23455(.O (g29570), .I1 (g28709), .I2 (g29175));
NR2X1 gate23456(.O (g29571), .I1 (g28710), .I2 (g29176));
NR2X1 gate23457(.O (g29574), .I1 (g28712), .I2 (g29180));
NR2X1 gate23458(.O (g29576), .I1 (g28713), .I2 (g29183));
NR2X1 gate23459(.O (g29577), .I1 (g28714), .I2 (g29186));
NR2X1 gate23460(.O (g29578), .I1 (g28715), .I2 (g29188));
NR2X1 gate23461(.O (g29579), .I1 (g29399), .I2 (g17001));
NR2X1 gate23462(.O (g29580), .I1 (g29403), .I2 (g17031));
NR2X1 gate23463(.O (g29581), .I1 (g29406), .I2 (g17065));
NR2X1 gate23464(.O (g29582), .I1 (g29409), .I2 (g17100));
NR2X1 gate23465(.O (g29606), .I1 (g13878), .I2 (g29248));
NR2X1 gate23466(.O (g29608), .I1 (g13892), .I2 (g29251));
NR2X1 gate23467(.O (g29609), .I1 (g13900), .I2 (g29252));
NR2X1 gate23468(.O (g29611), .I1 (g13913), .I2 (g29255));
NR2X1 gate23469(.O (g29612), .I1 (g13933), .I2 (g29256));
NR2X1 gate23470(.O (g29613), .I1 (g13941), .I2 (g29257));
NR2X1 gate23471(.O (g29616), .I1 (g13969), .I2 (g29259));
NR2X1 gate23472(.O (g29617), .I1 (g13989), .I2 (g29260));
NR2X1 gate23473(.O (g29618), .I1 (g13997), .I2 (g29261));
NR2X1 gate23474(.O (g29620), .I1 (g14039), .I2 (g29262));
NR2X1 gate23475(.O (g29621), .I1 (g14059), .I2 (g29263));
NR2X1 gate23476(.O (g29623), .I1 (g14130), .I2 (g29264));
NR2X1 gate23477(.O (g29663), .I1 (g29518), .I2 (g29284));
NR2X1 gate23478(.O (g29665), .I1 (g29521), .I2 (g29289));
NR2X1 gate23479(.O (g29667), .I1 (g29524), .I2 (g29294));
NR2X1 gate23480(.O (g29669), .I1 (g29528), .I2 (g29300));
NR2X1 gate23481(.O (g29670), .I1 (g29529), .I2 (g29302));
NR2X1 gate23482(.O (g29671), .I1 (g29534), .I2 (g29310));
NR2X1 gate23483(.O (g29672), .I1 (g29536), .I2 (g29312));
NR2X1 gate23484(.O (g29676), .I1 (g29540), .I2 (g29320));
NR2X1 gate23485(.O (g29677), .I1 (g29543), .I2 (g29321));
NR2X1 gate23486(.O (g29678), .I1 (g29545), .I2 (g29323));
NR2X1 gate23487(.O (g29679), .I1 (g29549), .I2 (g29329));
NR2X1 gate23488(.O (g29680), .I1 (g29553), .I2 (g29330));
NR2X1 gate23489(.O (g29681), .I1 (g29555), .I2 (g29332));
NR2X1 gate23490(.O (g29682), .I1 (g29557), .I2 (g29336));
NR2X1 gate23491(.O (g29683), .I1 (g29559), .I2 (g29337));
NR2X1 gate23492(.O (g29684), .I1 (g29562), .I2 (g29338));
NR2X1 gate23493(.O (g29685), .I1 (g29564), .I2 (g29341));
NR2X1 gate23494(.O (g29686), .I1 (g29566), .I2 (g29342));
NR2X1 gate23495(.O (g29687), .I1 (g29572), .I2 (g29344));
NR2X1 gate23496(.O (g29688), .I1 (g29575), .I2 (g29346));
NR2X1 gate23497(.O (g29703), .I1 (g29583), .I2 (g1917));
NR3X1 gate23498(.O (g29705), .I1 (g6104), .I2 (g29583), .I3 (g25339));
NR2X1 gate23499(.O (g29709), .I1 (g29583), .I2 (g1909));
NR3X1 gate23500(.O (g29710), .I1 (g6104), .I2 (g29583), .I3 (g25412));
NR3X1 gate23501(.O (g29713), .I1 (g6104), .I2 (g29583), .I3 (g25332));
NR2X1 gate23502(.O (g29717), .I1 (g29583), .I2 (g1910));
NR3X1 gate23503(.O (g29718), .I1 (g6104), .I2 (g29583), .I3 (g25409));
NR3X1 gate23504(.O (g29721), .I1 (g6104), .I2 (g29583), .I3 (g25323));
NR2X1 gate23505(.O (g29725), .I1 (g29583), .I2 (g1911));
NR2X1 gate23506(.O (g29727), .I1 (g29583), .I2 (g1912));
NR3X1 gate23507(.O (g29728), .I1 (g6104), .I2 (g29583), .I3 (g25401));
NR2X1 gate23508(.O (g29731), .I1 (g29583), .I2 (g1913));
NR3X1 gate23509(.O (g29732), .I1 (g6104), .I2 (g29583), .I3 (g25387));
NR2X1 gate23510(.O (g29735), .I1 (g23797), .I2 (g29583));
NR2X1 gate23511(.O (g29736), .I1 (g29583), .I2 (g25444));
NR2X1 gate23512(.O (g29740), .I1 (g29583), .I2 (g1914));
NR3X1 gate23513(.O (g29741), .I1 (g6104), .I2 (g29583), .I3 (g25376));
NR2X1 gate23514(.O (g29744), .I1 (g29583), .I2 (g24641));
NR2X1 gate23515(.O (g29747), .I1 (g29583), .I2 (g1916));
NR3X1 gate23516(.O (g29748), .I1 (g6104), .I2 (g29583), .I3 (g25363));
NR3X1 gate23517(.O (g29751), .I1 (g6104), .I2 (g29583), .I3 (g25352));
NR2X1 gate23518(.O (g29754), .I1 (g16178), .I2 (g29607));
NR2X1 gate23519(.O (g29755), .I1 (g16229), .I2 (g29610));
NR2X1 gate23520(.O (g29756), .I1 (g16284), .I2 (g29614));
NR2X1 gate23521(.O (g29757), .I1 (g16285), .I2 (g29615));
NR2X1 gate23522(.O (g29758), .I1 (g16335), .I2 (g29619));
NR2X1 gate23523(.O (g29759), .I1 (g16379), .I2 (g29622));
NR2X1 gate23524(.O (g29760), .I1 (g16411), .I2 (g29624));
NR3X1 gate23525(.O (g29761), .I1 (g28707), .I2 (g28711), .I3 (g29466));
NR2X1 gate23526(.O (g29762), .I1 (g16432), .I2 (g29625));
NR2X1 gate23527(.O (g29763), .I1 (g16438), .I2 (g29626));
NR2X1 gate23528(.O (g29764), .I1 (g16462), .I2 (g29464));
NR2X1 gate23529(.O (g29765), .I1 (g13492), .I2 (g29465));
NR2X1 gate23530(.O (g29766), .I1 (g29467), .I2 (g19142));
NR2X1 gate23531(.O (g29767), .I1 (g29468), .I2 (g19143));
NR2X1 gate23532(.O (g29768), .I1 (g29469), .I2 (g19146));
NR2X1 gate23533(.O (g29769), .I1 (g29470), .I2 (g19148));
NR2X1 gate23534(.O (g29770), .I1 (g29471), .I2 (g29196));
NR2X1 gate23535(.O (g29771), .I1 (g29472), .I2 (g29200));
NR2X1 gate23536(.O (g29772), .I1 (g29473), .I2 (g29203));
NR2X1 gate23537(.O (g29773), .I1 (g29474), .I2 (g29208));
NR2X1 gate23538(.O (g29774), .I1 (g29475), .I2 (g29211));
NR2X1 gate23539(.O (g29775), .I1 (g29476), .I2 (g29217));
NR2X1 gate23540(.O (g29776), .I1 (g29477), .I2 (g29220));
NR2X1 gate23541(.O (g29777), .I1 (g29478), .I2 (g29225));
NR2X1 gate23542(.O (g29778), .I1 (g29479), .I2 (g29229));
NR2X1 gate23543(.O (g29779), .I1 (g13943), .I2 (g29502));
NR2X1 gate23544(.O (g29780), .I1 (g29480), .I2 (g29232));
NR2X1 gate23545(.O (g29781), .I1 (g29481), .I2 (g29233));
NR2X1 gate23546(.O (g29782), .I1 (g29482), .I2 (g29234));
NR2X1 gate23547(.O (g29783), .I1 (g29483), .I2 (g29235));
NR2X1 gate23548(.O (g29784), .I1 (g29484), .I2 (g29236));
NR2X1 gate23549(.O (g29785), .I1 (g29485), .I2 (g29238));
NR2X1 gate23550(.O (g29786), .I1 (g29486), .I2 (g29239));
NR2X1 gate23551(.O (g29787), .I1 (g29487), .I2 (g29240));
NR2X1 gate23552(.O (g29788), .I1 (g29488), .I2 (g29241));
NR2X1 gate23553(.O (g29789), .I1 (g29489), .I2 (g29242));
NR2X1 gate23554(.O (g29791), .I1 (g29490), .I2 (g29243));
NR2X1 gate23555(.O (g29912), .I1 (g24676), .I2 (g29716));
NR2X1 gate23556(.O (g29914), .I1 (g24695), .I2 (g29724));
NR2X1 gate23557(.O (g29916), .I1 (g24712), .I2 (g29726));
NR2X1 gate23558(.O (g29918), .I1 (g29744), .I2 (g22367));
NR2X1 gate23559(.O (g29919), .I1 (g29736), .I2 (g22367));
NR2X1 gate23560(.O (g29920), .I1 (g24723), .I2 (g29739));
NR2X1 gate23561(.O (g29921), .I1 (g29736), .I2 (g22367));
NR2X1 gate23562(.O (g29922), .I1 (g29744), .I2 (g22367));
NR2X1 gate23563(.O (g29924), .I1 (g29710), .I2 (g22367));
NR2X1 gate23564(.O (g29926), .I1 (g29718), .I2 (g22367));
NR2X1 gate23565(.O (g29928), .I1 (g29673), .I2 (g22367));
NR2X1 gate23566(.O (g29929), .I1 (g29673), .I2 (g22367));
NR2X1 gate23567(.O (g29936), .I1 (g16049), .I2 (g29790));
NR2X1 gate23568(.O (g29939), .I1 (g16102), .I2 (g29792));
NR2X1 gate23569(.O (g29941), .I1 (g16182), .I2 (g29793));
NR2X1 gate23570(.O (g30010), .I1 (g29520), .I2 (g29942));
NR2X1 gate23571(.O (g30011), .I1 (g29522), .I2 (g29944));
NR2X1 gate23572(.O (g30012), .I1 (g29523), .I2 (g29945));
NR2X1 gate23573(.O (g30013), .I1 (g29525), .I2 (g29946));
NR2X1 gate23574(.O (g30014), .I1 (g29526), .I2 (g29947));
NR2X1 gate23575(.O (g30015), .I1 (g29527), .I2 (g29948));
NR2X1 gate23576(.O (g30016), .I1 (g29531), .I2 (g29949));
NR2X1 gate23577(.O (g30017), .I1 (g29532), .I2 (g29950));
NR2X1 gate23578(.O (g30018), .I1 (g29533), .I2 (g29951));
NR2X1 gate23579(.O (g30019), .I1 (g29538), .I2 (g29952));
NR2X1 gate23580(.O (g30020), .I1 (g29539), .I2 (g29953));
NR2X1 gate23581(.O (g30021), .I1 (g29541), .I2 (g29954));
NR2X1 gate23582(.O (g30022), .I1 (g29547), .I2 (g29955));
NR2X1 gate23583(.O (g30023), .I1 (g29548), .I2 (g29956));
NR2X1 gate23584(.O (g30024), .I1 (g29550), .I2 (g29957));
NR2X1 gate23585(.O (g30025), .I1 (g29558), .I2 (g29958));
NR2X1 gate23586(.O (g30026), .I1 (g29560), .I2 (g29959));
NR2X1 gate23587(.O (g30027), .I1 (g29565), .I2 (g29960));
NR2X1 gate23588(.O (g30028), .I1 (g29567), .I2 (g29961));
NR2X1 gate23589(.O (g30029), .I1 (g29573), .I2 (g29962));
NR2X1 gate23590(.O (g30030), .I1 (g24676), .I2 (g29923));
NR2X1 gate23591(.O (g30031), .I1 (g24695), .I2 (g29925));
NR2X1 gate23592(.O (g30032), .I1 (g24712), .I2 (g29927));
NR2X1 gate23593(.O (g30033), .I1 (g24723), .I2 (g29931));
NR2X1 gate23594(.O (g30053), .I1 (g29963), .I2 (g16286));
NR2X1 gate23595(.O (g30054), .I1 (g29964), .I2 (g16336));
NR2X1 gate23596(.O (g30055), .I1 (g29965), .I2 (g13326));
NR2X1 gate23597(.O (g30056), .I1 (g29966), .I2 (g13345));
NR2X1 gate23598(.O (g30057), .I1 (g29967), .I2 (g13368));
NR2X1 gate23599(.O (g30058), .I1 (g29968), .I2 (g13395));
NR2X1 gate23600(.O (g30059), .I1 (g29969), .I2 (g29811));
NR2X1 gate23601(.O (g30060), .I1 (g29970), .I2 (g11612));
NR2X1 gate23602(.O (g30061), .I1 (g29971), .I2 (g13493));
NR2X1 gate23603(.O (g30062), .I1 (g29810), .I2 (g29815));
NR2X1 gate23604(.O (g30063), .I1 (g29812), .I2 (g11637));
NR2X1 gate23605(.O (g30064), .I1 (g29813), .I2 (g13506));
NR2X1 gate23606(.O (g30065), .I1 (g29814), .I2 (g29817));
NR2X1 gate23607(.O (g30066), .I1 (g29816), .I2 (g13517));
NR2X1 gate23608(.O (g30067), .I1 (g29818), .I2 (g29820));
NR2X1 gate23609(.O (g30068), .I1 (g29819), .I2 (g29821));
NR2X1 gate23610(.O (g30069), .I1 (g29822), .I2 (g29828));
NR2X1 gate23611(.O (g30070), .I1 (g29827), .I2 (g29833));
NR2X1 gate23612(.O (g30071), .I1 (g29834), .I2 (g29839));
NR2X1 gate23613(.O (g30072), .I1 (g29910), .I2 (g8947));
NR2X1 gate23614(.O (g30245), .I1 (g16074), .I2 (g30077));
NR2X1 gate23615(.O (g30246), .I1 (g16107), .I2 (g30079));
NR2X1 gate23616(.O (g30247), .I1 (g16112), .I2 (g30080));
NR2X1 gate23617(.O (g30248), .I1 (g16139), .I2 (g30081));
NR2X1 gate23618(.O (g30249), .I1 (g16158), .I2 (g30082));
NR2X1 gate23619(.O (g30250), .I1 (g16163), .I2 (g30083));
NR2X1 gate23620(.O (g30251), .I1 (g16198), .I2 (g30085));
NR2X1 gate23621(.O (g30252), .I1 (g16217), .I2 (g30086));
NR2X1 gate23622(.O (g30253), .I1 (g16222), .I2 (g30087));
NR2X1 gate23623(.O (g30254), .I1 (g16242), .I2 (g30088));
NR2X1 gate23624(.O (g30255), .I1 (g16263), .I2 (g30089));
NR2X1 gate23625(.O (g30256), .I1 (g16282), .I2 (g30090));
NR2X1 gate23626(.O (g30257), .I1 (g16290), .I2 (g30091));
NR2X1 gate23627(.O (g30258), .I1 (g16291), .I2 (g30092));
NR2X1 gate23628(.O (g30259), .I1 (g16301), .I2 (g30093));
NR2X1 gate23629(.O (g30260), .I1 (g16322), .I2 (g30094));
NR2X1 gate23630(.O (g30261), .I1 (g16342), .I2 (g30095));
NR2X1 gate23631(.O (g30262), .I1 (g16343), .I2 (g30096));
NR2X1 gate23632(.O (g30263), .I1 (g16344), .I2 (g30097));
NR2X1 gate23633(.O (g30264), .I1 (g16348), .I2 (g30098));
NR2X1 gate23634(.O (g30265), .I1 (g16349), .I2 (g30099));
NR2X1 gate23635(.O (g30266), .I1 (g16359), .I2 (g30100));
NR2X1 gate23636(.O (g30267), .I1 (g16380), .I2 (g30101));
NR2X1 gate23637(.O (g30268), .I1 (g16382), .I2 (g30102));
NR2X1 gate23638(.O (g30269), .I1 (g16386), .I2 (g30103));
NR2X1 gate23639(.O (g30270), .I1 (g16387), .I2 (g30104));
NR2X1 gate23640(.O (g30271), .I1 (g16388), .I2 (g30105));
NR2X1 gate23641(.O (g30272), .I1 (g16392), .I2 (g30106));
NR2X1 gate23642(.O (g30273), .I1 (g16393), .I2 (g30107));
NR2X1 gate23643(.O (g30274), .I1 (g16403), .I2 (g30108));
NR2X1 gate23644(.O (g30275), .I1 (g16413), .I2 (g30109));
NR2X1 gate23645(.O (g30276), .I1 (g16415), .I2 (g30110));
NR2X1 gate23646(.O (g30277), .I1 (g16418), .I2 (g30111));
NR2X1 gate23647(.O (g30278), .I1 (g16420), .I2 (g30112));
NR2X1 gate23648(.O (g30279), .I1 (g16424), .I2 (g30113));
NR2X1 gate23649(.O (g30280), .I1 (g16425), .I2 (g30114));
NR2X1 gate23650(.O (g30281), .I1 (g16426), .I2 (g30115));
NR2X1 gate23651(.O (g30282), .I1 (g16430), .I2 (g30117));
NR2X1 gate23652(.O (g30283), .I1 (g16431), .I2 (g30118));
NR2X1 gate23653(.O (g30284), .I1 (g16444), .I2 (g29980));
NR2X1 gate23654(.O (g30285), .I1 (g16447), .I2 (g29981));
NR2X1 gate23655(.O (g30286), .I1 (g16449), .I2 (g29982));
NR2X1 gate23656(.O (g30287), .I1 (g16452), .I2 (g29983));
NR2X1 gate23657(.O (g30288), .I1 (g16454), .I2 (g29984));
NR2X1 gate23658(.O (g30289), .I1 (g16458), .I2 (g29985));
NR2X1 gate23659(.O (g30290), .I1 (g16459), .I2 (g29986));
NR2X1 gate23660(.O (g30291), .I1 (g16460), .I2 (g29987));
NR2X1 gate23661(.O (g30292), .I1 (g13477), .I2 (g29988));
NR2X1 gate23662(.O (g30293), .I1 (g13480), .I2 (g29989));
NR2X1 gate23663(.O (g30294), .I1 (g13483), .I2 (g29990));
NR2X1 gate23664(.O (g30295), .I1 (g13485), .I2 (g29991));
NR2X1 gate23665(.O (g30296), .I1 (g13488), .I2 (g29993));
NR2X1 gate23666(.O (g30297), .I1 (g13490), .I2 (g29994));
NR2X1 gate23667(.O (g30298), .I1 (g13496), .I2 (g29995));
NR2X1 gate23668(.O (g30299), .I1 (g13499), .I2 (g29996));
NR2X1 gate23669(.O (g30300), .I1 (g13502), .I2 (g30001));
NR2X1 gate23670(.O (g30301), .I1 (g13504), .I2 (g30002));
NR2X1 gate23671(.O (g30302), .I1 (g13513), .I2 (g30003));
NR2X1 gate23672(.O (g30303), .I1 (g13516), .I2 (g30005));
NR2X1 gate23673(.O (g30304), .I1 (g13527), .I2 (g30007));
NR2X1 gate23674(.O (g30338), .I1 (g14297), .I2 (g30225));
NR2X1 gate23675(.O (g30341), .I1 (g14328), .I2 (g30226));
NR2X1 gate23676(.O (g30356), .I1 (g14419), .I2 (g30227));
NR2X1 gate23677(.O (g30399), .I1 (g30116), .I2 (g30123));
NR2X1 gate23678(.O (g30400), .I1 (g29997), .I2 (g30127));
NR2X1 gate23679(.O (g30401), .I1 (g29998), .I2 (g30128));
NR2X1 gate23680(.O (g30402), .I1 (g29999), .I2 (g30129));
NR2X1 gate23681(.O (g30403), .I1 (g30004), .I2 (g30131));
NR2X1 gate23682(.O (g30404), .I1 (g30006), .I2 (g30132));
NR2X1 gate23683(.O (g30405), .I1 (g30008), .I2 (g30133));
NR2X1 gate23684(.O (g30406), .I1 (g30009), .I2 (g30138));
NR2X1 gate23685(.O (g30455), .I1 (g13953), .I2 (g30216));
NR2X1 gate23686(.O (g30468), .I1 (g14007), .I2 (g30217));
NR2X1 gate23687(.O (g30470), .I1 (g14023), .I2 (g30218));
NR2X1 gate23688(.O (g30482), .I1 (g14067), .I2 (g30219));
NR2X1 gate23689(.O (g30485), .I1 (g14098), .I2 (g30220));
NR2X1 gate23690(.O (g30487), .I1 (g14114), .I2 (g30221));
NR2X1 gate23691(.O (g30500), .I1 (g14182), .I2 (g30222));
NR2X1 gate23692(.O (g30503), .I1 (g14213), .I2 (g30223));
NR2X1 gate23693(.O (g30505), .I1 (g14229), .I2 (g30224));
NR2X1 gate23694(.O (g30566), .I1 (g14327), .I2 (g30398));
NR2X1 gate23695(.O (g30584), .I1 (g30412), .I2 (g2611));
NR3X1 gate23696(.O (g30588), .I1 (g6119), .I2 (g30412), .I3 (g25353));
NR2X1 gate23697(.O (g30593), .I1 (g30412), .I2 (g2603));
NR3X1 gate23698(.O (g30594), .I1 (g6119), .I2 (g30412), .I3 (g25419));
NR3X1 gate23699(.O (g30597), .I1 (g6119), .I2 (g30412), .I3 (g25341));
NR2X1 gate23700(.O (g30601), .I1 (g30412), .I2 (g2604));
NR3X1 gate23701(.O (g30602), .I1 (g6119), .I2 (g30412), .I3 (g25417));
NR3X1 gate23702(.O (g30605), .I1 (g6119), .I2 (g30412), .I3 (g25333));
NR2X1 gate23703(.O (g30608), .I1 (g30412), .I2 (g2605));
NR2X1 gate23704(.O (g30609), .I1 (g30412), .I2 (g2606));
NR3X1 gate23705(.O (g30610), .I1 (g6119), .I2 (g30412), .I3 (g25411));
NR2X1 gate23706(.O (g30613), .I1 (g30412), .I2 (g2607));
NR3X1 gate23707(.O (g30614), .I1 (g6119), .I2 (g30412), .I3 (g25403));
NR2X1 gate23708(.O (g30617), .I1 (g23850), .I2 (g30412));
NR2X1 gate23709(.O (g30618), .I1 (g30412), .I2 (g25449));
NR2X1 gate23710(.O (g30621), .I1 (g30412), .I2 (g2608));
NR3X1 gate23711(.O (g30622), .I1 (g6119), .I2 (g30412), .I3 (g25393));
NR2X1 gate23712(.O (g30625), .I1 (g30412), .I2 (g24660));
NR2X1 gate23713(.O (g30628), .I1 (g30412), .I2 (g2610));
NR3X1 gate23714(.O (g30629), .I1 (g6119), .I2 (g30412), .I3 (g25378));
NR3X1 gate23715(.O (g30632), .I1 (g6119), .I2 (g30412), .I3 (g25366));
NR2X1 gate23716(.O (g30635), .I1 (g16108), .I2 (g30407));
NR2X1 gate23717(.O (g30636), .I1 (g16140), .I2 (g30409));
NR2X1 gate23718(.O (g30637), .I1 (g16141), .I2 (g30410));
NR2X1 gate23719(.O (g30638), .I1 (g16159), .I2 (g30411));
NR2X1 gate23720(.O (g30639), .I1 (g16186), .I2 (g30436));
NR2X1 gate23721(.O (g30640), .I1 (g16187), .I2 (g30437));
NR2X1 gate23722(.O (g30641), .I1 (g16188), .I2 (g30438));
NR2X1 gate23723(.O (g30642), .I1 (g16199), .I2 (g30440));
NR2X1 gate23724(.O (g30643), .I1 (g16200), .I2 (g30441));
NR2X1 gate23725(.O (g30644), .I1 (g16218), .I2 (g30442));
NR2X1 gate23726(.O (g30645), .I1 (g16240), .I2 (g30444));
NR2X1 gate23727(.O (g30646), .I1 (g16241), .I2 (g30445));
NR2X1 gate23728(.O (g30647), .I1 (g16251), .I2 (g30447));
NR2X1 gate23729(.O (g30648), .I1 (g16252), .I2 (g30448));
NR2X1 gate23730(.O (g30649), .I1 (g16253), .I2 (g30449));
NR2X1 gate23731(.O (g30650), .I1 (g16264), .I2 (g30451));
NR2X1 gate23732(.O (g30651), .I1 (g16265), .I2 (g30452));
NR2X1 gate23733(.O (g30652), .I1 (g16283), .I2 (g30453));
NR2X1 gate23734(.O (g30653), .I1 (g16289), .I2 (g30454));
NR2X1 gate23735(.O (g30654), .I1 (g16299), .I2 (g30457));
NR2X1 gate23736(.O (g30655), .I1 (g16300), .I2 (g30458));
NR2X1 gate23737(.O (g30656), .I1 (g16310), .I2 (g30460));
NR2X1 gate23738(.O (g30657), .I1 (g16311), .I2 (g30461));
NR2X1 gate23739(.O (g30658), .I1 (g16312), .I2 (g30462));
NR2X1 gate23740(.O (g30659), .I1 (g16323), .I2 (g30464));
NR2X1 gate23741(.O (g30660), .I1 (g16324), .I2 (g30465));
NR2X1 gate23742(.O (g30661), .I1 (g16345), .I2 (g30467));
NR2X1 gate23743(.O (g30662), .I1 (g16347), .I2 (g30469));
NR2X1 gate23744(.O (g30663), .I1 (g16357), .I2 (g30472));
NR2X1 gate23745(.O (g30664), .I1 (g16358), .I2 (g30473));
NR2X1 gate23746(.O (g30665), .I1 (g16368), .I2 (g30475));
NR2X1 gate23747(.O (g30666), .I1 (g16369), .I2 (g30476));
NR2X1 gate23748(.O (g30667), .I1 (g16370), .I2 (g30477));
NR2X1 gate23749(.O (g30668), .I1 (g16381), .I2 (g30478));
NR2X1 gate23750(.O (g30669), .I1 (g16383), .I2 (g30481));
NR2X1 gate23751(.O (g30670), .I1 (g16389), .I2 (g30484));
NR2X1 gate23752(.O (g30671), .I1 (g16391), .I2 (g30486));
NR2X1 gate23753(.O (g30672), .I1 (g16401), .I2 (g30489));
NR2X1 gate23754(.O (g30673), .I1 (g16402), .I2 (g30490));
NR2X1 gate23755(.O (g30674), .I1 (g16414), .I2 (g30492));
NR2X1 gate23756(.O (g30675), .I1 (g16416), .I2 (g30495));
NR2X1 gate23757(.O (g30676), .I1 (g16419), .I2 (g30496));
NR2X1 gate23758(.O (g30677), .I1 (g16421), .I2 (g30499));
NR2X1 gate23759(.O (g30678), .I1 (g16427), .I2 (g30502));
NR2X1 gate23760(.O (g30679), .I1 (g16429), .I2 (g30504));
NR2X1 gate23761(.O (g30680), .I1 (g16443), .I2 (g30327));
NR2X1 gate23762(.O (g30681), .I1 (g16448), .I2 (g30330));
NR2X1 gate23763(.O (g30682), .I1 (g16450), .I2 (g30333));
NR2X1 gate23764(.O (g30683), .I1 (g16453), .I2 (g30334));
NR2X1 gate23765(.O (g30684), .I1 (g16455), .I2 (g30337));
NR3X1 gate23766(.O (g30685), .I1 (g29992), .I2 (g30000), .I3 (g30372));
NR2X1 gate23767(.O (g30686), .I1 (g16461), .I2 (g30340));
NR2X1 gate23768(.O (g30687), .I1 (g13479), .I2 (g30345));
NR2X1 gate23769(.O (g30688), .I1 (g13484), .I2 (g30348));
NR2X1 gate23770(.O (g30689), .I1 (g13486), .I2 (g30351));
NR2X1 gate23771(.O (g30690), .I1 (g13489), .I2 (g30352));
NR2X1 gate23772(.O (g30691), .I1 (g13491), .I2 (g30355));
NR2X1 gate23773(.O (g30692), .I1 (g13498), .I2 (g30361));
NR2X1 gate23774(.O (g30693), .I1 (g13503), .I2 (g30364));
NR2X1 gate23775(.O (g30694), .I1 (g13505), .I2 (g30367));
NR2X1 gate23776(.O (g30695), .I1 (g13515), .I2 (g30374));
NR2X1 gate23777(.O (g30699), .I1 (g13914), .I2 (g30387));
NR2X1 gate23778(.O (g30700), .I1 (g13952), .I2 (g30388));
NR2X1 gate23779(.O (g30701), .I1 (g13970), .I2 (g30389));
NR2X1 gate23780(.O (g30702), .I1 (g14006), .I2 (g30390));
NR2X1 gate23781(.O (g30703), .I1 (g14022), .I2 (g30391));
NR2X1 gate23782(.O (g30704), .I1 (g14040), .I2 (g30392));
NR2X1 gate23783(.O (g30705), .I1 (g14097), .I2 (g30393));
NR2X1 gate23784(.O (g30706), .I1 (g14113), .I2 (g30394));
NR2X1 gate23785(.O (g30707), .I1 (g14131), .I2 (g30395));
NR2X1 gate23786(.O (g30708), .I1 (g14212), .I2 (g30396));
NR2X1 gate23787(.O (g30709), .I1 (g14228), .I2 (g30397));
NR2X1 gate23788(.O (g30780), .I1 (g30625), .I2 (g22387));
NR2X1 gate23789(.O (g30783), .I1 (g30618), .I2 (g22387));
NR2X1 gate23790(.O (g30785), .I1 (g30618), .I2 (g22387));
NR2X1 gate23791(.O (g30786), .I1 (g30625), .I2 (g22387));
NR2X1 gate23792(.O (g30787), .I1 (g30594), .I2 (g22387));
NR2X1 gate23793(.O (g30788), .I1 (g30602), .I2 (g22387));
NR2X1 gate23794(.O (g30789), .I1 (g30575), .I2 (g22387));
NR2X1 gate23795(.O (g30790), .I1 (g30575), .I2 (g22387));
NR2X1 gate23796(.O (g30796), .I1 (g16069), .I2 (g30696));
NR2X1 gate23797(.O (g30798), .I1 (g16134), .I2 (g30697));
NR2X1 gate23798(.O (g30801), .I1 (g16237), .I2 (g30698));
NR2X1 gate23799(.O (g30929), .I1 (g30728), .I2 (g30736));
NR2X1 gate23800(.O (g30930), .I1 (g30735), .I2 (g30744));
NR2X1 gate23801(.O (g30931), .I1 (g30743), .I2 (g30750));
NR2X1 gate23802(.O (g30932), .I1 (g30754), .I2 (g30757));
NR2X1 gate23803(.O (g30933), .I1 (g30755), .I2 (g30758));
NR2X1 gate23804(.O (g30934), .I1 (g30759), .I2 (g30761));
NR2X1 gate23805(.O (g30935), .I1 (g30760), .I2 (g30762));
NR2X1 gate23806(.O (g30936), .I1 (g30763), .I2 (g30764));
NR2X1 gate23807(.O (g30954), .I1 (g30916), .I2 (g30944));
NR2X1 gate23808(.O (g30955), .I1 (g30918), .I2 (g30945));
NR2X1 gate23809(.O (g30956), .I1 (g30919), .I2 (g30946));
NR2X1 gate23810(.O (g30957), .I1 (g30920), .I2 (g30947));
NR2X1 gate23811(.O (g30958), .I1 (g30922), .I2 (g30948));
NR2X1 gate23812(.O (g30959), .I1 (g30923), .I2 (g30949));
NR2X1 gate23813(.O (g30960), .I1 (g30924), .I2 (g30950));
NR2X1 gate23814(.O (g30961), .I1 (g30925), .I2 (g30951));
NR3X1 gate23815(.O (g30970), .I1 (g30917), .I2 (g30921), .I3 (g30953));
endmodule