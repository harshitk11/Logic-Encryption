
module s5378_0 ( clk, n3065gat, n3066gat, n3067gat, n3068gat, n3069gat, 
        n3070gat, n3071gat, n3072gat, n3073gat, n3074gat, n3075gat, n3076gat, 
        n3077gat, n3078gat, n3079gat, n3080gat, n3081gat, n3082gat, n3083gat, 
        n3084gat, n3085gat, n3086gat, n3087gat, n3088gat, n3089gat, n3090gat, 
        n3091gat, n3092gat, n3093gat, n3094gat, n3095gat, n3097gat, n3098gat, 
        n3099gat, n3100gat, key_1, key_2, key_3, key_4, key_5, key_6, key_7, 
        key_8, key_9, key_10, key_11, key_12, key_13, key_14, key_15, key_16, 
        key_17, key_18, key_19, key_20, key_21, key_22, key_23, key_24, key_25, 
        key_26, key_27, key_28, key_29, key_30, key_31, key_32, key_33, key_34, 
        key_35, key_36, key_37, key_38, key_39, key_40, key_41, key_42, key_43, 
        key_44, key_45, key_46, key_47, key_48, key_49, key_50, key_51, key_52, 
        key_53, key_54, key_55, key_56, key_57, key_58, key_59, key_60, key_61, 
        key_62, key_63, key_64, key_65, key_66, key_67, key_68, key_69, key_70, 
        key_71, key_72, key_73, key_74, key_75, key_76, key_77, key_78, key_79, 
        key_80, key_81, key_82, key_83, key_84, key_85, key_86, key_87, key_88, 
        key_89, key_90, key_91, key_92, key_93, key_94, key_95, key_96, key_97, 
        key_98, key_99, key_100, key_101, key_102, key_103, key_104, key_105, 
        key_106, key_107, key_108, key_109, key_110, key_111, key_112, key_113, 
        key_114, key_115, key_116, key_117, key_118, key_119, key_120, key_121, 
        key_122, key_123, key_124, key_125, key_126, key_127, key_128, 
        n3104gat, n3105gat, n3106gat, n3107gat, n3108gat, n3109gat, n3110gat, 
        n3111gat, n3112gat, n3113gat, n3114gat, n3115gat, n3116gat, n3117gat, 
        n3118gat, n3119gat, n3120gat, n3121gat, n3122gat, n3123gat, n3124gat, 
        n3125gat, n3126gat, n3127gat, n3128gat, n3129gat, n3130gat, n3131gat, 
        n3132gat, n3133gat, n3134gat, n3135gat, n3136gat, n3137gat, n3138gat, 
        n3139gat, n3140gat, n3141gat, n3142gat, n3143gat, n3144gat, n3145gat, 
        n3146gat, n3147gat, n3148gat, n3149gat, n3150gat, n3151gat, n3152gat, 
        test_si, test_so, test_se );
  input clk, n3065gat, n3066gat, n3067gat, n3068gat, n3069gat, n3070gat,
         n3071gat, n3072gat, n3073gat, n3074gat, n3075gat, n3076gat, n3077gat,
         n3078gat, n3079gat, n3080gat, n3081gat, n3082gat, n3083gat, n3084gat,
         n3085gat, n3086gat, n3087gat, n3088gat, n3089gat, n3090gat, n3091gat,
         n3092gat, n3093gat, n3094gat, n3095gat, n3097gat, n3098gat, n3099gat,
         n3100gat, key_1, key_2, key_3, key_4, key_5, key_6, key_7, key_8,
         key_9, key_10, key_11, key_12, key_13, key_14, key_15, key_16, key_17,
         key_18, key_19, key_20, key_21, key_22, key_23, key_24, key_25,
         key_26, key_27, key_28, key_29, key_30, key_31, key_32, key_33,
         key_34, key_35, key_36, key_37, key_38, key_39, key_40, key_41,
         key_42, key_43, key_44, key_45, key_46, key_47, key_48, key_49,
         key_50, key_51, key_52, key_53, key_54, key_55, key_56, key_57,
         key_58, key_59, key_60, key_61, key_62, key_63, key_64, key_65,
         key_66, key_67, key_68, key_69, key_70, key_71, key_72, key_73,
         key_74, key_75, key_76, key_77, key_78, key_79, key_80, key_81,
         key_82, key_83, key_84, key_85, key_86, key_87, key_88, key_89,
         key_90, key_91, key_92, key_93, key_94, key_95, key_96, key_97,
         key_98, key_99, key_100, key_101, key_102, key_103, key_104, key_105,
         key_106, key_107, key_108, key_109, key_110, key_111, key_112,
         key_113, key_114, key_115, key_116, key_117, key_118, key_119,
         key_120, key_121, key_122, key_123, key_124, key_125, key_126,
         key_127, key_128, test_si, test_se;
  output n3104gat, n3105gat, n3106gat, n3107gat, n3108gat, n3109gat, n3110gat,
         n3111gat, n3112gat, n3113gat, n3114gat, n3115gat, n3116gat, n3117gat,
         n3118gat, n3119gat, n3120gat, n3121gat, n3122gat, n3123gat, n3124gat,
         n3125gat, n3126gat, n3127gat, n3128gat, n3129gat, n3130gat, n3131gat,
         n3132gat, n3133gat, n3134gat, n3135gat, n3136gat, n3137gat, n3138gat,
         n3139gat, n3140gat, n3141gat, n3142gat, n3143gat, n3144gat, n3145gat,
         n3146gat, n3147gat, n3148gat, n3149gat, n3150gat, n3151gat, n3152gat,
         test_so;
  wire   n398gat, n402gat, n919gat, n846gat, n394gat, n703gat, n722gat,
         n726gat, n271gat, n160gat, n337gat, n842gat, n341gat, n2522gat,
         n1821gat, n283gat, n165gat, n279gat, n1026gat, n275gat, n2476gat,
         n1298gat, n2468gat, n2526gat, n2464gat, n2102gat, n1763gat, n1197gat,
         n667gat, n1834gat, n1767gat, n2084gat, n2021gat, n2182gat, n2095gat,
         n2040gat, n2266gat, n463gat, n384gat, n470gat, n148gat, n1771gat,
         n1675gat, n1456gat, n1525gat, key_out_4, key_out_6, key_out_5,
         key_out_7, key_out_8, key_out_9, key_out_10, key_out_11, key_out_12,
         key_out_23, key_out_20, key_out_18, key_out_19, key_out_37,
         key_out_24, key_out_46, key_out_32, key_out_106, key_out_17, n748gat,
         n43gat, n55gat, key_out_81, key_out_82, key_out_83, key_out_84,
         key_out_85, key_out_88, key_out_89, key_out_90, n933gat, n504gat,
         n2913gat, n2920gat, n2905gat, n2898gat, n567gat, n2989gat,
         key_out_122, key_out_123, key_out_124, key_out_125, key_out_126,
         key_out_127, key_out_128, n2909gat, n2908gat, n2971gat, key_out_108,
         key_out_110, key_out_111, key_out_112, key_out_114, key_out_115,
         key_out_117, key_out_118, key_out_119, n3010gat, n3016gat, n2579gat,
         n2646gat, n2613gat, n2983gat, n2917gat, n2892gat, n2900gat, n2929gat,
         n2925gat, n2916gat, n2899gat, n2926gat, n2924gat, n2923gat, n3147gat,
         n3142gat, n1620gat, n1827gat, n1606gat, n1610gat, n1793gat, n1516gat,
         n1565gat, n1696gat, n2009gat, n1636gat, n2163gat, n2015gat, n2017gat,
         n2194gat, n2057gat, n2556gat, n2539gat, n2436gat, n2387gat, n2330gat,
         n2396gat, n2198gat, n2197gat, n2196gat, n1882gat, n1613gat, n1391gat,
         n1927gat, n1567gat, n1564gat, n1915gat, n1800gat, n1593gat, n189,
         n191, n192, n196, n197, n220, n221, n240, n690, n711, n712, n720,
         n731, n733, n775, n776, n778, n3139gat, n780, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n806, n807, n811,
         n812, n813, n814, n815, n817, n818, n819, n821, n822, n824, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465;
  assign n3148gat = n3147gat;
  assign n3115gat = n3147gat;
  assign n3112gat = n3147gat;
  assign n3141gat = n3142gat;
  assign n3140gat = n3139gat;

  DFZX1 gate1 ( .D(key_out_17), .TD(test_si), .SEL(test_se), .CK(clk), .Q(
        n1465), .QB(n852) );
  DFZX1 gate2 ( .D(key_out_4), .TD(n1465), .SEL(test_se), .CK(clk), .Q(n398gat) );
  DFZX1 gate4 ( .D(key_out_6), .TD(n398gat), .SEL(test_se), .CK(clk), .Q(
        n402gat) );
  DFZX1 gate6 ( .D(key_out_5), .TD(n402gat), .SEL(test_se), .CK(clk), .Q(
        n919gat) );
  DFZX1 gate8 ( .D(key_out_7), .TD(n919gat), .SEL(test_se), .CK(clk), .Q(
        n846gat) );
  DFZX1 gate10 ( .D(key_out_4), .TD(n846gat), .SEL(test_se), .CK(clk), .Q(
        n394gat) );
  DFZX1 gate12 ( .D(key_out_6), .TD(n394gat), .SEL(test_se), .CK(clk), .Q(
        n703gat) );
  DFZX1 gate14 ( .D(key_out_5), .TD(n703gat), .SEL(test_se), .CK(clk), .Q(
        n722gat) );
  DFZX1 gate16 ( .D(key_out_7), .TD(n722gat), .SEL(test_se), .CK(clk), .Q(
        n726gat) );
  DFZX1 gate18 ( .D(n748gat), .TD(n726gat), .SEL(test_se), .CK(clk), .Q(n1464), 
        .QB(n776) );
  DFZX1 gate19 ( .D(key_out_8), .TD(n1464), .SEL(test_se), .CK(clk), .Q(
        n271gat) );
  DFZX1 gate21 ( .D(key_out_9), .TD(n271gat), .SEL(test_se), .CK(clk), .Q(
        n160gat), .QB(n1354) );
  DFZX1 gate23 ( .D(key_out_10), .TD(n160gat), .SEL(test_se), .CK(clk), .Q(
        n337gat) );
  DFZX1 gate25 ( .D(key_out_11), .TD(n337gat), .SEL(test_se), .CK(clk), .Q(
        n842gat) );
  DFZX1 gate27 ( .D(key_out_12), .TD(n842gat), .SEL(test_se), .CK(clk), .Q(
        n341gat) );
  DFZX1 gate29 ( .D(n43gat), .TD(n341gat), .SEL(test_se), .CK(clk), .Q(
        n2522gat) );
  DFZX1 gate30 ( .D(n1620gat), .TD(n2522gat), .SEL(test_se), .CK(clk), .Q(
        n1363), .QB(n787) );
  DFZX1 gate31 ( .D(n787), .TD(n1363), .SEL(test_se), .CK(clk), .Q(n1463), 
        .QB(n775) );
  DFZX1 gate32 ( .D(n1827gat), .TD(n1463), .SEL(test_se), .CK(clk), .Q(
        n1821gat) );
  DFZX1 gate33 ( .D(n1827gat), .TD(n1821gat), .SEL(test_se), .CK(clk), .Q(
        n1379), .QB(n865) );
  DFZX1 gate34 ( .D(n788), .TD(n1379), .SEL(test_se), .CK(clk), .Q(n1462), 
        .QB(n789) );
  DFZX1 gate35 ( .D(n789), .TD(n1462), .SEL(test_se), .CK(clk), .Q(n1461), 
        .QB(n690) );
  DFZX1 gate36 ( .D(key_out_8), .TD(n1461), .SEL(test_se), .CK(clk), .Q(
        n283gat) );
  DFZX1 gate38 ( .D(key_out_9), .TD(n283gat), .SEL(test_se), .CK(clk), .Q(
        n165gat) );
  DFZX1 gate40 ( .D(key_out_10), .TD(n165gat), .SEL(test_se), .CK(clk), .Q(
        n279gat) );
  DFZX1 gate42 ( .D(key_out_11), .TD(n279gat), .SEL(test_se), .CK(clk), .Q(
        n1026gat) );
  DFZX1 gate44 ( .D(key_out_12), .TD(n1026gat), .SEL(test_se), .CK(clk), .Q(
        n275gat) );
  DFZX1 gate46 ( .D(n55gat), .TD(n275gat), .SEL(test_se), .CK(clk), .Q(
        n2476gat) );
  DFZX1 gate47 ( .D(key_out_81), .TD(n2476gat), .SEL(test_se), .CK(clk), .Q(
        n1355) );
  DFZX1 gate48 ( .D(key_out_82), .TD(n1355), .SEL(test_se), .CK(clk), .Q(n1348) );
  DFZX1 gate49 ( .D(key_out_83), .TD(n1348), .SEL(test_se), .CK(clk), .Q(n1460), .QB(n844) );
  DFZX1 gate50 ( .D(key_out_84), .TD(n1460), .SEL(test_se), .CK(clk), .Q(n1423) );
  DFZX1 gate51 ( .D(key_out_85), .TD(n1423), .SEL(test_se), .CK(clk), .Q(n1424) );
  DFZX1 gate52 ( .D(key_out_17), .TD(n1424), .SEL(test_se), .CK(clk), .Q(
        n1298gat) );
  DFZX1 gate54 ( .D(key_out_88), .TD(n1298gat), .SEL(test_se), .CK(clk), .Q(
        n1346) );
  DFZX1 gate55 ( .D(key_out_89), .TD(n1346), .SEL(test_se), .CK(clk), .Q(n1344), .QB(n862) );
  DFZX1 gate56 ( .D(key_out_90), .TD(n1344), .SEL(test_se), .CK(clk), .Q(n1342) );
  DFZX1 gate57 ( .D(n933gat), .TD(n1342), .SEL(test_se), .CK(clk), .Q(n2468gat) );
  DFZX1 gate58 ( .D(key_out_6), .TD(n2468gat), .SEL(test_se), .CK(clk), .Q(
        n1418) );
  DFZX1 gate59 ( .D(key_out_4), .TD(n1418), .SEL(test_se), .CK(clk), .Q(n1419)
         );
  DFZX1 gate60 ( .D(key_out_7), .TD(n1419), .SEL(test_se), .CK(clk), .Q(n1459), 
        .QB(n859) );
  DFZX1 gate61 ( .D(key_out_5), .TD(n1459), .SEL(test_se), .CK(clk), .Q(n1338)
         );
  DFZX1 gate62 ( .D(n2923gat), .TD(n1338), .SEL(test_se), .CK(clk), .Q(n1349), 
        .QB(n790) );
  DFZX1 gate63 ( .D(n2917gat), .TD(n1349), .SEL(test_se), .CK(clk), .Q(n1350), 
        .QB(n791) );
  DFZX1 gate64 ( .D(n2924gat), .TD(n1350), .SEL(test_se), .CK(clk), .Q(n1380), 
        .QB(n792) );
  DFZX1 gate65 ( .D(n2926gat), .TD(n1380), .SEL(test_se), .CK(clk), .Q(n1337), 
        .QB(n793) );
  DFZX1 gate66 ( .D(n2892gat), .TD(n1337), .SEL(test_se), .CK(clk), .Q(n1458), 
        .QB(n794) );
  DFZX1 gate67 ( .D(n504gat), .TD(n1458), .SEL(test_se), .CK(clk), .Q(n2526gat) );
  DFZX1 gate68 ( .D(n2913gat), .TD(n2526gat), .SEL(test_se), .CK(clk), .Q(
        n1420) );
  DFZX1 gate69 ( .D(n2920gat), .TD(n1420), .SEL(test_se), .CK(clk), .Q(n1347)
         );
  DFZX1 gate70 ( .D(n2905gat), .TD(n1347), .SEL(test_se), .CK(clk), .Q(n1381), 
        .QB(n863) );
  DFZX1 gate71 ( .D(n2900gat), .TD(n1381), .SEL(test_se), .CK(clk), .Q(n1421), 
        .QB(n795) );
  DFZX1 gate72 ( .D(n2925gat), .TD(n1421), .SEL(test_se), .CK(clk), .Q(n1422), 
        .QB(n796) );
  DFZX1 gate73 ( .D(n2929gat), .TD(n1422), .SEL(test_se), .CK(clk), .Q(n1351), 
        .QB(n797) );
  DFZX1 gate74 ( .D(n2898gat), .TD(n1351), .SEL(test_se), .CK(clk), .Q(n1345)
         );
  DFZX1 gate75 ( .D(n2916gat), .TD(n1345), .SEL(test_se), .CK(clk), .Q(n1343), 
        .QB(n798) );
  DFZX1 gate76 ( .D(n2899gat), .TD(n1343), .SEL(test_se), .CK(clk), .Q(n1341), 
        .QB(n799) );
  DFZX1 gate77 ( .D(n567gat), .TD(n1341), .SEL(test_se), .CK(clk), .Q(n2464gat) );
  DFZX1 gate78 ( .D(n2396gat), .TD(n2464gat), .SEL(test_se), .CK(clk), .Q(
        n1382), .QB(n800) );
  DFZX1 gate79 ( .D(n2198gat), .TD(n1382), .SEL(test_se), .CK(clk), .Q(n1383), 
        .QB(n801) );
  DFZX1 gate80 ( .D(n2196gat), .TD(n1383), .SEL(test_se), .CK(clk), .Q(n1457), 
        .QB(n802) );
  DFZX1 gate81 ( .D(n196), .TD(n1457), .SEL(test_se), .CK(clk), .Q(n1384), 
        .QB(n803) );
  DFZX1 gate82 ( .D(n2197gat), .TD(n1384), .SEL(test_se), .CK(clk), .Q(n1385), 
        .QB(n804) );
  DFZX1 gate83 ( .D(n2539gat), .TD(n1385), .SEL(test_se), .CK(clk), .Q(n1375)
         );
  DFZX1 gate84 ( .D(n2330gat), .TD(n1375), .SEL(test_se), .CK(clk), .Q(n1386), 
        .QB(n851) );
  DFZX1 gate85 ( .D(n2387gat), .TD(n1386), .SEL(test_se), .CK(clk), .Q(n1387), 
        .QB(n840) );
  DFZX1 gate86 ( .D(n2556gat), .TD(n1387), .SEL(test_se), .CK(clk), .Q(n1388)
         );
  DFZX1 gate87 ( .D(n2436gat), .TD(n1388), .SEL(test_se), .CK(clk), .Q(n1389)
         );
  DFZX1 gate88 ( .D(n1606gat), .TD(n1389), .SEL(test_se), .CK(clk), .Q(
        n2102gat) );
  DFZX1 gate89 ( .D(n1882gat), .TD(n2102gat), .SEL(test_se), .CK(clk), .Q(
        n1390) );
  DFZX1 gate90 ( .D(n1610gat), .TD(n1390), .SEL(test_se), .CK(clk), .Q(
        n1763gat) );
  DFZX1 gate91 ( .D(n2989gat), .TD(n1763gat), .SEL(test_se), .CK(clk), .Q(
        n1391) );
  DFZX1 gate92 ( .D(key_out_122), .TD(n1391), .SEL(test_se), .CK(clk), .Q(
        n1367) );
  DFZX1 gate93 ( .D(key_out_123), .TD(n1367), .SEL(test_se), .CK(clk), .Q(
        n1368) );
  DFZX1 gate94 ( .D(key_out_124), .TD(n1368), .SEL(test_se), .CK(clk), .Q(
        n1371) );
  DFZX1 gate95 ( .D(key_out_125), .TD(n1371), .SEL(test_se), .CK(clk), .Q(
        n1456), .QB(n841) );
  DFZX1 gate96 ( .D(key_out_126), .TD(n1456), .SEL(test_se), .CK(clk), .Q(
        n1392) );
  DFZX1 gate97 ( .D(key_out_127), .TD(n1392), .SEL(test_se), .CK(clk), .Q(
        n1372), .QB(n861) );
  DFZX1 gate98 ( .D(key_out_128), .TD(n1372), .SEL(test_se), .CK(clk), .Q(
        n1369) );
  DFZX1 gate99 ( .D(n2909gat), .TD(n1369), .SEL(test_se), .CK(clk), .Q(n1370)
         );
  DFZX1 gate100 ( .D(n2908gat), .TD(n1370), .SEL(test_se), .CK(clk), .Q(
        n1197gat) );
  DFZX1 gate101 ( .D(n2971gat), .TD(n1197gat), .SEL(test_se), .CK(clk), .Q(
        n1455), .QB(n1332) );
  DFZX1 gate102 ( .D(key_out_108), .TD(n1455), .SEL(test_se), .CK(clk), .Q(
        n667gat) );
  DFZX1 gate103 ( .D(key_out_110), .TD(n667gat), .SEL(test_se), .CK(clk), .Q(
        n1356), .QB(n858) );
  DFZX1 gate104 ( .D(key_out_111), .TD(n1356), .SEL(test_se), .CK(clk), .Q(
        n1393) );
  DFZX1 gate105 ( .D(key_out_112), .TD(n1393), .SEL(test_se), .CK(clk), .Q(
        n1425) );
  DFZX1 gate106 ( .D(key_out_114), .TD(n1425), .SEL(test_se), .CK(clk), .Q(
        n1340) );
  DFZX1 gate107 ( .D(key_out_115), .TD(n1340), .SEL(test_se), .CK(clk), .Q(
        n1339), .QB(n864) );
  DFZX1 gate108 ( .D(key_out_117), .TD(n1339), .SEL(test_se), .CK(clk), .Q(
        n1454), .QB(n843) );
  DFZX1 gate109 ( .D(key_out_118), .TD(n1454), .SEL(test_se), .CK(clk), .Q(
        n1394), .QB(n856) );
  DFZX1 gate110 ( .D(key_out_119), .TD(n1394), .SEL(test_se), .CK(clk), .Q(
        n1395) );
  DFZX1 gate111 ( .D(n3010gat), .TD(n1395), .SEL(test_se), .CK(clk), .Q(n1331)
         );
  DFZX1 gate112 ( .D(n3016gat), .TD(n1331), .SEL(test_se), .CK(clk), .Q(n1453), 
        .QB(n733) );
  DFZX1 gate113 ( .D(n785), .TD(n1453), .SEL(test_se), .CK(clk), .Q(n1452), 
        .QB(n806) );
  DFZX1 gate114 ( .D(n2579gat), .TD(n1452), .SEL(test_se), .CK(clk), .Q(n1451), 
        .QB(n1377) );
  DFZX1 gate115 ( .D(key_out_106), .TD(n1451), .SEL(test_se), .CK(clk), .Q(
        n1426), .QB(n807) );
  DFZX1 gate116 ( .D(n197), .TD(n1426), .SEL(test_se), .CK(clk), .Q(n1427), 
        .QB(n3128gat) );
  DFZX1 gate117 ( .D(n2194gat), .TD(n1427), .SEL(test_se), .CK(clk), .Q(n1374), 
        .QB(n3127gat) );
  DFZX1 gate118 ( .D(n2057gat), .TD(n1374), .SEL(test_se), .CK(clk), .Q(n1373), 
        .QB(n3126gat) );
  DFZX1 gate119 ( .D(n2646gat), .TD(n1373), .SEL(test_se), .CK(clk), .Q(n1378)
         );
  DFZX1 gate120 ( .D(n786), .TD(n1378), .SEL(test_se), .CK(clk), .Q(n1396), 
        .QB(n811) );
  DFZX1 gate121 ( .D(n2613gat), .TD(n1396), .SEL(test_se), .CK(clk), .Q(n1450), 
        .QB(n731) );
  DFZX1 gate122 ( .D(n191), .TD(n1450), .SEL(test_se), .CK(clk), .Q(n1834gat)
         );
  DFZX1 gate123 ( .D(n192), .TD(n1834gat), .SEL(test_se), .CK(clk), .Q(
        n1767gat) );
  DFZX1 gate124 ( .D(n3149gat), .TD(n1767gat), .SEL(test_se), .CK(clk), .Q(
        n2084gat) );
  DFZX1 gate125 ( .D(key_out_23), .TD(n2084gat), .SEL(test_se), .CK(clk), .Q(
        n1366), .QB(n845) );
  DFZX1 gate126 ( .D(key_out_37), .TD(n1366), .SEL(test_se), .CK(clk), .Q(
        n1397), .QB(n846) );
  DFZX1 gate127 ( .D(n221), .TD(n1397), .SEL(test_se), .CK(clk), .Q(n1398), 
        .QB(n853) );
  DFZX1 gate128 ( .D(n220), .TD(n1398), .SEL(test_se), .CK(clk), .Q(n1399), 
        .QB(n838) );
  DFZX1 gate129 ( .D(key_out_24), .TD(n1399), .SEL(test_se), .CK(clk), .Q(
        n1400), .QB(n842) );
  DFZX1 gate130 ( .D(n800), .TD(n1400), .SEL(test_se), .CK(clk), .Q(n1401), 
        .QB(n836) );
  DFZX1 gate131 ( .D(n801), .TD(n1401), .SEL(test_se), .CK(clk), .Q(n1402), 
        .QB(n848) );
  DFZX1 gate132 ( .D(n803), .TD(n1402), .SEL(test_se), .CK(clk), .Q(n1403), 
        .QB(n839) );
  DFZX1 gate133 ( .D(n804), .TD(n1403), .SEL(test_se), .CK(clk), .Q(n1365), 
        .QB(n847) );
  DFZX1 gate134 ( .D(n802), .TD(n1365), .SEL(test_se), .CK(clk), .Q(n1404), 
        .QB(n837) );
  DFZX1 gate135 ( .D(n1793gat), .TD(n1404), .SEL(test_se), .CK(clk), .Q(n1449), 
        .QB(n720) );
  DFZX1 gate136 ( .D(n782), .TD(n1449), .SEL(test_se), .CK(clk), .Q(n2021gat)
         );
  DFZX1 gate137 ( .D(n1516gat), .TD(n2021gat), .SEL(test_se), .CK(clk), .Q(
        n1405) );
  DFZX1 gate138 ( .D(key_out_46), .TD(n1405), .SEL(test_se), .CK(clk), .Q(
        n1358) );
  DFZX1 gate139 ( .D(n780), .TD(n1358), .SEL(test_se), .CK(clk), .Q(n1357) );
  DFZX1 gate140 ( .D(n1565gat), .TD(n1357), .SEL(test_se), .CK(clk), .Q(n1448), 
        .QB(n815) );
  DFZX1 gate141 ( .D(n815), .TD(n1448), .SEL(test_se), .CK(clk), .Q(n1406) );
  DFZX1 gate142 ( .D(n783), .TD(n1406), .SEL(test_se), .CK(clk), .Q(n1447), 
        .QB(n1333) );
  DFZX1 gate143 ( .D(key_out_18), .TD(n1447), .SEL(test_se), .CK(clk), .Q(
        n1407) );
  DFZX1 gate144 ( .D(key_out_19), .TD(n1407), .SEL(test_se), .CK(clk), .Q(
        n1360) );
  DFZX1 gate145 ( .D(key_out_20), .TD(n1360), .SEL(test_se), .CK(clk), .Q(
        n1376), .QB(n855) );
  DFZX1 gate146 ( .D(n778), .TD(n1376), .SEL(test_se), .CK(clk), .Q(n2182gat)
         );
  DFZX1 gate147 ( .D(n2983gat), .TD(n2182gat), .SEL(test_se), .CK(clk), .Q(
        n1446), .QB(n817) );
  DFZX1 gate148 ( .D(n817), .TD(n1446), .SEL(test_se), .CK(clk), .Q(n1361), 
        .QB(n818) );
  DFZX1 gate149 ( .D(n818), .TD(n1361), .SEL(test_se), .CK(clk), .Q(n1445), 
        .QB(n819) );
  DFZX1 gate150 ( .D(n819), .TD(n1445), .SEL(test_se), .CK(clk), .Q(n1364), 
        .QB(n854) );
  DFZX1 gate151 ( .D(n1696gat), .TD(n1364), .SEL(test_se), .CK(clk), .Q(n1408), 
        .QB(n821) );
  DFZX1 gate152 ( .D(n2009gat), .TD(n1408), .SEL(test_se), .CK(clk), .Q(n1444), 
        .QB(n3106gat) );
  DFZX1 gate153 ( .D(n821), .TD(n1444), .SEL(test_se), .CK(clk), .Q(n1443), 
        .QB(n824) );
  DFZX1 gate154 ( .D(n1636gat), .TD(n1443), .SEL(test_se), .CK(clk), .Q(n1352)
         );
  DFZX1 gate155 ( .D(n813), .TD(n1352), .SEL(test_se), .CK(clk), .Q(n1353) );
  DFZX1 gate159 ( .D(n822), .TD(n1353), .SEL(test_se), .CK(clk), .Q(n2095gat)
         );
  DFZX1 gate160 ( .D(key_out_32), .TD(n2095gat), .SEL(test_se), .CK(clk), .Q(
        n1442), .QB(n827) );
  DFZX1 gate161 ( .D(n827), .TD(n1442), .SEL(test_se), .CK(clk), .Q(n1359) );
  DFZX1 gate162 ( .D(n2163gat), .TD(n1359), .SEL(test_se), .CK(clk), .Q(n1409)
         );
  DFZX1 gate163 ( .D(n189), .TD(n1409), .SEL(test_se), .CK(clk), .Q(n2040gat)
         );
  DFZX1 gate164 ( .D(n2015gat), .TD(n2040gat), .SEL(test_se), .CK(clk), .Q(
        n1441), .QB(n828) );
  DFZX1 gate165 ( .D(n828), .TD(n1441), .SEL(test_se), .CK(clk), .Q(n1410), 
        .QB(n829) );
  DFZX1 gate166 ( .D(n2017gat), .TD(n1410), .SEL(test_se), .CK(clk), .Q(n1440), 
        .QB(n830) );
  DFZX1 gate167 ( .D(n830), .TD(n1440), .SEL(test_se), .CK(clk), .Q(n1439), 
        .QB(n712) );
  DFZX1 gate168 ( .D(n807), .TD(n1439), .SEL(test_se), .CK(clk), .Q(n2266gat)
         );
  DFZX1 gate169 ( .D(n829), .TD(n2266gat), .SEL(test_se), .CK(clk), .Q(n1438), 
        .QB(n831) );
  DFZX1 gate170 ( .D(n831), .TD(n1438), .SEL(test_se), .CK(clk), .Q(n1437), 
        .QB(n832) );
  DFZX1 gate171 ( .D(n832), .TD(n1437), .SEL(test_se), .CK(clk), .Q(n1362), 
        .QB(n833) );
  DFZX1 gate172 ( .D(n833), .TD(n1362), .SEL(test_se), .CK(clk), .Q(n1436), 
        .QB(n834) );
  DFZX1 gate173 ( .D(n834), .TD(n1436), .SEL(test_se), .CK(clk), .Q(n1435), 
        .QB(n711) );
  DFZX1 gate174 ( .D(n811), .TD(n1435), .SEL(test_se), .CK(clk), .Q(n1329) );
  DFZX1 gate175 ( .D(n806), .TD(n1329), .SEL(test_se), .CK(clk), .Q(n1328) );
  DFZX1 gate176 ( .D(n794), .TD(n1328), .SEL(test_se), .CK(clk), .Q(n1411) );
  DFZX1 gate177 ( .D(n791), .TD(n1411), .SEL(test_se), .CK(clk), .Q(n1434), 
        .QB(n849) );
  DFZX1 gate178 ( .D(n795), .TD(n1434), .SEL(test_se), .CK(clk), .Q(n1433), 
        .QB(n850) );
  DFZX1 gate179 ( .D(n797), .TD(n1433), .SEL(test_se), .CK(clk), .Q(n1412) );
  DFZX1 gate180 ( .D(n796), .TD(n1412), .SEL(test_se), .CK(clk), .Q(n463gat)
         );
  DFZX1 gate181 ( .D(n798), .TD(n463gat), .SEL(test_se), .CK(clk), .Q(n1413)
         );
  DFZX1 gate182 ( .D(n799), .TD(n1413), .SEL(test_se), .CK(clk), .Q(n384gat)
         );
  DFZX1 gate183 ( .D(n792), .TD(n384gat), .SEL(test_se), .CK(clk), .Q(n1414)
         );
  DFZX1 gate184 ( .D(n793), .TD(n1414), .SEL(test_se), .CK(clk), .Q(n470gat)
         );
  DFZX1 gate185 ( .D(n790), .TD(n470gat), .SEL(test_se), .CK(clk), .Q(n148gat)
         );
  DFZX1 gate186 ( .D(n824), .TD(n148gat), .SEL(test_se), .CK(clk), .Q(n1432), 
        .QB(n835) );
  DFZX1 gate187 ( .D(n835), .TD(n1432), .SEL(test_se), .CK(clk), .Q(n1330) );
  DFZX1 gate188 ( .D(n1613gat), .TD(n1330), .SEL(test_se), .CK(clk), .Q(
        n1771gat) );
  DFZX1 gate189 ( .D(n1391gat), .TD(n1771gat), .SEL(test_se), .CK(clk), .Q(
        n1336) );
  DFZX1 gate190 ( .D(n1927gat), .TD(n1336), .SEL(test_se), .CK(clk), .Q(n1335)
         );
  DFZX1 gate191 ( .D(n814), .TD(n1335), .SEL(test_se), .CK(clk), .Q(n1675gat)
         );
  DFZX1 gate192 ( .D(n240), .TD(n1675gat), .SEL(test_se), .CK(clk), .Q(n1334)
         );
  DFZX1 gate193 ( .D(n1567gat), .TD(n1334), .SEL(test_se), .CK(clk), .Q(n1415), 
        .QB(n857) );
  DFZX1 gate194 ( .D(n1564gat), .TD(n1415), .SEL(test_se), .CK(clk), .Q(
        n1456gat) );
  DFZX1 gate195 ( .D(n812), .TD(n1456gat), .SEL(test_se), .CK(clk), .Q(
        n1525gat) );
  DFZX1 gate196 ( .D(n1915gat), .TD(n1525gat), .SEL(test_se), .CK(clk), .Q(
        n1431), .QB(n860) );
  DFZX1 gate197 ( .D(n1800gat), .TD(n1431), .SEL(test_se), .CK(clk), .Q(n1417)
         );
  DFZX1 gate198 ( .D(n1593gat), .TD(n1417), .SEL(test_se), .CK(clk), .Q(
        test_so), .QB(n1416) );
  INVCKX2 U670 ( .I(n1243), .O(n1233) );
  OAI12X1 U671 ( .B1(n784), .B2(n1428), .A1(n1243), .O(n1326) );
  TIE0X1 U672 ( .O(n1428) );
  TIE1X1 U673 ( .O(n3147gat) );
  INVCKX1 U674 ( .I(n866), .O(n822) );
  AOI33X1 U675 ( .A1(n867), .A2(n868), .A3(n869), .B1(n870), .B2(n871), .B3(
        n872), .O(n866) );
  NR2X1 U676 ( .I1(n838), .I2(n873), .O(n812) );
  OR2B1XLP U677 ( .I1(n874), .B1(n875), .O(n786) );
  XOR2X1 U678 ( .I1(n876), .I2(n1329), .O(n875) );
  OAI112X1 U679 ( .C1(n846), .C2(n877), .A1(n878), .B1(n838), .O(n876) );
  ND2X1 U680 ( .I1(n879), .I2(n196), .O(n785) );
  XOR2X1 U681 ( .I1(n880), .I2(n1328), .O(n879) );
  ND3X1 U682 ( .I1(n881), .I2(n839), .I3(n882), .O(n880) );
  ND3X1 U683 ( .I1(n883), .I2(n884), .I3(n885), .O(n782) );
  AN4B1XLP U684 ( .I1(n886), .I2(n1410), .I3(n1359), .B1(n887), .O(n3146gat)
         );
  AO13X1 U685 ( .B1(n1330), .B2(n888), .B3(n889), .A1(key_out_32), .O(n887) );
  NR3X1 U686 ( .I1(n827), .I2(n832), .I3(n831), .O(n886) );
  AOI12X1 U687 ( .B1(n1330), .B2(n889), .A1(n189), .O(n3145gat) );
  OAI112X1 U688 ( .C1(n1352), .C2(n890), .A1(n891), .B1(n892), .O(n3139gat) );
  MXL2XLP U689 ( .A(n893), .B(n894), .S(n2989gat), .OB(n892) );
  NR2X1 U690 ( .I1(n1353), .I2(n860), .O(n894) );
  OAI13X1 U691 ( .B1(n1525gat), .B2(n1405), .B3(n895), .A1(n896), .O(n893) );
  MXL2XLP U692 ( .A(n897), .B(n1416), .S(n1417), .OB(n896) );
  AOI12X1 U693 ( .B1(key_out_46), .B2(n898), .A1(n1353), .O(n897) );
  OAI112X1 U694 ( .C1(n899), .C2(n865), .A1(n888), .B1(n900), .O(n891) );
  NR3X1 U695 ( .I1(n901), .I2(n1408), .I3(n3098gat), .O(n900) );
  AN2X1 U696 ( .I1(n3097gat), .I2(n902), .O(n899) );
  AOI33X1 U697 ( .A1(n903), .A2(n904), .A3(n905), .B1(n906), .B2(n860), .B3(
        n907), .O(n890) );
  NR2X1 U698 ( .I1(n1415), .I2(n908), .O(n905) );
  INVCKX1 U699 ( .I(n909), .O(n904) );
  ND2X1 U700 ( .I1(n910), .I2(n911), .O(n3016gat) );
  AN4B1XLP U701 ( .I1(n2522gat), .I2(n2526gat), .I3(n2464gat), .B1(n1332), .O(
        n911) );
  AN4B1XLP U702 ( .I1(n2476gat), .I2(n2468gat), .I3(n1331), .B1(n3090gat), .O(
        n910) );
  AOI112X1 U703 ( .C1(n2182gat), .C2(n912), .A1(n913), .B1(n914), .O(n2983gat)
         );
  OR4B2XLP U704 ( .I1(n1407), .I2(n1360), .B1(n855), .B2(n1333), .O(n912) );
  OAI12X1 U705 ( .B1(n915), .B2(n1456gat), .A1(n916), .O(n3142gat) );
  MXL2XLP U706 ( .A(n917), .B(n918), .S(n2989gat), .OB(n916) );
  NR2X1 U707 ( .I1(n1334), .I2(n857), .O(n918) );
  OAI23X1 U708 ( .B1(n1675gat), .B2(n1405), .B3(n895), .A1(n1335), .A2(n919), 
        .O(n917) );
  AOI112X1 U709 ( .C1(n1336), .C2(n780), .A1(n3149gat), .B1(n920), .O(n919) );
  AOI13X1 U710 ( .B1(n2989gat), .B2(n857), .B3(n903), .A1(n907), .O(n915) );
  ND2X1 U711 ( .I1(n898), .I2(n895), .O(n903) );
  OAI22X1 U712 ( .A1(n921), .A2(n922), .B1(n923), .B2(n924), .O(n3133gat) );
  AOI222X1 U713 ( .A1(n925), .A2(n794), .B1(n926), .B2(n927), .C1(n928), .C2(
        n861), .O(n924) );
  OAI22X1 U714 ( .A1(n929), .A2(n922), .B1(n923), .B2(n930), .O(n3130gat) );
  OA222X1 U715 ( .A1(n931), .A2(n1349), .B1(n932), .B2(n933), .C1(n934), .C2(
        n1367), .O(n930) );
  OAI22X1 U716 ( .A1(n935), .A2(n922), .B1(n923), .B2(n936), .O(n3129gat) );
  AOI222X1 U717 ( .A1(n925), .A2(n793), .B1(n926), .B2(n937), .C1(n928), .C2(
        n3116gat), .O(n936) );
  OAI22X1 U718 ( .A1(n938), .A2(n922), .B1(n923), .B2(n939), .O(n3136gat) );
  AOI222X1 U719 ( .A1(n926), .A2(n940), .B1(n928), .B2(n841), .C1(n925), .C2(
        n859), .O(n939) );
  OAI22X1 U720 ( .A1(n941), .A2(n922), .B1(n923), .B2(n942), .O(n3137gat) );
  OA222X1 U721 ( .A1(n932), .A2(n943), .B1(n934), .B2(n1392), .C1(n931), .C2(
        n1338), .O(n942) );
  OAI22X1 U722 ( .A1(n944), .A2(n922), .B1(n923), .B2(n945), .O(n3132gat) );
  OA222X1 U723 ( .A1(n931), .A2(n1350), .B1(n932), .B2(n946), .C1(n934), .C2(
        n1368), .O(n945) );
  OAI22X1 U724 ( .A1(n947), .A2(n922), .B1(n923), .B2(n948), .O(n3134gat) );
  OA222X1 U725 ( .A1(n932), .A2(n949), .B1(n934), .B2(n1370), .C1(n931), .C2(
        n1419), .O(n948) );
  OAI22X1 U726 ( .A1(n950), .A2(n922), .B1(n923), .B2(n951), .O(n3131gat) );
  OA222X1 U727 ( .A1(n931), .A2(n1380), .B1(n932), .B2(n952), .C1(n934), .C2(
        n1371), .O(n951) );
  OAI22X1 U728 ( .A1(n953), .A2(n922), .B1(n923), .B2(n954), .O(n3135gat) );
  OA222X1 U729 ( .A1(n932), .A2(n955), .B1(n934), .B2(n1369), .C1(n931), .C2(
        n1418), .O(n954) );
  OA12X1 U730 ( .B1(n872), .B2(n956), .A1(n957), .O(n923) );
  MXL2XLP U731 ( .A(n958), .B(n959), .S(n872), .OB(n922) );
  INVCKX1 U732 ( .I(n956), .O(n959) );
  OAI12X1 U733 ( .B1(n960), .B2(n961), .A1(n962), .O(n956) );
  AN4B1XLP U734 ( .I1(n963), .I2(n962), .I3(n964), .B1(n965), .O(n958) );
  OAI222X1 U735 ( .A1(n966), .A2(n967), .B1(n968), .B2(n969), .C1(n970), .C2(
        n971), .O(n2929gat) );
  XNR2X1 U736 ( .I1(n1412), .I2(n972), .O(n969) );
  MXL2XLP U737 ( .A(n973), .B(n974), .S(n975), .OB(n2926gat) );
  XOR2X1 U738 ( .I1(n470gat), .I2(n976), .O(n974) );
  NR2X1 U739 ( .I1(n977), .I2(n978), .O(n976) );
  AOI12X1 U740 ( .B1(n1414), .B2(n849), .A1(n1411), .O(n977) );
  OAI222X1 U741 ( .A1(n973), .A2(n967), .B1(n979), .B2(n968), .C1(n970), .C2(
        n980), .O(n2925gat) );
  XOR2X1 U742 ( .I1(n463gat), .I2(n981), .O(n979) );
  NR2X1 U743 ( .I1(n982), .I2(n972), .O(n981) );
  AOI12X1 U744 ( .B1(n1413), .B2(n850), .A1(n1412), .O(n982) );
  MXL2XLP U745 ( .A(n983), .B(n984), .S(n975), .OB(n2924gat) );
  XNR2X1 U746 ( .I1(n1414), .I2(n985), .O(n984) );
  MXL2XLP U747 ( .A(n986), .B(n987), .S(n975), .OB(n2923gat) );
  XOR2X1 U748 ( .I1(n148gat), .I2(n988), .O(n987) );
  NR2X1 U749 ( .I1(n1414), .I2(n985), .O(n988) );
  ND2X1 U750 ( .I1(n989), .I2(n849), .O(n985) );
  OAI22X1 U751 ( .A1(n970), .A2(n990), .B1(n991), .B2(n967), .O(n2920gat) );
  MXL2XLP U752 ( .A(n991), .B(n992), .S(n975), .OB(n2917gat) );
  XNR2X1 U753 ( .I1(n849), .I2(n989), .O(n992) );
  NR2X1 U754 ( .I1(n978), .I2(n1411), .O(n989) );
  OAI222X1 U755 ( .A1(n993), .A2(n967), .B1(n968), .B2(n994), .C1(n970), .C2(
        n995), .O(n2916gat) );
  XNR2X1 U756 ( .I1(n1413), .I2(n996), .O(n994) );
  OAI22X1 U757 ( .A1(n970), .A2(n997), .B1(n986), .B2(n967), .O(n2913gat) );
  OAI12X1 U758 ( .B1(n998), .B2(n999), .A1(n1000), .O(n2909gat) );
  OAI12X1 U759 ( .B1(n973), .B2(n999), .A1(n1000), .O(n2908gat) );
  OAI22X1 U760 ( .A1(n970), .A2(n1001), .B1(n983), .B2(n967), .O(n2905gat) );
  OAI222X1 U761 ( .A1(n1002), .A2(n967), .B1(n968), .B2(n1003), .C1(n970), 
        .C2(n1004), .O(n2900gat) );
  XNR2X1 U762 ( .I1(n850), .I2(n1005), .O(n1003) );
  OAI222X1 U763 ( .A1(n998), .A2(n967), .B1(n1006), .B2(n968), .C1(n970), .C2(
        n1007), .O(n2899gat) );
  ND2X1 U764 ( .I1(n970), .I2(n967), .O(n968) );
  XOR2X1 U765 ( .I1(n384gat), .I2(n1008), .O(n1006) );
  NR2X1 U766 ( .I1(n1413), .I2(n996), .O(n1008) );
  ND2X1 U767 ( .I1(n1005), .I2(n850), .O(n996) );
  NR2X1 U768 ( .I1(n972), .I2(n1412), .O(n1005) );
  OAI22X1 U769 ( .A1(n970), .A2(n1009), .B1(n1010), .B2(n967), .O(n2898gat) );
  ND3X1 U770 ( .I1(n872), .I2(n870), .I3(n1011), .O(n967) );
  INVCKX1 U771 ( .I(n1012), .O(n872) );
  MXL2XLP U772 ( .A(n1010), .B(n1013), .S(n975), .OB(n2892gat) );
  AOI13X1 U773 ( .B1(n1011), .B2(n1012), .B3(n870), .A1(n1014), .O(n975) );
  INVCKX1 U774 ( .I(n970), .O(n1014) );
  ND3X1 U775 ( .I1(n869), .I2(n1015), .I3(n867), .O(n970) );
  INVCKX1 U776 ( .I(n1016), .O(n869) );
  AN4B1XLP U777 ( .I1(n1017), .I2(n1018), .I3(n960), .B1(n1019), .O(n870) );
  XNR2X1 U778 ( .I1(n1411), .I2(n978), .O(n1013) );
  ND2X1 U779 ( .I1(n1020), .I2(n1021), .O(n3104gat) );
  AOI23X1 U780 ( .B1(n3094gat), .B2(n1022), .B3(n1023), .A1(n1024), .A2(n1018), 
        .O(n1020) );
  INVCKX1 U781 ( .I(n1025), .O(n1023) );
  ND2X1 U782 ( .I1(n1026), .I2(n1027), .O(n3105gat) );
  AOI23X1 U783 ( .B1(n1015), .B2(n1016), .B3(n867), .A1(n1028), .A2(n1018), 
        .O(n1026) );
  INVCKX1 U784 ( .I(n1029), .O(n867) );
  ND2X1 U785 ( .I1(n1030), .I2(n2613gat), .O(n3143gat) );
  ND2X1 U786 ( .I1(n1371), .I2(n1031), .O(n3109gat) );
  ND2X1 U787 ( .I1(n1367), .I2(n1032), .O(n3108gat) );
  OAI12X1 U788 ( .B1(n935), .B2(n957), .A1(n2646gat), .O(n3125gat) );
  INVCKX1 U789 ( .I(n1033), .O(n935) );
  OAI122X1 U790 ( .B1(n1422), .B2(n931), .C1(n1424), .C2(n932), .A1(n1034), 
        .O(n1033) );
  AOI122X1 U791 ( .B1(n1035), .B2(n1036), .C1(n928), .C2(n1037), .A1(n1038), 
        .O(n1034) );
  AOI112X1 U792 ( .C1(n852), .C2(n1039), .A1(n1040), .B1(n1041), .O(n1038) );
  OAI12X1 U793 ( .B1(n941), .B2(n957), .A1(n2971gat), .O(n3124gat) );
  XNR2X1 U794 ( .I1(n1197gat), .I2(n3116gat), .O(n2971gat) );
  OA112X1 U795 ( .C1(n1042), .C2(n932), .A1(n1043), .B1(n1044), .O(n941) );
  OA22X1 U796 ( .A1(n1045), .A2(n1046), .B1(n931), .B2(n1351), .O(n1044) );
  AOI23X1 U797 ( .B1(n1047), .B2(n852), .B3(n1048), .A1(n1049), .A2(n928), .O(
        n1043) );
  OAI12X1 U798 ( .B1(n938), .B2(n957), .A1(n3010gat), .O(n3123gat) );
  XNR2X1 U799 ( .I1(n667gat), .I2(n1037), .O(n3010gat) );
  INVCKX1 U800 ( .I(n1050), .O(n938) );
  OAI122X1 U801 ( .B1(n934), .B2(n1051), .C1(n1421), .C2(n931), .A1(n1052), 
        .O(n1050) );
  MAOI1X1 U802 ( .A1(n1035), .A2(n1053), .B1(n932), .B2(n1423), .O(n1052) );
  OAI12X1 U803 ( .B1(n953), .B2(n957), .A1(n504gat), .O(n3122gat) );
  XOR3X1 U804 ( .I1(n1054), .I2(n1055), .I3(n1350), .O(n504gat) );
  XOR4XLP U805 ( .I1(n1419), .I2(n859), .I3(n794), .I4(n1418), .O(n1055) );
  XOR4XLP U806 ( .I1(n1349), .I2(n1380), .I3(n1337), .I4(n1338), .O(n1054) );
  AOI122X1 U807 ( .B1(n856), .B2(n928), .C1(n798), .C2(n925), .A1(n1056), .O(
        n953) );
  OAI22X1 U808 ( .A1(n1045), .A2(n1057), .B1(n932), .B2(n1344), .O(n1056) );
  OAI12X1 U809 ( .B1(n947), .B2(n957), .A1(n567gat), .O(n3121gat) );
  XOR3X1 U810 ( .I1(n1058), .I2(n1059), .I3(n1347), .O(n567gat) );
  XOR4XLP U811 ( .I1(n1421), .I2(n1422), .I3(n1381), .I4(n1420), .O(n1059) );
  XOR4XLP U812 ( .I1(n1345), .I2(n1351), .I3(n1341), .I4(n1343), .O(n1058) );
  INVCKX1 U813 ( .I(n1060), .O(n947) );
  OAI122X1 U814 ( .B1(n1395), .B2(n934), .C1(n1341), .C2(n931), .A1(n1061), 
        .O(n1060) );
  MAOI1X1 U815 ( .A1(n1035), .A2(n1062), .B1(n932), .B2(n1342), .O(n1061) );
  OAI12X1 U816 ( .B1(n921), .B2(n957), .A1(n55gat), .O(n3120gat) );
  XNR3X1 U817 ( .I1(n1063), .I2(key_91), .I3(n1064), .O(n55gat) );
  XOR4XLP U818 ( .I1(key_98), .I2(n1065), .I3(n943), .I4(n937), .O(n1064) );
  XNR2X1 U819 ( .I1(n1026gat), .I2(key_96), .O(n937) );
  AOI12X1 U820 ( .B1(n1066), .B2(n927), .A1(n1067), .O(n1065) );
  MXL2XLP U821 ( .A(n1068), .B(n1069), .S(n949), .OB(n1067) );
  OR2X1 U822 ( .I1(n927), .I2(n1066), .O(n1069) );
  XOR2X1 U823 ( .I1(n955), .I2(n927), .O(n1068) );
  XOR4XLP U824 ( .I1(n933), .I2(n946), .I3(n940), .I4(n952), .O(n1063) );
  AOI122X1 U825 ( .B1(n1070), .B2(n1035), .C1(n843), .C2(n928), .A1(n1071), 
        .O(n921) );
  OAI22X1 U826 ( .A1(n931), .A2(n1345), .B1(n932), .B2(n1346), .O(n1071) );
  INVCKX1 U827 ( .I(n934), .O(n928) );
  OAI12X1 U828 ( .B1(n944), .B2(n957), .A1(n933gat), .O(n3119gat) );
  OAI22X1 U829 ( .A1(n1072), .A2(n1073), .B1(n1074), .B2(n1075), .O(n933gat)
         );
  XNR2X1 U830 ( .I1(n1073), .I2(key_41), .O(n1075) );
  AOI22X1 U831 ( .A1(n1076), .A2(n1077), .B1(n1078), .B2(n1079), .O(n1074) );
  XOR4XLP U832 ( .I1(n1342), .I2(n1344), .I3(n1346), .I4(key_87), .O(n1073) );
  AOI22X1 U833 ( .A1(n1079), .A2(n1077), .B1(n1076), .B2(n1078), .O(n1072) );
  XNR2X1 U834 ( .I1(n1079), .I2(key_42), .O(n1076) );
  XNR2X1 U835 ( .I1(n1078), .I2(key_43), .O(n1077) );
  XOR4XLP U836 ( .I1(n1348), .I2(n1355), .I3(n844), .I4(key_80), .O(n1078) );
  XNR3X1 U837 ( .I1(n1423), .I2(n1424), .I3(n1042), .O(n1079) );
  INVCKX1 U838 ( .I(n1080), .O(n944) );
  OAI122X1 U839 ( .B1(n1081), .B2(n1045), .C1(n1393), .C2(n934), .A1(n1082), 
        .O(n1080) );
  OA22X1 U840 ( .A1(n931), .A2(n1347), .B1(n932), .B2(n1348), .O(n1082) );
  XOR2X1 U841 ( .I1(n160gat), .I2(key_102), .O(n1081) );
  ND2X1 U842 ( .I1(n2579gat), .I2(n1030), .O(n3144gat) );
  INVCKX1 U843 ( .I(n1083), .O(n1030) );
  OAI122X1 U844 ( .B1(n1405), .B2(n1084), .C1(n1085), .C2(n720), .A1(n1086), 
        .O(n1083) );
  AOI33X1 U845 ( .A1(n920), .A2(n804), .A3(n1087), .B1(n852), .B2(n824), .B3(
        n888), .O(n1086) );
  MXL2XLP U846 ( .A(n1088), .B(n1089), .S(n802), .OB(n1087) );
  ND2X1 U847 ( .I1(n1090), .I2(n1091), .O(n1089) );
  XNR2X1 U848 ( .I1(n1046), .I2(n1037), .O(n1091) );
  XOR4XLP U849 ( .I1(n858), .I2(n1393), .I3(n1092), .I4(n1093), .O(n1037) );
  XOR4XLP U850 ( .I1(key_109), .I2(n1094), .I3(key_116), .I4(key_113), .O(
        n1093) );
  MAOI1X1 U851 ( .A1(n1051), .A2(n864), .B1(n1049), .B2(n1340), .O(n1094) );
  INVCKX1 U852 ( .I(n1095), .O(n1049) );
  XOR4XLP U853 ( .I1(n843), .I2(n1394), .I3(n1425), .I4(n1395), .O(n1092) );
  AOI12X1 U854 ( .B1(n1090), .B2(n858), .A1(n1096), .O(n1088) );
  MXL2XLP U855 ( .A(n1097), .B(n1098), .S(n803), .OB(n1096) );
  AOI122X1 U856 ( .B1(n1099), .B2(n856), .C1(n1100), .C2(n843), .A1(n1101), 
        .O(n1098) );
  OAI22X1 U857 ( .A1(n1425), .A2(n1102), .B1(n1095), .B2(n1103), .O(n1101) );
  XOR2X1 U858 ( .I1(n1339), .I2(key_45), .O(n1095) );
  OA222X1 U859 ( .A1(n1103), .A2(n1051), .B1(n1104), .B2(n1395), .C1(n1105), 
        .C2(n1393), .O(n1097) );
  XOR2X1 U860 ( .I1(n1340), .I2(key_44), .O(n1051) );
  AOI23X1 U861 ( .B1(n1106), .B2(n802), .B3(n1385), .A1(n1107), .A2(n1108), 
        .O(n1085) );
  OAI122X1 U862 ( .B1(n1109), .B2(n1105), .C1(n1110), .C2(n1103), .A1(n1111), 
        .O(n1108) );
  AOI112X1 U863 ( .C1(n1099), .C2(n1112), .A1(n1113), .B1(n1114), .O(n1111) );
  AOI12X1 U864 ( .B1(n2084gat), .B2(n1115), .A1(n1116), .O(n1114) );
  INVCKX1 U865 ( .I(n1090), .O(n1116) );
  AOI112X1 U866 ( .C1(n1115), .C2(n898), .A1(n1102), .B1(n1384), .O(n1113) );
  OAI122X1 U867 ( .B1(n1345), .B2(n1117), .C1(n1346), .C2(n1118), .A1(n1119), 
        .O(n1112) );
  OA22X1 U868 ( .A1(n1120), .A2(n1347), .B1(n1121), .B2(n1348), .O(n1119) );
  ND2X1 U869 ( .I1(n800), .I2(n801), .O(n1103) );
  AOI122X1 U870 ( .B1(n1122), .B2(n798), .C1(n1123), .C2(n862), .A1(n1124), 
        .O(n1110) );
  OAI22X1 U871 ( .A1(n1342), .A2(n1121), .B1(n1341), .B2(n1120), .O(n1124) );
  AOI122X1 U872 ( .B1(n1122), .B2(n863), .C1(n1123), .C2(n844), .A1(n1125), 
        .O(n1109) );
  OAI22X1 U873 ( .A1(n1355), .A2(n1121), .B1(n1420), .B2(n1120), .O(n1125) );
  OAI122X1 U874 ( .B1(n1126), .B2(n1104), .C1(n1127), .C2(n1105), .A1(n1128), 
        .O(n1106) );
  AOI22X1 U875 ( .A1(n1129), .A2(n1090), .B1(n1130), .B2(n1131), .O(n1128) );
  OAI22X1 U876 ( .A1(n1042), .A2(n1118), .B1(n1351), .B2(n1117), .O(n1131) );
  XOR2X1 U877 ( .I1(n1298gat), .I2(key_86), .O(n1042) );
  MXL2XLP U878 ( .A(n1421), .B(n1423), .S(n3149gat), .OB(n1129) );
  INVCKX1 U879 ( .I(n1132), .O(n1127) );
  OAI122X1 U880 ( .B1(n1120), .B2(n1349), .C1(n1117), .C2(n1380), .A1(n1133), 
        .O(n1132) );
  OA22X1 U881 ( .A1(n952), .A2(n1118), .B1(n933), .B2(n1121), .O(n1133) );
  XOR2X1 U882 ( .I1(n283gat), .I2(key_92), .O(n933) );
  INVCKX1 U883 ( .I(n1123), .O(n1118) );
  XOR2X1 U884 ( .I1(n279gat), .I2(key_94), .O(n952) );
  INVCKX1 U885 ( .I(n1122), .O(n1117) );
  INVCKX1 U886 ( .I(n1099), .O(n1104) );
  NR2X1 U887 ( .I1(n801), .I2(n1382), .O(n1099) );
  AOI122X1 U888 ( .B1(n1122), .B2(n794), .C1(n1123), .C2(n927), .A1(n1134), 
        .O(n1126) );
  OAI22X1 U889 ( .A1(n946), .A2(n1121), .B1(n1350), .B2(n1120), .O(n1134) );
  ND2X1 U890 ( .I1(n1384), .I2(n1135), .O(n1120) );
  ND2X1 U891 ( .I1(n1384), .I2(n3149gat), .O(n1121) );
  XOR2X1 U892 ( .I1(n165gat), .I2(key_93), .O(n946) );
  XNR2X1 U893 ( .I1(n275gat), .I2(key_99), .O(n927) );
  NR2X1 U894 ( .I1(n1384), .I2(n1135), .O(n1123) );
  NR2X1 U895 ( .I1(n3149gat), .I2(n1384), .O(n1122) );
  INVCKX1 U896 ( .I(n1136), .O(n1084) );
  OAI23X1 U897 ( .B1(n2989gat), .B2(n1353), .B3(n1135), .A1(n1137), .A2(n1352), 
        .O(n1136) );
  INVCKX1 U898 ( .I(n907), .O(n1137) );
  XNR2X1 U899 ( .I1(n1138), .I2(key_34), .O(n907) );
  ND2X1 U900 ( .I1(n3149gat), .I2(n2989gat), .O(n1138) );
  INVCKX1 U901 ( .I(n3149gat), .O(n1135) );
  OAI12X1 U902 ( .B1(n950), .B2(n957), .A1(n43gat), .O(n3118gat) );
  XOR4XLP U903 ( .I1(n1139), .I2(n1140), .I3(n1036), .I4(n1141), .O(n43gat) );
  XOR4XLP U904 ( .I1(n1142), .I2(n1046), .I3(n1057), .I4(n1143), .O(n1141) );
  XNR2X1 U905 ( .I1(n842gat), .I2(key_104), .O(n1036) );
  MUX4X1 U906 ( .A(n1144), .B(n1145), .C(n1145), .D(n1144), .S0(n1146), .S1(
        n1147), .O(n1140) );
  XOR2X1 U907 ( .I1(n1354), .I2(key_102), .O(n1147) );
  INVCKX1 U908 ( .I(n1070), .O(n1139) );
  XNR2X1 U909 ( .I1(n341gat), .I2(key_105), .O(n1070) );
  INVCKX1 U910 ( .I(n1148), .O(n950) );
  OAI122X1 U911 ( .B1(n1425), .B2(n934), .C1(n1381), .C2(n931), .A1(n1149), 
        .O(n1148) );
  AOI22X1 U912 ( .A1(n1035), .A2(n1144), .B1(n926), .B2(n844), .O(n1149) );
  INVCKX1 U913 ( .I(n932), .O(n926) );
  OAI12X1 U914 ( .B1(n929), .B2(n957), .A1(n748gat), .O(n3117gat) );
  XOR4XLP U915 ( .I1(n1150), .I2(n1151), .I3(n1152), .I4(n1153), .O(n748gat)
         );
  XOR4XLP U916 ( .I1(key_73), .I2(key_72), .I3(n3089gat), .I4(key_74), .O(
        n1153) );
  XNR2X1 U917 ( .I1(n1012), .I2(n871), .O(n1152) );
  MXL2XLP U918 ( .A(n1154), .B(n1155), .S(n1156), .OB(n1151) );
  XNR2X1 U919 ( .I1(n1157), .I2(n1158), .O(n1155) );
  AOI12X1 U920 ( .B1(n1158), .B2(n1157), .A1(n962), .O(n1154) );
  OAI112X1 U921 ( .C1(n963), .C2(n964), .A1(n962), .B1(n1156), .O(n957) );
  INVCKX1 U922 ( .I(n1159), .O(n929) );
  OAI122X1 U923 ( .B1(n1356), .B2(n934), .C1(n1420), .C2(n931), .A1(n1160), 
        .O(n1159) );
  MAOI1X1 U924 ( .A1(n1035), .A2(n1146), .B1(n932), .B2(n1355), .O(n1160) );
  ND2X1 U925 ( .I1(n1047), .I2(n1040), .O(n932) );
  INVCKX1 U926 ( .I(n1045), .O(n1035) );
  ND2X1 U927 ( .I1(n1041), .I2(n1040), .O(n1045) );
  INVCKX1 U928 ( .I(n1048), .O(n1040) );
  INVCKX1 U929 ( .I(n925), .O(n931) );
  NR2X1 U930 ( .I1(n1039), .I2(n1048), .O(n925) );
  INVCKX1 U931 ( .I(n1161), .O(n1039) );
  ND2X1 U932 ( .I1(n1041), .I2(n1048), .O(n934) );
  AOI22X1 U933 ( .A1(n1012), .A2(n1162), .B1(n1163), .B2(n1150), .O(n1048) );
  NR2X1 U934 ( .I1(n1161), .I2(n1047), .O(n1041) );
  NR2X1 U935 ( .I1(n964), .I2(n960), .O(n1047) );
  NR2X1 U936 ( .I1(n1156), .I2(n1164), .O(n960) );
  NR2X1 U937 ( .I1(n1165), .I2(n1011), .O(n964) );
  NR2X1 U938 ( .I1(n961), .I2(n963), .O(n1161) );
  NR2X1 U939 ( .I1(n1165), .I2(n1019), .O(n963) );
  INVCKX1 U940 ( .I(n1150), .O(n1019) );
  INVCKX1 U941 ( .I(n1162), .O(n1165) );
  NR2X1 U942 ( .I1(n1011), .I2(n1164), .O(n961) );
  OAI112X1 U943 ( .C1(n1022), .C2(n1166), .A1(n1167), .B1(n1168), .O(n3152gat)
         );
  INVCKX1 U944 ( .I(n1028), .O(n1167) );
  NR3X1 U945 ( .I1(n871), .I2(n1156), .I3(n1169), .O(n1028) );
  ND2X1 U946 ( .I1(n1015), .I2(n1016), .O(n1166) );
  ND2X1 U947 ( .I1(n1170), .I2(n1372), .O(n3111gat) );
  ND2X1 U948 ( .I1(n1368), .I2(n1171), .O(n3110gat) );
  OAI112X1 U949 ( .C1(n1172), .C2(n1025), .A1(n1173), .B1(n1174), .O(n3151gat)
         );
  INVCKX1 U950 ( .I(n1024), .O(n1173) );
  NR3X1 U951 ( .I1(n965), .I2(n1011), .I3(n1169), .O(n1024) );
  ND2X1 U952 ( .I1(n1369), .I2(n1175), .O(n3113gat) );
  ND2X1 U953 ( .I1(n1176), .I2(n1177), .O(n3114gat) );
  XNR2X1 U954 ( .I1(n841), .I2(key_21), .O(n1177) );
  OAI12X1 U955 ( .B1(n1409), .B2(n1178), .A1(n1179), .O(n3150gat) );
  INVCKX1 U956 ( .I(n1144), .O(n1178) );
  XNR2X1 U957 ( .I1(n1145), .I2(key_121), .O(n1144) );
  XOR2X1 U958 ( .I1(n337gat), .I2(key_103), .O(n1145) );
  OA12X1 U959 ( .B1(n1180), .B2(n1181), .A1(n1182), .O(n2646gat) );
  XOR2X1 U960 ( .I1(n1183), .I2(key_13), .O(n1182) );
  OAI112X1 U961 ( .C1(n1373), .C2(key_out_18), .A1(n1184), .B1(n1181), .O(
        n1183) );
  OAI22X1 U962 ( .A1(n1426), .A2(n1185), .B1(n1186), .B2(n1187), .O(n1181) );
  AOI12X1 U963 ( .B1(n1426), .B2(n1188), .A1(n1427), .O(n1186) );
  INVCKX1 U964 ( .I(key_107), .O(n1188) );
  NR2X1 U965 ( .I1(key_107), .I2(n1427), .O(n1185) );
  OA12X1 U966 ( .B1(key_out_18), .B2(n1373), .A1(n1184), .O(n1180) );
  OR2X1 U967 ( .I1(key_out_19), .I2(n1374), .O(n1184) );
  MUX2X1 U968 ( .A(n1189), .B(n1190), .S(n1396), .O(n2613gat) );
  XOR2X1 U969 ( .I1(n1191), .I2(n1192), .O(n1190) );
  OAI22X1 U970 ( .A1(n1389), .A2(key_out_24), .B1(n1388), .B2(key_out_23), .O(
        n1192) );
  XOR2X1 U971 ( .I1(n1191), .I2(n1193), .O(n1189) );
  OAI22X1 U972 ( .A1(n1388), .A2(n1389), .B1(key_out_23), .B2(key_out_24), .O(
        n1193) );
  OAI22X1 U973 ( .A1(n1375), .A2(n1194), .B1(n1195), .B2(n220), .O(n1191) );
  AOI22X1 U974 ( .A1(n1196), .A2(n1197), .B1(n840), .B2(n851), .O(n1195) );
  AOI22X1 U975 ( .A1(n1196), .A2(n840), .B1(n1197), .B2(n851), .O(n1194) );
  XOR4XLP U976 ( .I1(n801), .I2(n1198), .I3(n1384), .I4(n1199), .O(n2579gat)
         );
  OR2B1XLP U977 ( .I1(n1107), .B1(n1200), .O(n1199) );
  NR2X1 U978 ( .I1(n804), .I2(n802), .O(n1107) );
  XNR2X1 U979 ( .I1(n806), .I2(n800), .O(n1198) );
  NR2X1 U980 ( .I1(n874), .I2(n1021), .O(n2556gat) );
  XNR2X1 U981 ( .I1(n878), .I2(n1400), .O(n1021) );
  OR3X1 U982 ( .I1(n1201), .I2(n1202), .I3(n1203), .O(n878) );
  NR2X1 U983 ( .I1(n1168), .I2(n874), .O(n2539gat) );
  AN2X1 U984 ( .I1(n1204), .I2(n838), .O(n1168) );
  NR2X1 U985 ( .I1(n1027), .I2(n874), .O(n2436gat) );
  INVCKX1 U986 ( .I(n1205), .O(n1027) );
  OAI23X1 U987 ( .B1(n1201), .B2(n1202), .B3(n845), .A1(n1206), .A2(n1203), 
        .O(n1205) );
  XOR2X1 U988 ( .I1(n1366), .I2(key_14), .O(n1203) );
  AN2X1 U989 ( .I1(n1207), .I2(n846), .O(n1206) );
  INVCKX1 U990 ( .I(n1208), .O(n240) );
  NR2X1 U991 ( .I1(n1209), .I2(n1171), .O(n2396gat) );
  XNR2X1 U992 ( .I1(n836), .I2(n1210), .O(n1171) );
  NR2X1 U993 ( .I1(n1179), .I2(n874), .O(n2387gat) );
  OA22X1 U994 ( .A1(n1202), .A2(n846), .B1(n1207), .B2(n1201), .O(n1179) );
  XOR2X1 U995 ( .I1(n1397), .I2(key_38), .O(n1201) );
  XNR2X1 U996 ( .I1(n1207), .I2(key_36), .O(n1202) );
  NR2X1 U997 ( .I1(n877), .I2(n1204), .O(n1207) );
  NR2X1 U998 ( .I1(n1174), .I2(n874), .O(n2330gat) );
  ND2X1 U999 ( .I1(n914), .I2(n197), .O(n874) );
  AN3X1 U1000 ( .I1(n1211), .I2(n1212), .I3(n1213), .O(n914) );
  MXL2XLP U1001 ( .A(n1214), .B(n1215), .S(n1406), .OB(n1213) );
  NR2X1 U1002 ( .I1(n908), .I2(n1208), .O(n1215) );
  OAI112X1 U1003 ( .C1(n1357), .C2(n1358), .A1(n908), .B1(n1216), .O(n1212) );
  OR4B2XLP U1004 ( .I1(n1357), .I2(n1358), .B1(n814), .B2(n908), .O(n1211) );
  NR3X1 U1005 ( .I1(n1217), .I2(n1397), .I3(n845), .O(n814) );
  OA12X1 U1006 ( .B1(n853), .B2(n1204), .A1(n877), .O(n1174) );
  XOR2X1 U1007 ( .I1(n1398), .I2(key_27), .O(n877) );
  XOR2X1 U1008 ( .I1(n1399), .I2(key_26), .O(n1204) );
  INVCKX1 U1009 ( .I(n1196), .O(n221) );
  XOR2X1 U1010 ( .I1(n1386), .I2(key_29), .O(n1196) );
  XNR2X1 U1011 ( .I1(n1375), .I2(key_25), .O(n220) );
  NR2X1 U1012 ( .I1(n1170), .I2(n1209), .O(n2198gat) );
  NR2X1 U1013 ( .I1(n1209), .I2(n1032), .O(n2197gat) );
  XNR2X1 U1014 ( .I1(n881), .I2(n1365), .O(n1032) );
  NR2X1 U1015 ( .I1(n1209), .I2(n1031), .O(n2196gat) );
  ND2X1 U1016 ( .I1(n881), .I2(n1218), .O(n1031) );
  AO12X1 U1017 ( .B1(n836), .B2(n1210), .A1(n837), .O(n1218) );
  ND3X1 U1018 ( .I1(n837), .I2(n836), .I3(n1210), .O(n881) );
  NR2X1 U1019 ( .I1(n1176), .I2(n1219), .O(n2194gat) );
  AN2X1 U1020 ( .I1(n1407), .I2(n1376), .O(n1176) );
  AN4B2X1 U1021 ( .I1(n1220), .I2(n1364), .B1(n1221), .B2(n1359), .O(n2163gat)
         );
  NR2X1 U1022 ( .I1(n1219), .I2(n1175), .O(n2057gat) );
  XOR2X1 U1023 ( .I1(n1360), .I2(n1222), .O(n1175) );
  NR2X1 U1024 ( .I1(n1407), .I2(n1376), .O(n1222) );
  NR3X1 U1025 ( .I1(n2040gat), .I2(n1361), .I3(n1408), .O(n2015gat) );
  AOI112X1 U1026 ( .C1(n1408), .C2(n854), .A1(n1223), .B1(n1224), .O(n2009gat)
         );
  INVCKX1 U1027 ( .I(n2017gat), .O(n1223) );
  NR2X1 U1028 ( .I1(n902), .I2(n1221), .O(n2017gat) );
  INVCKX1 U1029 ( .I(n1209), .O(n196) );
  ND2X1 U1030 ( .I1(n197), .I2(n913), .O(n1209) );
  MXL2XLP U1031 ( .A(n1225), .B(n1226), .S(n908), .OB(n913) );
  AN4B2X1 U1032 ( .I1(n837), .I2(n847), .B1(n1403), .B2(n1227), .O(n1226) );
  ND2X1 U1033 ( .I1(n1401), .I2(n1402), .O(n1227) );
  NR2X1 U1034 ( .I1(n1221), .I2(n1228), .O(n1927gat) );
  INVCKX1 U1035 ( .I(n885), .O(n192) );
  NR2X1 U1036 ( .I1(n1208), .I2(n1229), .O(n1915gat) );
  ND2X1 U1037 ( .I1(n1230), .I2(n845), .O(n1208) );
  INVCKX1 U1038 ( .I(n883), .O(n191) );
  INVCKX1 U1039 ( .I(n884), .O(n189) );
  NR2X1 U1040 ( .I1(n778), .I2(n783), .O(n884) );
  ND2X1 U1041 ( .I1(n1231), .I2(n898), .O(n778) );
  INVCKX1 U1042 ( .I(n920), .O(n898) );
  AN4B2X1 U1043 ( .I1(n1053), .I2(n1143), .B1(n1232), .B2(n1409), .O(n920) );
  AN3B2X1 U1044 ( .I1(n1233), .B1(n711), .B2(n1362), .O(n1882gat) );
  NR2X1 U1045 ( .I1(n3099gat), .I2(n775), .O(n1827gat) );
  NR2X1 U1046 ( .I1(n1228), .I2(n1229), .O(n1800gat) );
  OR4B2XLP U1047 ( .I1(n1404), .I2(n1234), .B1(n836), .B2(n839), .O(n1229) );
  ND2X1 U1048 ( .I1(n1365), .I2(n1402), .O(n1234) );
  NR2X1 U1049 ( .I1(n1235), .I2(n1236), .O(n1793gat) );
  AN2B1XLP U1050 ( .I1(n888), .B1(n889), .O(n3107gat) );
  AN2X1 U1051 ( .I1(n1408), .I2(n1771gat), .O(n889) );
  AN4B1XLP U1052 ( .I1(n1237), .I2(n1238), .I3(n783), .B1(n840), .O(n3138gat)
         );
  NR2X1 U1053 ( .I1(n885), .I2(n1239), .O(n1696gat) );
  ND3X1 U1054 ( .I1(n1046), .I2(n1053), .I3(n1240), .O(n885) );
  AN4B1XLP U1055 ( .I1(n1397), .I2(n845), .I3(n2989gat), .B1(n1217), .O(
        n1636gat) );
  NR2X1 U1056 ( .I1(n1241), .I2(n1242), .O(n1620gat) );
  NR2X1 U1057 ( .I1(n1239), .I2(n883), .O(n1613gat) );
  ND3X1 U1058 ( .I1(n1053), .I2(n1241), .I3(n1240), .O(n883) );
  AN2B1XLP U1059 ( .I1(n1606gat), .B1(n1239), .O(n1610gat) );
  OR3B2X1 U1060 ( .I1(n901), .B1(n1233), .B2(n1363), .O(n1239) );
  AN2B1XLP U1061 ( .I1(n690), .B1(n788), .O(n901) );
  ND2X1 U1062 ( .I1(n1379), .I2(n1821gat), .O(n788) );
  AN2B1XLP U1063 ( .I1(n1146), .B1(n1409), .O(n1606gat) );
  XNR2X1 U1064 ( .I1(n271gat), .I2(key_79), .O(n1146) );
  NR3X1 U1065 ( .I1(n854), .I2(n1217), .I3(n1244), .O(n1593gat) );
  INVCKX1 U1066 ( .I(n1245), .O(n1217) );
  AN2B1XLP U1067 ( .I1(n813), .B1(n1236), .O(n1567gat) );
  AN4B2X1 U1068 ( .I1(n1398), .I2(n1400), .B1(n1397), .B2(n1246), .O(n813) );
  ND2X1 U1069 ( .I1(n1399), .I2(n1366), .O(n1246) );
  NR3X1 U1070 ( .I1(n1236), .I2(n1399), .I3(n873), .O(n1565gat) );
  OR3X1 U1071 ( .I1(n1244), .I2(n842), .I3(n1398), .O(n873) );
  OR4B2XLP U1072 ( .I1(n1404), .I2(n1247), .B1(n836), .B2(n848), .O(n1236) );
  ND2X1 U1073 ( .I1(n1365), .I2(n1403), .O(n1247) );
  NR3X1 U1074 ( .I1(n1248), .I2(n1221), .I3(n1225), .O(n1564gat) );
  AN4B2X1 U1075 ( .I1(n837), .I2(n847), .B1(n839), .B2(n882), .O(n1225) );
  ND2X1 U1076 ( .I1(n1401), .I2(n848), .O(n882) );
  AN4B1XLP U1077 ( .I1(n1249), .I2(n847), .I3(n3149gat), .B1(n1235), .O(n1221)
         );
  AOI12X1 U1078 ( .B1(n908), .B2(n1216), .A1(n1214), .O(n1235) );
  INVCKX1 U1079 ( .I(n1248), .O(n1214) );
  INVCKX1 U1080 ( .I(n1228), .O(n1216) );
  ND2X1 U1081 ( .I1(n1230), .I2(n1366), .O(n1228) );
  AN4B1XLP U1082 ( .I1(n838), .I2(n846), .I3(n1400), .B1(n1398), .O(n1230) );
  INVCKX1 U1083 ( .I(n2989gat), .O(n908) );
  ND3X1 U1084 ( .I1(n1834gat), .I2(n1767gat), .I3(n1390), .O(n3149gat) );
  MXL2XLP U1085 ( .A(n1250), .B(n1251), .S(n836), .OB(n1249) );
  OAI112X1 U1086 ( .C1(n1252), .C2(n1253), .A1(n1066), .B1(n1404), .O(n1251)
         );
  OR2X1 U1087 ( .I1(n1254), .I2(n1255), .O(n1253) );
  MXL2XLP U1088 ( .A(n1256), .B(n1170), .S(n837), .OB(n1250) );
  NR2X1 U1089 ( .I1(n1066), .I2(n1257), .O(n1256) );
  AOI112X1 U1090 ( .C1(n1254), .C2(n949), .A1(n1252), .B1(n1255), .O(n1257) );
  AN3X1 U1091 ( .I1(n1258), .I2(n1210), .I3(n1259), .O(n1255) );
  NR2X1 U1092 ( .I1(n1402), .I2(n1403), .O(n1210) );
  MUX2X1 U1093 ( .A(n1260), .B(n1261), .S(n1402), .O(n1252) );
  AN3B2X1 U1094 ( .I1(n1258), .B1(n1403), .B2(n1259), .O(n1261) );
  NR3X1 U1095 ( .I1(n1262), .I2(n1258), .I3(n839), .O(n1260) );
  NR3X1 U1096 ( .I1(n1258), .I2(n1259), .I3(n1263), .O(n1254) );
  INVCKX1 U1097 ( .I(n1262), .O(n1259) );
  ND2X1 U1098 ( .I1(n949), .I2(n940), .O(n1262) );
  XNR2X1 U1099 ( .I1(n846gat), .I2(key_95), .O(n940) );
  INVCKX1 U1100 ( .I(n1264), .O(n949) );
  NR2X1 U1101 ( .I1(n1264), .I2(n943), .O(n1258) );
  XOR2X1 U1102 ( .I1(n919gat), .I2(key_97), .O(n943) );
  NR2X1 U1103 ( .I1(n1264), .I2(n955), .O(n1066) );
  XOR2X1 U1104 ( .I1(n402gat), .I2(key_100), .O(n955) );
  XNR2X1 U1105 ( .I1(n398gat), .I2(key_101), .O(n1264) );
  ND2X1 U1106 ( .I1(n1265), .I2(n2989gat), .O(n1248) );
  OAI12X1 U1107 ( .B1(n1390), .B2(n1763gat), .A1(n2102gat), .O(n2989gat) );
  XOR2X1 U1108 ( .I1(key_30), .I2(n1266), .O(n1265) );
  AN4B1XLP U1109 ( .I1(n1398), .I2(n842), .I3(n838), .B1(n1244), .O(n1266) );
  AN4B1XLP U1110 ( .I1(n847), .I2(n1267), .I3(n1245), .B1(n1244), .O(n1516gat)
         );
  ND2X1 U1111 ( .I1(n1397), .I2(n1366), .O(n1244) );
  NR3X1 U1112 ( .I1(n842), .I2(n1399), .I3(n853), .O(n1245) );
  NR3X1 U1113 ( .I1(n1263), .I2(n836), .I3(n837), .O(n1267) );
  INVCKX1 U1114 ( .I(n1170), .O(n1263) );
  NR2X1 U1115 ( .I1(n839), .I2(n848), .O(n1170) );
  AN4B2X1 U1116 ( .I1(n1090), .I2(n804), .B1(n802), .B2(n1268), .O(n1391gat)
         );
  ND2X1 U1117 ( .I1(n1237), .I2(n1387), .O(n1268) );
  NR2X1 U1118 ( .I1(n1102), .I2(n803), .O(n1090) );
  XOR4XLP U1119 ( .I1(n1371), .I2(n1269), .I3(n861), .I4(n1270), .O(n3116gat)
         );
  XOR4XLP U1120 ( .I1(n1369), .I2(n1370), .I3(n1367), .I4(n1368), .O(n1270) );
  AOI12X1 U1121 ( .B1(n1392), .B2(key_22), .A1(n1271), .O(n1269) );
  MXL2XLP U1122 ( .A(n1272), .B(n1273), .S(n841), .OB(n1271) );
  OR2B1XLP U1123 ( .I1(key_22), .B1(n1272), .O(n1273) );
  NR2X1 U1124 ( .I1(n1392), .I2(key_21), .O(n1272) );
  XOR2X1 U1125 ( .I1(n1274), .I2(key_90), .O(key_out_90) );
  OAI22X1 U1126 ( .A1(n998), .A2(n1275), .B1(n1276), .B2(n1007), .O(n1274) );
  XOR2X1 U1127 ( .I1(key_9), .I2(n1277), .O(key_out_9) );
  XOR2X1 U1128 ( .I1(n1278), .I2(key_89), .O(key_out_89) );
  OAI22X1 U1129 ( .A1(n993), .A2(n1275), .B1(n1276), .B2(n995), .O(n1278) );
  XOR2X1 U1130 ( .I1(n1279), .I2(key_88), .O(key_out_88) );
  OAI22X1 U1131 ( .A1(n1010), .A2(n1275), .B1(n1276), .B2(n1009), .O(n1279) );
  XOR2X1 U1132 ( .I1(n1280), .I2(key_85), .O(key_out_85) );
  OAI22X1 U1133 ( .A1(n973), .A2(n1275), .B1(n1276), .B2(n980), .O(n1280) );
  XOR2X1 U1134 ( .I1(n1281), .I2(key_84), .O(key_out_84) );
  OAI22X1 U1135 ( .A1(n1002), .A2(n1275), .B1(n1276), .B2(n1004), .O(n1281) );
  XOR2X1 U1136 ( .I1(n1282), .I2(key_83), .O(key_out_83) );
  OAI22X1 U1137 ( .A1(n983), .A2(n1275), .B1(n1276), .B2(n1001), .O(n1282) );
  XOR2X1 U1138 ( .I1(n1283), .I2(key_82), .O(key_out_82) );
  OAI22X1 U1139 ( .A1(n991), .A2(n1275), .B1(n1276), .B2(n990), .O(n1283) );
  XOR2X1 U1140 ( .I1(n1284), .I2(key_81), .O(key_out_81) );
  OAI22X1 U1141 ( .A1(n986), .A2(n1275), .B1(n1276), .B2(n997), .O(n1284) );
  XOR2X1 U1142 ( .I1(key_8), .I2(n1285), .O(key_out_8) );
  XOR2X1 U1143 ( .I1(key_7), .I2(n1286), .O(key_out_7) );
  XOR2X1 U1144 ( .I1(key_6), .I2(n1287), .O(key_out_6) );
  XOR2X1 U1145 ( .I1(key_5), .I2(n1288), .O(key_out_5) );
  INVCKX1 U1146 ( .I(n906), .O(key_out_46) );
  XOR2X1 U1147 ( .I1(n1405), .I2(key_46), .O(n906) );
  XOR2X1 U1148 ( .I1(key_4), .I2(n1289), .O(key_out_4) );
  INVCKX1 U1149 ( .I(n1197), .O(key_out_37) );
  XOR2X1 U1150 ( .I1(n1387), .I2(key_37), .O(n1197) );
  XNR2X1 U1151 ( .I1(n1388), .I2(key_24), .O(key_out_24) );
  INVCKX1 U1152 ( .I(n1187), .O(key_out_20) );
  XOR2X1 U1153 ( .I1(n1427), .I2(key_20), .O(n1187) );
  XNR2X1 U1154 ( .I1(n1373), .I2(key_19), .O(key_out_19) );
  XNR2X1 U1155 ( .I1(n1374), .I2(key_18), .O(key_out_18) );
  XOR2X1 U1156 ( .I1(n1290), .I2(key_17), .O(key_out_17) );
  OAI22X1 U1157 ( .A1(n966), .A2(n1275), .B1(n1276), .B2(n971), .O(n1290) );
  XNR2X1 U1158 ( .I1(n3095gat), .I2(key_2), .O(n1276) );
  XNR2X1 U1159 ( .I1(n3093gat), .I2(key_15), .O(n1275) );
  XOR2X1 U1160 ( .I1(n1291), .I2(key_128), .O(key_out_128) );
  OAI12X1 U1161 ( .B1(n993), .B2(n999), .A1(n1000), .O(n1291) );
  XOR2X1 U1162 ( .I1(n1292), .I2(key_127), .O(key_out_127) );
  OAI12X1 U1163 ( .B1(n1010), .B2(n999), .A1(n1000), .O(n1292) );
  XOR2X1 U1164 ( .I1(n1293), .I2(key_126), .O(key_out_126) );
  OAI12X1 U1165 ( .B1(n966), .B2(n999), .A1(n1000), .O(n1293) );
  XOR2X1 U1166 ( .I1(n1294), .I2(key_125), .O(key_out_125) );
  OAI12X1 U1167 ( .B1(n1002), .B2(n999), .A1(n1000), .O(n1294) );
  XOR2X1 U1168 ( .I1(n1295), .I2(key_124), .O(key_out_124) );
  OAI12X1 U1169 ( .B1(n983), .B2(n999), .A1(n1000), .O(n1295) );
  XOR2X1 U1170 ( .I1(n1296), .I2(key_123), .O(key_out_123) );
  OAI12X1 U1171 ( .B1(n991), .B2(n999), .A1(n1000), .O(n1296) );
  XOR2X1 U1172 ( .I1(n1297), .I2(key_122), .O(key_out_122) );
  OAI12X1 U1173 ( .B1(n986), .B2(n999), .A1(n1000), .O(n1297) );
  XNR2X1 U1174 ( .I1(n1298), .I2(key_1), .O(n999) );
  OAI23X1 U1175 ( .B1(n1299), .B2(n1011), .B3(n1169), .A1(n1029), .A2(n1025), 
        .O(n1298) );
  ND2X1 U1176 ( .I1(n868), .I2(n1016), .O(n1025) );
  ND2X1 U1177 ( .I1(n1300), .I2(n1012), .O(n1016) );
  XNR2X1 U1178 ( .I1(n1015), .I2(key_28), .O(n868) );
  ND2X1 U1179 ( .I1(n1300), .I2(n1150), .O(n1015) );
  ND2X1 U1180 ( .I1(n3094gat), .I2(n1172), .O(n1029) );
  INVCKX1 U1181 ( .I(n1022), .O(n1172) );
  ND2X1 U1182 ( .I1(n1300), .I2(n871), .O(n1022) );
  XNR2X1 U1183 ( .I1(n1301), .I2(key_63), .O(n1300) );
  ND3X1 U1184 ( .I1(n1017), .I2(n1162), .I3(n1156), .O(n1301) );
  INVCKX1 U1185 ( .I(n965), .O(n1156) );
  OR4B2XLP U1186 ( .I1(n1150), .I2(n1164), .B1(n1012), .B2(n1017), .O(n1169)
         );
  AN2X1 U1187 ( .I1(n962), .I2(n888), .O(n1017) );
  XNR2X1 U1188 ( .I1(n3106gat), .I2(key_33), .O(n888) );
  NR2X1 U1189 ( .I1(n1157), .I2(n1158), .O(n962) );
  XOR2X1 U1190 ( .I1(n3084gat), .I2(key_66), .O(n1158) );
  XOR2X1 U1191 ( .I1(n3083gat), .I2(key_69), .O(n1157) );
  XOR2X1 U1192 ( .I1(n3088gat), .I2(key_71), .O(n1012) );
  INVCKX1 U1193 ( .I(n1163), .O(n1164) );
  XOR2X1 U1194 ( .I1(n3087gat), .I2(key_68), .O(n1150) );
  INVCKX1 U1195 ( .I(n871), .O(n1011) );
  XOR2X1 U1196 ( .I1(n3086gat), .I2(key_70), .O(n871) );
  ND2X1 U1197 ( .I1(n965), .I2(n1018), .O(n1299) );
  OR2X1 U1198 ( .I1(n3092gat), .I2(n3091gat), .O(n1018) );
  XOR2X1 U1199 ( .I1(n3085gat), .I2(key_67), .O(n965) );
  XOR2X1 U1200 ( .I1(key_12), .I2(n1302), .O(key_out_12) );
  XOR2X1 U1201 ( .I1(n1303), .I2(key_119), .O(key_out_119) );
  OAI122X1 U1202 ( .B1(n998), .B2(n1304), .C1(n1305), .C2(n1007), .A1(n1000), 
        .O(n1303) );
  INVCKX1 U1203 ( .I(n3078gat), .O(n1007) );
  XNR2X1 U1204 ( .I1(n1289), .I2(key_56), .O(n998) );
  XOR2X1 U1205 ( .I1(n3069gat), .I2(key_57), .O(n1289) );
  XOR2X1 U1206 ( .I1(n1306), .I2(key_118), .O(key_out_118) );
  OAI122X1 U1207 ( .B1(n993), .B2(n1304), .C1(n1305), .C2(n995), .A1(n1000), 
        .O(n1306) );
  INVCKX1 U1208 ( .I(n3079gat), .O(n995) );
  XNR2X1 U1209 ( .I1(n1287), .I2(key_52), .O(n993) );
  XOR2X1 U1210 ( .I1(n3070gat), .I2(key_59), .O(n1287) );
  XOR2X1 U1211 ( .I1(n1307), .I2(key_117), .O(key_out_117) );
  OAI122X1 U1212 ( .B1(n1010), .B2(n1304), .C1(n1305), .C2(n1009), .A1(n1000), 
        .O(n1307) );
  INVCKX1 U1213 ( .I(n3077gat), .O(n1009) );
  XNR2X1 U1214 ( .I1(n1302), .I2(key_51), .O(n1010) );
  XOR2X1 U1215 ( .I1(n3068gat), .I2(key_64), .O(n1302) );
  XOR2X1 U1216 ( .I1(n1308), .I2(key_115), .O(key_out_115) );
  OAI122X1 U1217 ( .B1(n966), .B2(n1304), .C1(n1305), .C2(n971), .A1(n1000), 
        .O(n1308) );
  INVCKX1 U1218 ( .I(n3081gat), .O(n971) );
  XNR2X1 U1219 ( .I1(n1288), .I2(key_53), .O(n966) );
  XOR2X1 U1220 ( .I1(n3072gat), .I2(key_58), .O(n1288) );
  XOR2X1 U1221 ( .I1(n1309), .I2(key_114), .O(key_out_114) );
  OAI122X1 U1222 ( .B1(n1002), .B2(n1304), .C1(n1305), .C2(n1004), .A1(n1000), 
        .O(n1309) );
  INVCKX1 U1223 ( .I(n3080gat), .O(n1004) );
  XNR2X1 U1224 ( .I1(n1286), .I2(key_54), .O(n1002) );
  XOR2X1 U1225 ( .I1(n3071gat), .I2(key_62), .O(n1286) );
  XOR2X1 U1226 ( .I1(n1310), .I2(key_112), .O(key_out_112) );
  OAI122X1 U1227 ( .B1(n983), .B2(n1304), .C1(n1305), .C2(n1001), .A1(n1000), 
        .O(n1310) );
  INVCKX1 U1228 ( .I(n3075gat), .O(n1001) );
  XNR2X1 U1229 ( .I1(n1311), .I2(key_49), .O(n983) );
  XOR2X1 U1230 ( .I1(n1312), .I2(key_111), .O(key_out_111) );
  OAI122X1 U1231 ( .B1(n991), .B2(n1304), .C1(n1305), .C2(n990), .A1(n1000), 
        .O(n1312) );
  INVCKX1 U1232 ( .I(n3076gat), .O(n990) );
  XNR2X1 U1233 ( .I1(n1277), .I2(key_48), .O(n991) );
  XOR2X1 U1234 ( .I1(n3067gat), .I2(key_65), .O(n1277) );
  XOR2X1 U1235 ( .I1(n1313), .I2(key_110), .O(key_out_110) );
  OAI122X1 U1236 ( .B1(n986), .B2(n1304), .C1(n1305), .C2(n997), .A1(n1000), 
        .O(n1313) );
  INVCKX1 U1237 ( .I(n3074gat), .O(n997) );
  XNR2X1 U1238 ( .I1(n1285), .I2(key_50), .O(n986) );
  XOR2X1 U1239 ( .I1(n3065gat), .I2(key_60), .O(n1285) );
  XOR2X1 U1240 ( .I1(key_11), .I2(n1314), .O(key_out_11) );
  XOR2X1 U1241 ( .I1(n1315), .I2(key_108), .O(key_out_108) );
  OAI122X1 U1242 ( .B1(n1305), .B2(n980), .C1(n973), .C2(n1304), .A1(n1000), 
        .O(n1315) );
  XOR2X1 U1243 ( .I1(n1316), .I2(key_120), .O(n1000) );
  OR4B2XLP U1244 ( .I1(n1385), .I2(n895), .B1(n840), .B2(n1317), .O(n1316) );
  NR3X1 U1245 ( .I1(n1318), .I2(n909), .I3(n1238), .O(n1317) );
  NR3X1 U1246 ( .I1(n1200), .I2(n1384), .I3(n1102), .O(n1238) );
  INVCKX1 U1247 ( .I(n1130), .O(n1102) );
  NR2X1 U1248 ( .I1(n801), .I2(n800), .O(n1130) );
  NR3X1 U1249 ( .I1(n1105), .I2(n1200), .I3(n803), .O(n909) );
  ND2X1 U1250 ( .I1(n802), .I2(n804), .O(n1200) );
  INVCKX1 U1251 ( .I(n1100), .O(n1105) );
  NR2X1 U1252 ( .I1(n800), .I2(n1383), .O(n1100) );
  MXL2XLP U1253 ( .A(n1319), .B(n1237), .S(n1391), .OB(n1318) );
  AN4B2X1 U1254 ( .I1(n1388), .I2(n1389), .B1(n851), .B2(n1375), .O(n1237) );
  AN4B1XLP U1255 ( .I1(n1375), .I2(n1388), .I3(key_out_23), .B1(n1386), .O(
        n1319) );
  XNR2X1 U1256 ( .I1(n1389), .I2(key_23), .O(key_out_23) );
  INVCKX1 U1257 ( .I(n780), .O(n895) );
  OR2B1XLP U1258 ( .I1(n783), .B1(n1231), .O(n780) );
  OA13X1 U1259 ( .B1(n1242), .B2(n1409), .B3(n1046), .A1(n1115), .O(n1231) );
  OR4B2XLP U1260 ( .I1(n1232), .I2(n1241), .B1(n1142), .B2(n1320), .O(n1115)
         );
  NR2X1 U1261 ( .I1(n1409), .I2(n1143), .O(n1320) );
  ND3X1 U1262 ( .I1(n1143), .I2(n1142), .I3(n1057), .O(n1242) );
  INVCKX1 U1263 ( .I(n1062), .O(n1143) );
  ND2X1 U1264 ( .I1(n978), .I2(n972), .O(n783) );
  ND3X1 U1265 ( .I1(n1046), .I2(n1142), .I3(n1240), .O(n972) );
  INVCKX1 U1266 ( .I(n1241), .O(n1046) );
  ND3X1 U1267 ( .I1(n1142), .I2(n1241), .I3(n1240), .O(n978) );
  NR3X1 U1268 ( .I1(n1057), .I2(n1409), .I3(n1062), .O(n1240) );
  XNR2X1 U1269 ( .I1(n394gat), .I2(key_75), .O(n1062) );
  INVCKX1 U1270 ( .I(n1232), .O(n1057) );
  XNR2X1 U1271 ( .I1(n703gat), .I2(key_77), .O(n1232) );
  XNR2X1 U1272 ( .I1(n722gat), .I2(key_76), .O(n1241) );
  INVCKX1 U1273 ( .I(n1053), .O(n1142) );
  XNR2X1 U1274 ( .I1(n726gat), .I2(key_78), .O(n1053) );
  XNR2X1 U1275 ( .I1(n1163), .I2(key_16), .O(n1304) );
  XOR2X1 U1276 ( .I1(n3093gat), .I2(key_40), .O(n1163) );
  XNR2X1 U1277 ( .I1(n1314), .I2(key_47), .O(n973) );
  XOR2X1 U1278 ( .I1(n3073gat), .I2(key_55), .O(n1314) );
  INVCKX1 U1279 ( .I(n3082gat), .O(n980) );
  XNR2X1 U1280 ( .I1(n1162), .I2(key_3), .O(n1305) );
  XOR2X1 U1281 ( .I1(n3095gat), .I2(key_35), .O(n1162) );
  XOR2X1 U1282 ( .I1(n1321), .I2(key_106), .O(key_out_106) );
  ND2X1 U1283 ( .I1(n197), .I2(n1322), .O(n1321) );
  XOR2X1 U1284 ( .I1(n2266gat), .I2(n1323), .O(n1322) );
  ND2X1 U1285 ( .I1(n1407), .I2(n855), .O(n1323) );
  INVCKX1 U1286 ( .I(n1219), .O(n197) );
  OAI112X1 U1287 ( .C1(n902), .C2(n712), .A1(n1324), .B1(n1325), .O(n1219) );
  AN2X1 U1288 ( .I1(n1410), .I2(n1220), .O(n1325) );
  INVCKX1 U1289 ( .I(n1224), .O(n1220) );
  XNR2X1 U1290 ( .I1(n1326), .I2(key_31), .O(n1224) );
  XNR2X1 U1291 ( .I1(n3100gat), .I2(key_39), .O(n1243) );
  OR4B2XLP U1292 ( .I1(n733), .I2(n776), .B1(n1327), .B2(n1378), .O(n784) );
  NR2X1 U1293 ( .I1(n1377), .I2(n731), .O(n1327) );
  INVCKX1 U1294 ( .I(key_out_32), .O(n1324) );
  XNR2X1 U1295 ( .I1(n2095gat), .I2(key_32), .O(key_out_32) );
  AN2X1 U1296 ( .I1(n1390), .I2(n2021gat), .O(n902) );
  XOR2X1 U1297 ( .I1(key_10), .I2(n1311), .O(key_out_10) );
  XOR2X1 U1298 ( .I1(n3066gat), .I2(key_61), .O(n1311) );
endmodule

