module s13207(clk, g43, g49, g633, g634, g635, g645, g647, g648, g690, g694, g698, g702, g722, g723, g751, g752, g753, g754, g755, g756, g757, g781, g941, g962, g1000, g1008, g1016, g1080, g1234, g1553, g1554, g786, g1206, g929, g955, g795, g1194, g1198, g1202, g24, g1203, g1196, g29, g22, g28, g10, g23, g37, g26, g1, g27, g42, g11, g32, g41, g31, g45, g9, g44, g21, g30, g25, g206, g291, g372, g453, g534, g594, g785, g1006, g1015, g1017, g1246, g1724, g1783, g1798, g1804, g1810, g1817, g1824, g1829, g1870, g1871, g1894, g1911, g1944, g2662, g2844, g2888, g3077, g3096, g3130, g3159, g3191, g3829, g3859, g3860, g4267, g4316, g4370, g4371, g4372, g4373, g4655, g4657, g4660, g4661, g4663, g4664, g5143, g5164, g5571, g5669, g5678, g5682, g5684, g5687, g5729, g6207, g6212, g6223, g6236, g6269, g6425, g6648, g6653, g6675, g6849, g6850, g6895, g6909, g7048, g7063, g7103, g7283, g7284, g7285, g7286, g7287, g7288, g7289, g7290, g7291, g7292, g7293, g7294, g7295, g7298, g7423, g7424, g7425, g7474, g7504, g7505, g7506, g7507, g7508, g7514, g7729, g7730, g7731, g7732, g8216, g8217, g8218, g8219, g8234, g8661, g8663, g8872, g8958, g9128, g9132, g9204, g9280, g9297, g9299, g9305, g9308, g9310, g9312, g9314, g9378, g7763, g1205, g3856, g3857, g3854, g1193, g1197, g1201, g6294, g6376, g1195, g6300, g6292, g6298, g6291, g6293, g6304, g6296, g6289, g6297, g6306, g6290, g6303, g6305, g6302, g6308, g6288, g6307, g6299, g6301, g6295);
input clk, g43, g49, g633, g634, g635, g645, g647, g648, g690, g694, g698, g702, g722, g723, g751, g752, g753, g754, g755, g756, g757, g781, g941, g962, g1000, g1008, g1016, g1080, g1234, g1553, g1554, g786, g1206, g929, g955, g795, g1194, g1198, g1202, g24, g1203, g1196, g29, g22, g28, g10, g23, g37, g26, g1, g27, g42, g11, g32, g41, g31, g45, g9, g44, g21, g30, g25;
output g206, g291, g372, g453, g534, g594, g785, g1006, g1015, g1017, g1246, g1724, g1783, g1798, g1804, g1810, g1817, g1824, g1829, g1870, g1871, g1894, g1911, g1944, g2662, g2844, g2888, g3077, g3096, g3130, g3159, g3191, g3829, g3859, g3860, g4267, g4316, g4370, g4371, g4372, g4373, g4655, g4657, g4660, g4661, g4663, g4664, g5143, g5164, g5571, g5669, g5678, g5682, g5684, g5687, g5729, g6207, g6212, g6223, g6236, g6269, g6425, g6648, g6653, g6675, g6849, g6850, g6895, g6909, g7048, g7063, g7103, g7283, g7284, g7285, g7286, g7287, g7288, g7289, g7290, g7291, g7292, g7293, g7294, g7295, g7298, g7423, g7424, g7425, g7474, g7504, g7505, g7506, g7507, g7508, g7514, g7729, g7730, g7731, g7732, g8216, g8217, g8218, g8219, g8234, g8661, g8663, g8872, g8958, g9128, g9132, g9204, g9280, g9297, g9299, g9305, g9308, g9310, g9312, g9314, g9378, g7763, g1205, g3856, g3857, g3854, g1193, g1197, g1201, g6294, g6376, g1195, g6300, g6292, g6298, g6291, g6293, g6304, g6296, g6289, g6297, g6306, g6290, g6303, g6305, g6302, g6308, g6288, g6307, g6299, g6301, g6295;
wire clk, g43, g49, g633, g634, g635, g645, g647, g648, g690, g694, g698, g702, g722, g723, g751, g752, g753, g754, g755, g756, g757, g781, g941, g962, g1000, g1008, g1016, g1080, g1234, g1553, g1554, g786, g1206, g929, g955, g795, g1194, g1198, g1202, g24, g1203, g1196, g29, g22, g28, g10, g23, g37, g26, g1, g27, g42, g11, g32, g41, g31, g45, g9, g44, g21, g30, g25;
wire g397, g1271, g312, g273, g452, g948, g629, g207, g1541, g1153, g940;
wire g976, g498, g314, g1092, g454, g196, g535, g292, g772, g1375, g689;
wire g183, g359, g1384, g1339, g20, g1424, g767, g393, g1077, g1231, g294;
wire g1477, g4, g608, g1205, g465, g774, g921, g1304, g243, g1499, g80;
wire g1444, g1269, g600, g423, g771, g803, g843, g315, g455, g906, g622;
wire g891, g1014, g984, g117, g137, g527, g1513, g278, g1378, g718, g598;
wire g1182, g1288, g1382, g179, g624, g48, g362, g878, g270, g763, g710;
wire g730, g295, g1037, g1102, g483, g775, g621, g1364, g1454, g1296, g5;
wire g1532, g587, g741, g13, g606, g1012, g52, g646, g1412, g327, g1189;
wire g1389, g1029, g1371, g1429, g398, g985, g354, g619, g113, g133, g180;
wire g1138, g1309, g889, g390, g625, g417, g681, g437, g351, g1201, g109;
wire g1049, g1098, g200, g240, g479, g126, g596, g1268, g222, g420, g3;
wire g58, g172, g387, g840, g365, g1486, g1504, g1185, g1385, g583, g822;
wire g1025, g969, g768, g174, g685, g1087, g355, g911, g1226, g99, g1045;
wire g1173, g1373, g186, g760, g959, g1369, g1007, g1459, g758, g480, g396;
wire g612, g38, g632, g1415, g1227, g246, g449, g517, g118, g138, g16;
wire g284, g142, g219, g426, g1388, g806, g846, g1428, g579, g1030, g614;
wire g1430, g1247, g669, g110, g130, g225, g281, g819, g1308, g611, g631;
wire g1217, g104, g1365, g825, g1333, g474, g1396, g141, g1509, g766, g1018;
wire g588, g1467, g317, g457, g486, g471, g1381, g1197, g513, g1397, g533;
wire g1021, g1421, g952, g1263, g580, g615, g1257, g46, g402, g998, g1041;
wire g297, g954, g105, g145, g212, g1368, g232, g990, g475, g33, g951;
wire g799, g812, g567, g313, g333, g168, g214, g234, g652, g1126, g1400;
wire g1326, g92, g309, g211, g834, g231, g557, g1383, g1220, g158, g627;
wire g661, g77, g831, g1327, g293, g1146, g89, g150, g773, g859, g1240;
wire g518, g1472, g1443, g436, g405, g1034, g1147, g374, g98, g563, g510;
wire g530, g215, g235, g1013, g6, g55, g1317, g504, g665, g544, g371;
wire g62, g792, g468, g815, g1460, g553, g623, g501, g1190, g1390, g74;
wire g1156, g318, g458, g342, g1250, g1163, g1363, g1432, g1053, g252, g330;
wire g264, g1157, g1357, g375, g68, g852, g261, g516, g536, g979, g778;
wire g199, g1292, g290, g1084, g1439, g770, g1276, g890, g1004, g1404, g93;
wire g2, g287, g560, g1224, g1320, g617, g316, g336, g933, g456, g345;
wire g628, g8, g887, g789, g173, g550, g255, g949, g1244, g620, g1435;
wire g477, g926, g368, g855, g1214, g1110, g1310, g296, g972, g1402, g1236;
wire g896, g613, g566, g1394, g1489, g883, g47, g971, g609, g103, g1254;
wire g556, g1409, g626, g1229, g782, g237, g942, g228, g706, g746, g1462;
wire g963, g129, g837, g599, g1192, g828, g1392, g492, g95, g944, g195;
wire g1431, g1252, g356, g953, g1176, g1376, g1005, g1405, g901, g1270, g1225;
wire g1073, g1324, g1069, g443, g1377, g377, g618, g602, g213, g233, g1199;
wire g1399, g83, g888, g573, g399, g1245, g507, g547, g108, g610, g630;
wire g1207, g249, g65, g916, g936, g478, g604, g945, g1114, g100, g429;
wire g809, g849, g1408, g1336, g601, g122, g1065, g1122, g1228, g495, g1322;
wire g1230, g1033, g267, g1195, g1395, g373, g274, g1266, g714, g734, g1142;
wire g1342, g769, g1081, g1481, g1097, g543, g1154, g1354, g489, g874, g121;
wire g591, g616, g1267, g1312, g605, g182, g1401, g950, g1329, g408, g871;
wire g759, g146, g202, g440, g476, g184, g1149, g1398, g210, g394, g86;
wire g570, g275, g303, g125, g181, g1524, g595, g1319, g863, g1211, g966;
wire g1186, g1386, g875, g1170, g1370, g201, g1325, g1280, g1106, g1061, g1387;
wire g762, g1461, g378, g1200, g1514, g1403, g1345, g1191, g1391, g185, g1307;
wire g1159, g1223, g446, g1416, g395, g764, g1251, g216, g236, g205, g540;
wire g576, g1537, g727, g999, g761, g1272, g1243, g1328, g1130, g1330, g114;
wire g134, g1166, g524, g1366, g348, g1148, g1348, g1155, g1260, g7, g258;
wire g521, g300, g765, g1118, g1167, g1318, g1367, g677, g376, g1057, g973;
wire g1193, g1393, g1549, g1321, g1253, g1519, g584, g539, g324, g432, g1158;
wire g321, g1311, g414, g1374, g94, g1284, g1545, g1380, g673, g607, g306;
wire g943, g162, g411, g866, g1204, g1300, g384, g339, g459, g1323, g381;
wire g1528, g1351, g597, g1372, g154, g435, g970, g1134, g995, g190, g1313;
wire g603, g1494, g462, g1160, g1360, g1450, g187, g1179, g1379, g12, g71;
wire g1658, g1777, I9325, I7758, g5652, I13502, g6895, g3880, g6837, I15824, g5843;
wire I6112, g7189, g8970, I6267, g6062, I16126, I10519, I15181, I11443, I12436, I10675;
wire g2547, I7365, I10154, g1611, I11278, g7171, I14154, I12274, g8224, g5834, g5971;
wire g3978, I6676, g3612, I8520, g2892, I13469, I12346, I9636, I14637, g6788, g1799;
wire g3935, I5933, g9207, I13039, I15426, g5598, g1674, g7281, g3982, g4666, I15190;
wire g2945, g5121, g3128, g3629, g7297, g5670, I11815, g6842, g3130, g9088, g8789;
wire g3542, I12292, g6298, g2709, I11677, g6392, g4648, I8829, I15546, g1680, I15211;
wire g2340, I12409, g4655, g7745, g7138, I6703, g5938, g8771, g2478, g5813, g7338;
wire g2907, g1744, g9215, g7109, g6854, I12635, g7309, g1802, I10439, g2959, I14728;
wire I8733, I14439, g2517, g4010, I7662, I9446, I8974, g5740, g5519, g9114, g1558;
wire I7290, g2876, g9314, I11884, I9145, I6468, g5606, I8796, g7759, I14349, I11410;
wire I12164, g695, g6708, I13410, I15625, g6520, g1901, g6219, g6640, I8980, g3902;
wire I12891, I11479, I11666, g5687, g2915, I13666, g6252, g6812, g4372, g7049, g3512;
wire I13478, g5586, g6958, I15943, g4618, I6716, g6376, g4667, I5981, I8177, I7847;
wire I16055, g9336, g2310, g7715, g1600, g1574, g1864, g4566, I11556, g7098, I5997;
wire g6829, g7498, g2663, I12108, g6765, g3529, g8959, I6198, g4693, I13580, g4134;
wire g3649, I14139, I9416, I12283, g8482, g5525, g3851, g5645, I5353, g2402, I7950;
wire g2824, g1580, g2236, g7584, g4555, g9065, I9642, g7539, I15411, I15527, I10415;
wire I13084, g9322, g3964, g4792, g9230, g6225, I8781, I8898, g6073, g2877, g6796;
wire g1736, I12091, g4621, g5607, g9033, g7162, g7268, g7019, I11740, g7362, g5158;
wire I13740, I9654, I15894, g6324, I7723, g4113, g6069, g2556, g1889, I7101, I5901;
wire g2222, I13676, g9096, I8291, I13373, g2928, g4202, g8663, I7605, I15714, g5587;
wire g2930, I15315, I11800, g1871, g4908, g6377, g6206, g5311, g2899, g9195, g4094;
wire I11936, g3872, I15202, g3652, g4567, g7728, g7486, g3843, g3989, I6186, g7730;
wire I9612, I10608, g5174, g8762, g7504, I15978, I14115, g7185, g4776, I7041, g6849;
wire I9935, g4593, I11964, g3549, g3834, g3971, g7070, g2295, I14052, g2237, g7470;
wire I15741, g8657, g6781, g7425, g5180, g2844, I8215, g6898, g1838, g5591, g6900;
wire g8222, I8886, g5832, I14813, g1795, g6797, g1737, g2394, g9248, g1809, I10973;
wire I14798, g6245, g4360, I7368, g9255, g9081, I12948, I13909, I15735, g4521, I14184;
wire g1672, I14674, g8464, g6291, I12702, g2557, g4050, g4641, I11908, I12757, g9097;
wire g2966, g5794, I5889, g1643, I11569, g7131, g6344, g2471, g7006, g7331, I15196;
wire I6636, I14732, g2242, g6207, g3909, I11747, I12564, g8563, g2948, I11242, g7766;
wire g6819, g7105, g3519, I10761, g7305, I7856, I7734, g2955, g7487, g5628, g1742;
wire g6088, g6852, g5515, I12397, g6488, g4658, g7748, g4777, I10400, g5100, I9512;
wire I13807, I11974, I12062, I14400, g2350, g9112, g7755, g9218, g1926, I9823, g9312;
wire g2038, g4882, I14214, I12933, I9366, g7226, I11230, I11293, I10207, I13293, I12508;
wire I11638, g6886, I6446, g4611, g291, I14005, g7045, I11416, I10538, I6003, I9148;
wire I13416, I5795, g9129, g2769, g7173, g9329, g6314, g7091, g7491, g6870, g3860;
wire g2918, g3341, g1983, g6825, g6650, g7169, g7283, g1572, g8955, I6695, g4541;
wire g7059, g7920, g7578, g6008, I11835, g3691, I11014, g7459, g9221, I12205, I9463;
wire g7718, g7767, g4153, g4680, I7688, g6136, g4353, I11586, I12912, g6336, I14100;
wire I6223, g8038, g6768, I8913, g7582, g6594, g1961, g3879, g4802, g7261, I14683;
wire g3962, g5151, g7793, g3158, g3659, g6806, g5648, I6416, g3506, g7015, I12592;
wire g4558, g9068, I7126, I5926, I7400, I8859, I7326, I6115, I6251, g2921, g6065;
wire g6887, g6122, I10882, g6228, I5754, g3587, g6322, I11275, I9457, g8918, I16180;
wire g6230, g7246, g8967, I13746, I13493, I9393, g4511, I15660, g2895, g6033, g2837;
wire g7721, g5839, I9834, g4092, I13035, g3985, I12731, I11806, g4600, I7383, g4574;
wire g6096, g6496, g1679, I8097, g5172, g5278, g6845, g7502, I15550, g9198, g3545;
wire I8354, g738, g6195, g5618, g6137, g6891, g5143, g1831, g6337, g3591, g3832;
wire g4580, g9241, I7588, g3853, I14725, g7188, g5988, g2842, I9938, I10758, g1805;
wire g6807, g1916, g5693, g7216, g1749, g2298, I14082, g6859, g2392, I13193, g2485;
wire I11362, g7028, I13362, g3931, I8218, I15773, I6629, g4623, g7247, g1798, I6130;
wire g4076, g9319, I10940, g2941, I9606, g6342, g3905, I13475, g5621, I14848, g6255;
wire g6815, I10804, I6800, I9687, g3630, g6481, I14804, g7741, g4651, g5113, g6692;
wire g6097, I11437, I15839, g2520, I15930, g2640, g9211, g6354, g4285, I8727, g9186;
wire I5679, g4500, g9386, g6960, I15965, I7944, g1579, g1869, g7108, I10135, g7308;
wire I11347, g2958, I13347, g9026, I5831, g2376, g5494, g3750, I9570, I10406, I9341;
wire I10962, g1752, I14406, g3973, I9525, I11781, I12768, I15619, g9370, g1917, I9645;
wire I15557, g2829, g9125, g4024, I11236, g2286, g6783, g7758, g7066, I10500, I16168;
wire g7589, I6090, g2911, g4795, I8932, I5422, g7466, g4809, g6267, g6312, g3969;
wire I6166, I14049, g9280, I11821, I12881, g1786, g7365, g7048, I7347, g9083, g2270;
wire g4477, g7448, I13063, g7711, g4523, g6676, I11790, g6293, I13264, I6148, g7055;
wire g8219, g4643, g3666, I9158, I13137, I6348, g2225, g6129, g8640, g7455, g6329;
wire g6761, g2073, g5160, g7133, I7697, g9106, g7333, I13873, g9306, g6828, g1770;
wire g7774, g5521, g8958, g6830, g4634, g3648, g3875, g2324, g3530, I9111, g7196;
wire g4742, g9061, I15601, g9187, g4104, I10605, I11422, g6592, g3655, I15187, I14273;
wire I11209, I13422, I14106, I13209, g2540, I9615, g6221, I12003, g8765, g7538, I13834;
wire I6463, I10463, I16084, g2177, g7780, g9027, g5724, g2377, I14463, I12779, g5179;
wire g6703, g7509, g4926, I15937, g9200, I11021, I14234, g3884, g3839, g2287, g7018;
wire g4273, g7067, g8974, I7317, g5658, I15791, g7418, g6624, g7467, g6953, I6118;
wire I14795, g8225, g5835, g7290, g4613, g6068, g1888, I6872, g9145, g4044, g6468;
wire I12945, I9591, g4444, g1787, I6652, I11607, I6057, I12826, I12999, I11320, I15666;
wire I13320, I6457, g7493, g1675, g6677, g7256, I13274, I7775, g5611, g8324, g4572;
wire I7922, g2898, I15478, g2900, g6866, I12672, I7581, I13122, g9107, g4543, I10421;
wire I11464, g5799, I13565, I9794, I6834, g9307, g2510, g639, g2245, g6149, g3988;
wire I6686, g6349, g5674, g8177, g3693, I11034, g9223, I14163, g2291, I14012, I11641;
wire g6848, I15580, I13797, I12331, g5541, g3548, g1684, g1745, g6198, g1639, g2344;
wire g6855, g6398, I10541, I6121, g7263, g2207, g5153, g5680, I12897, I12448, I12961;
wire I9515, I9630, I14789, g2259, g9115, g4014, I7079, I12505, g9315, g1808, g4885;
wire I13635, g5744, g8199, g9047, g5802, g4660, g2923, I12717, g1707, I14325, I10829;
wire g8781, I10535, I5389, I5706, g8898, g4903, g7562, I15178, I10946, g8797, g6524;
wire I14828, g6644, g8510, I13164, I5371, g7723, I14121, g2215, I15953, g6319, g7101;
wire g2886, g3908, g7301, I7356, I13891, I15654, g4036, g6152, g6258, g6352, g6818;
wire g1575, g1865, I8483, g6867, g3567, I15417, g1715, g2314, I9440, I14291, I12433;
wire g4335, I9123, I15334, g7751, g2870, g5492, I12148, I13109, g4382, g1833, g5600;
wire I13537, g5574, I8790, g6211, g2825, g2650, g6186, g6386, I12646, g7585, g9017;
wire I9666, I15762, I12343, g4805, g6975, g4916, g4022, g3965, I5963, g1584, g6599;
wire g1896, g7441, I15423, g6026, I9528, g6426, I6860, g3264, I7053, I6341, I10506;
wire g5580, I9648, g9234, I10028, g9128, g6614, g6370, I14028, g3933, I8904, g9330;
wire g6325, g6821, g3521, g4560, I8446, g3050, g3641, I15909, I15543, g5736, g2943;
wire g6984, g7168, g6939, g3996, I11796, I12412, I8841, g5623, g7772, g6083, g7058;
wire I5957, g2887, g4873, g4632, g7531, g4095, g5076, g8870, I8763, g4037, g6483;
wire I12229, I9884, g2934, g5476, g7743, g4653, I6358, g4102, g6636, I15568, I15747;
wire I5865, g9213, g6106, g5175, g4579, I10649, I12011, g6306, I5715, g7505, g5871;
wire g3878, g8008, g4719, g6790, g7734, I6587, g3777, g7411, I9372, I10491, I15814;
wire g3835, I16116, g6387, I11522, g2096, I9618, I12582, g5285, g6461, g8768, I13663;
wire g3882, g2496, I7626, g4917, I15974, I6615, g6756, g8972, I10770, I12310, g1897;
wire g9090, g6622, g7474, I8757, g6027, g7992, g4265, g3611, g6427, g2137, g2891;
wire g5184, I15638, g9366, g2913, I12379, g5139, g5384, g6904, I12958, g9056, g8065;
wire I8315, I8811, g6446, g8228, g3981, g5024, g6514, I6239, g3674, g2807, I5362;
wire I11326, I9555, g5795, g5737, I15391, g6403, I13326, g5809, I5419, I9804, I10262;
wire I7683, g3997, I12742, g6345, g6841, I15510, I11040, I11948, I8874, g2266, g6763;
wire I7778, I16142, g6391, g1006, g4296, I6853, g3238, I9621, g5477, g9260, g5523;
wire I12681, I10719, g6637, g5643, I15014, g1801, g4553, g9063, g6307, I15586, I15007;
wire I8880, I14718, g3802, g7688, g6359, g6223, g2481, g8913, g1748, g2692, g4012;
wire g6858, g5742, g5551, g5099, g2497, I12690, g2354, I16165, g2960, g4706, I9567;
wire I7526, I5897, I14573, I10247, g3901, g7000, I13509, I15720, g9318, g9367, I11933;
wire g7126, I8935, I5425, g4029, g6251, g6315, g6811, g6642, g4371, I11851, g3511;
wire g5754, g9057, I16006, g7760, I14388, I7850, g9193, g3092, I14777, g3492, g4281;
wire g6874, g5613, I14251, g3574, g3864, g8342, I15340, g2267, g2312, g6654, g5444;
wire g5269, I7702, I15684, g8481, I12128, g1578, g1868, I9360, g2401, I7919, I10032;
wire g1718, g7779, g2293, g6880, g4684, I9050, I11452, g6595, g4639, I5682, I5766;
wire I11047, I13574, g2329, I6440, g7023, g9121, g4963, g2761, I5801, g9321, g8960;
wire g7423, g1582, I11912, I11311, I13912, I13311, g2828, I12298, I6323, I14061, g1793;
wire I7561, g7588, I10766, g2727, g4808, g6978, g6612, g7161, g1015, g5729, g3968;
wire g6243, g7361, I15193, I13051, I13072, g2746, I12737, g2221, g3076, g7127, g8783;
wire g7327, I12232, g1664, I6151, g1246, g2703, g8218, I8823, g5014, g206, g6328;
wire g6130, g7146, g6542, g6330, g7346, g7633, g1721, I11350, g3871, I7970, I13350;
wire I15475, g2932, g7103, I9271, g3651, g7303, I7925, g8676, g2624, g2953, I15222;
wire g6800, g3285, I13152, g8761, g4604, I10451, I10472, I13846, g3500, I14451, g7732;
wire I5407, I13731, I5920, I6839, I5868, I7320, g2677, g7753, g5178, g5679, I11413;
wire I5718, g7508, I13413, g6213, I5535, g2866, g4584, I12445, g4539, g8746, g8221;
wire g5335, g5831, g3838, g1689, g2149, g2349, I12499, g7043, g9141, g5182, I10776;
wire I12316, I9132, I6143, I9209, g7116, g1671, I7987, g5805, g5916, g5022, g2699;
wire g4019, g6090, g4362, I11929, I12989, g3077, g7034, g5749, g6490, g6823, g7434;
wire I14825, g3523, I14370, g6366, I12722, g7565, I7299, I5664, g3643, I12924, I13583;
wire g2241, g1564, g7147, I16122, I10151, I10172, g7347, I15516, I9558, g5798, I14151;
wire g1826, I12271, I14172, g6148, g6649, I14996, g6348, I8989, g8677, g7533, g3634;
wire I8193, g6155, I14844, g6851, g6355, I11787, I14394, I12753, g8866, g7210, g2644;
wire g3499, I8971, I12145, g1638, I11302, I7738, g5873, I13302, g5037, g9111, I12199;
wire g7013, g9311, g5437, I11827, g5653, g7413, I13743, g3926, g5302, I14420, I15208;
wire g2818, g6063, g4070, I12529, g2867, g3754, I9600, g8198, g8747, g4025, I14318;
wire g5719, I12696, g9374, I14227, I5689, I7959, g1758, g1589, I14025, I7517, I11803;
wire I7082, g2893, I15726, g7117, g6279, g5917, g7317, I14058, g6720, I5428, g6118;
wire g6167, g6318, g1571, g3983, g6367, g9180, g6872, g7601, I15607, g9380, g3862;
wire g5042, g1711, g2274, g6652, I12161, g4678, g3712, g8524, g6843, I15530, g5786;
wire g4006, g2170, g1827, g2614, g9020, g7775, g5164, g6393, g4635, g5364, I15565;
wire g2325, g2821, I12259, I10377, g1774, I12708, g7581, I11662, I10739, g4087, g4105;
wire g8152, I9076, g5054, g6834, g4801, g8867, I9889, I14739, g2939, g3961, g7060;
wire I11890, g1803, g7460, I15641, I6160, g5725, g4748, I11482, g6598, g3927, I5609;
wire I11248, g1780, I12244, I11710, I13710, g2636, g7739, g3014, I9651, g6321, g4226;
wire g8386, I5883, g2106, g8975, g3946, g2306, I13779, g9204, I15408, I15635, g6625;
wire g1662, g2790, g7937, I7762, I12810, g6232, I11778, g3903, g9100, I12068, I10427;
wire g7479, g9300, g5412, I10366, g6253, g6938, I14427, I5466, g6813, g7294, g4373;
wire g3513, I9139, g6909, g7190, g2622, I11945, I12337, I5365, I5861, I11356, I13356;
wire g1816, g5171, g4602, g7501, I11380, I10403, g5787, g4007, g2904, I14403, g7156;
wire g5956, g6552, g7356, g4920, g6606, g4578, I11090, I7928, I11998, g8544, g3831;
wire I11233, g2514, g4718, g8483, I8962, I7064, I11672, g1847, I9672, I15711, I13672;
wire I7899, g4535, g2403, g8636, g1685, g2145, g6687, g2345, g2841, I7785, g7704;
wire g4582, g3805, g3916, g9323, g6586, g8790, g2695, g4015, g2637, I11449, I12918;
wire g5684, g8061, g5745, I15492, g5639, I14127, g7163, g3947, I11897, g2307, I11961;
wire g7032, g2536, g5109, I13897, g8756, g3798, g5309, g7432, g6141, g6860, g2359;
wire g4664, I9499, g6341, I11404, g3560, g9351, g2223, I7844, I15982, g5808, g1562;
wire I6680, g6645, I16040, g4721, I14103, I11212, g2016, I7731, g5759, g8514, g3873;
wire g3632, g3095, g1817, g3495, g3653, I8180, I12322, g8145, g2522, I14181, g7157;
wire g2642, I8832, g6879, g7357, g6607, I12532, g3579, g3869, g6962, I8853, g6659;
wire I12158, g6358, g6506, g1751, I5847, I12561, I16183, g5604, I12295, g3917, g2654;
wire I10190, g1585, g4689, g6587, g9372, I15522, I15663, I14190, I9543, g6111, g8223;
wire g6311, g5833, I7814, I13646, g9235, g4028, g2880, I7350, I6574, g2595, I6864;
wire I11971, g4030, g8016, g8757, g5584, g1673, g6374, I14211, g9134, I15553, I13369;
wire g2272, I14088, g4564, I11368, g8642, I5562, I12364, I7769, g5162, g3770, g5268;
wire I9014, g5362, I10497, I15536, g1772, g6380, I9660, g6591, I15702, I13850, g6832;
wire I5817, g2982, g8874, g3532, I7967, g7778, g1743, g2234, g6853, g2128, g4638;
wire g2629, g6020, g2328, I10987, I12289, I5605, I10250, g7735, g4609, g6507, g4308;
wire g1011, I13228, g9113, g6794, g1856, I12571, g9313, I11011, I5751, g5086, g8880;
wire g3189, I13716, g5730, g7475, I16072, g3990, g2554, I14338, g5185, g4589, I10969;
wire g9094, g7627, g3888, I15062, g6905, g3029, g7292, g3787, g8017, g6628, I15933;
wire g7526, g5470, g5897, g3956, g5025, g6515, I11627, g6630, g4571, I12687, g3675;
wire I12976, g1573, g1863, g6300, I13112, g7603, I11050, I11958, g7039, I9422, I8351;
wire g8234, g4455, g2902, g7439, I12643, I5368, I11386, g1569, g453, I5772, g2490;
wire I6024, I5531, g2366, I12669, g7583, g7702, g4196, g5678, I6795, I10503, g3684;
wire g3639, g4803, g6973, g5006, g3338, g8800, g3963, g9360, I15574, g4538, g1688;
wire g2148, I15205, g2649, g4780, g1857, g2348, I7788, g9050, g5682, g5766, g5087;
wire g1976, g6969, I15912, I9095, g5801, g3808, g7276, g5487, I14315, I6643, I11793;
wire I11428, I12424, I13428, g3707, g6323, I14819, g4662, g2698, g4018, I12558, I14202;
wire I8172, I14257, I9579, g2964, I14055, I16020, g9379, I7392, g5755, I15592, I15756;
wire g7527, I14070, g3957, I12544, I6099, I9752, g4093, g8512, I8282, I16046, g1760;
wire g4493, g7764, g6351, g6648, g6875, g7546, g3865, I10384, g6655, g5445, g5173;
wire I11317, g3604, I13317, g5491, g3498, I14067, I14094, g4381, g8649, g6010, g3833;
wire I11129, g2872, g1924, g5169, g4685, g4197, I10801, g6410, g7224, I7520, g4021;
wire g5007, I13057, I14801, g2652, g1779, g2057, I7640, I12124, I12678, g6884, g2843;
wire g7120, g5059, g6839, g2457, g5578, g5868, g7320, g2989, g3539, g3896, I11245;
wire g5459, I14019, g2393, g5718, I12460, I12939, I11323, g1977, I11299, I13323, I14196;
wire I13299, I14695, g7277, g1588, I11533, g2834, g2971, I13533, g8063, g5582, I15405;
wire g6278, g8463, g2686, g6372, g7789, g5261, g3019, g9132, g5793, I12065, I8202;
wire g9332, g6618, g1665, g6143, g7516, I7765, g6343, g4562, g6235, g5015, g3052;
wire g9209, g9353, I7911, I10457, I8094, g7771, I14457, g6566, g4631, I13737, g372;
wire I15583, g7299, g4257, g6693, g6134, g8619, g7547, g6334, g4301, g5246, g2625;
wire g8872, g2232, g4605, g3086, g2253, g2938, g3728, I14001, I13261, I11880, g6555;
wire g6804, I7473, g2909, I6946, I10256, g6792, I11512, g1732, I9675, I13512, g3881;
wire I5383, I10280, g8971, g7738, g4585, I8264, g6621, g1944, g3897, g4041, I12915;
wire g9092, I8360, g6313, g7078, g7340, I7377, I10157, I13831, I6036, I14157, I12277;
wire I6178, g4673, g6202, g8670, I9684, g7035, I13499, I15803, I9639, g7517, I7287;
wire g6094, I14231, I9791, I6831, g5028, g4669, g1565, I8724, g5671, I11722, I12782;
wire I13722, I16090, I6805, g3635, I13924, I5633, g1681, g6776, I7781, I6422, g6593;
wire g4890, I12352, I13432, g2525, g3801, I14763, I13271, g2645, I8835, g5826, I12418;
wire I7797, g8606, I12170, g4011, I11461, g9076, g5741, g7110, I5732, g6264, g7310;
wire I11031, I13031, g5638, g6360, g2879, I13199, I11736, I11887, g9375, I7344, g2962;
wire g5609, I15003, I8799, g2659, g6050, I12167, g2506, g1820, I6437, I11696, g7236;
wire I6302, g3091, I13843, I16026, g7762, g3491, g4080, I14076, I14085, g4573, I11764;
wire g5758, I13764, g6724, I11365, g2275, g2311, I9539, g6179, I13365, g5466, g4713;
wire I10243, g6379, I11132, g7590, g9184, I13869, I5565, g2615, g6878, g5165, g4569;
wire g5571, g3920, I12022, g3578, g3868, g2174, g6289, g6777, I8802, g6658, g2374;
wire g5448, g1922, I9162, g7556, I13161, I10773, g5055, I12313, g6835, g2985, I9419;
wire I10268, g1581, g5827, I12748, g6882, I6042, I15651, I15672, g3582, g2284, I5914;
wire I13225, g7064, g2239, I7314, I10180, I16148, g1597, g9077, g2180, g5846, g2380;
wire I13258, I12900, I7870, I8901, g2832, I12466, g5396, I5413, g1784, g6799, I6054;
wire g2020, I10930, I15513, I11043, I6454, I12101, I6770, g6674, I13244, g7563, g8111;
wire g5780, g4000, I10694, g4126, I10965, g6997, g7295, g2794, I11069, g9104, I5936;
wire g9099, I6532, g9304, g2931, g3721, g6238, I6553, g5662, I13810, g8174, g6332;
wire I15717, I11955, g5418, g5467, I9025, g6353, g7194, I13879, I9425, g655, g2905;
wire I6012, g6744, g7731, g6802, g8284, g2628, g3502, g8545, I6189, g2630, g5493;
wire g8180, I14279, g4608, g4924, I5775, g7966, g2100, g3940, I10469, I11967, I11994;
wire g7471, I15723, g9044, g1942, I6029, g4023, I8736, I10286, I6371, g1704, g5181;
wire I12008, I9678, I15433, g5847, I6956, g6901, I14039, g4588, I11425, g5685, g5197;
wire I13425, g5397, I8889, g6511, g703, I11458, I15811, I10815, I12454, g2973, g1810;
wire g3430, g4665, I12712, g4051, g6092, I13918, I15971, I8871, I14187, g7150, I14677;
wire g7350, g6864, I7195, g2969, I13444, g6714, g7773, g4146, g7009, g4633, g2323;
wire I10937, I6963, g1568, I6109, I6791, g4103, I12567, I6309, g4303, I11086, I7807;
wire g3910, I12238, g7769, I10169, I7859, g4696, g1912, g5631, g7836, I14169, g5723;
wire g4732, g5101, I12382, I5356, g2528, I14410, g2351, g2648, I8838, I12176, I8024;
wire I12675, g6736, g8750, I10479, g6968, g2655, g8973, g1929, I12154, I5942, I9369;
wire g7229, g6623, g7993, I7255, g6076, I14015, I9407, g6889, I11656, I13656, g3589;
wire g8040, I11353, g9036, g4443, I13353, I11680, g8969, I8477, g9178, g9378, I13144;
wire g4116, g6375, g6871, g4316, I5954, g2884, g3861, g5041, g3048, g4034, I9582;
wire I8205, g6651, g9182, I5432, g4565, g8666, g9382, I15959, I15379, I8742, g2372;
wire g3774, I13631, I5568, g8875, g3846, g2618, g1683, I16129, g6384, g2235, g2343;
wire g6139, g5168, I12439, g5669, g4697, g6339, g4914, I14531, g2282, I7112, g1778;
wire g1894, g5058, g6838, g4596, I8754, g6024, I14178, g4013, g2134, g6795, g3780;
wire I10186, g6737, g2334, I15681, g6809, I8273, I12349, g5743, I6419, I10373, g1782;
wire I7676, g2548, I7293, I12906, I15429, I7129, I13023, g1661, I7329, I11224, g6672;
wire g2555, g6231, g3018, I11308, g2804, I12304, g9095, I13308, g5734, g1949, g6523;
wire I9502, g3994, I8983, g9102, g9208, I15765, g9302, I8862, g6205, I14334, g8172;
wire I15690, g2621, I8712, I7592, g5074, g3093, I6728, I8543, g5474, g1646, g7298;
wire g4601, I7746, g6634, g8667, I13816, g8235, g2313, g6742, g1603, g6104, I14964;
wire g6304, I15504, g2202, I12138, g4922, I10587, I13752, I11374, g3847, g2908, g5480;
wire I6425, g5713, g4581, I12415, g3700, g9042, g2494, I7953, g6754, g1583, g5569;
wire g4597, I9564, I5894, I11669, g7708, I13669, g9233, g7520, g8792, I11260, g6613;
wire g3950, g4784, I10569, g4739, I11392, g1952, I9910, g6269, g5688, I6006, I15533;
wire g2965, g6983, g1616, I14747, g7176, I5475, I7716, g6572, g6862, I11559, g4079;
wire I11525, I11488, I13559, g3562, I12484, I9609, g2264, g6712, g7405, g4668, I6087;
wire I6305, g3631, g7829, g2360, g2933, g3723, I12609, g7286, g7765, I7198, I10807;
wire g5000, I5646, g8094, I14807, g2641, I14974, I9217, I10639, g4501, g6729, g6961;
wire I13544, g3605, I13865, g2996, I9466, g5760, g9189, g7733, I12921, I13713, g9389;
wire g1970, I6226, g7270, I8805, I10265, I8916, g1925, g8776, g2724, g7225, g7610;
wire g9029, g6014, I14416, g2379, I13610, I12813, I16145, g6885, I6045, g4704, I13042;
wire g6660, g6946, I13255, g2878, I13189, I7644, g5183, I13679, g7124, I12973, g5608;
wire I9333, g2289, g6903, g2777, g9281, g5779, I10579, I9774, g4250, g2882, I11686;
wire I11939, I7867, g9297, I13460, g4032, I11383, g2271, I9396, I13383, g1789, g7206;
wire I6578, I6868, I5616, g6036, I13267, g6378, I6767, g5161, I16132, I10442, I15498;
wire g1987, g1771, I7211, g7287, I14442, g6135, I5404, g4568, I7386, g5665, g9109;
wire g5051, g6335, g6831, g9309, g3531, g5127, g2674, g6288, g6382, I16161, g8179;
wire I9018, g3743, I7599, I15924, I6015, I12400, g4357, g5146, g6805, g5633, I11218;
wire I12214, g7781, g2238, g2332, I10430, I13837, g3856, g2680, I14430, g2209, g2353;
wire I9493, g4929, g9201, I12328, I15753, g5696, g8882, g1945, g6947, g7510, g7245;
wire g6798, I12538, g1738, g3074, I16043, g5732, g7291, g3992, I14035, I15199, I10684;
wire I11455, g4626, I8233, I11470, g5240, g7344, I13617, g5072, g9098, I13915, g8799;
wire I12241, I14142, g1907, g5472, I9021, g6873, g7207, g6632, g6095, g3080, g8674;
wire g6037, g3573, I15696, g3863, I5789, g1959, g2901, g7259, g6653, I13277, g6102;
wire g6208, g6302, g8541, I13075, g2511, I7061, g6869, g1876, I12771, I11467, I11494;
wire I13595, g7488, I12235, g2092, g5434, I10193, I11037, I14130, I14193, g6752, g5147;
wire I13782, I11984, g8802, I11419, I6428, g9019, g9362, I13419, g3857, g7951, I8706;
wire g3976, I15225, I15708, I13822, I10475, I9301, g7114, I11266, g4661, g6786, I7145;
wire I6564, g4075, I5945, I8787, g4475, g5596, g1663, I6826, g6364, g7870, g5013;
wire g4627, I5709, g8511, g9086, g1824, I5478, g6296, I11194, g4646, I7107, g2623;
wire g6725, I9585, I10347, I10253, g5820, I7359, g9185, g4084, g4603, I5435, g7336;
wire I13524, I15657, g9385, g8864, I15068, g7768, g1590, g1877, I11401, g6553, g9070;
wire g7594, I8745, I10236, g2375, g2871, I12725, g3220, I15337, g2651, I6217, g6012;
wire g1556, I13118, g3779, g4583, I11864, I14175, g2285, I7115, g6189, I8808, g6389;
wire I7811, I16158, I9669, I13749, g7887, g7122, g4919, g3977, I6571, g6888, I6048;
wire I10516, g5581, I14264, g3588, I9531, g2184, I6711, g6371, g1785, g6787, g8968;
wire g2384, I11704, g5060, I13704, I11305, g9331, g6956, I13305, g5460, g5597, I11254;
wire g7433, g6675, g4616, I11809, I11900, g4561, g3051, I13900, I6333, I13466, I9505;
wire g1563, g2424, I12141, g2795, I8449, I12652, g9087, g9105, g5784, g4004, I15010;
wire I15918, g9305, g5739, I8865, g7496, g4527, g7550, g6297, g3999, g4647, g8175;
wire I8715, I7595, g8871, g3633, g2672, g2231, g7137, I14208, g8651, g2477, I16017;
wire g2643, g6684, I12135, g6639, g5668, g6338, I15598, I6509, g5294, g4503, g5840;
wire g6963, I7978, g6791, g2205, I12406, g6309, g5190, g4925, I5657, I12361, I7417;
wire g3732, I6018, g1557, g2634, g3753, I10614, g6808, I9573, g9045, I10436, g724;
wire I14614, g7266, g2551, I14436, g2104, g3944, I11693, g5156, g9373, g9091, g4120;
wire I16023, I7629, g6759, I10274, I14073, I6093, I8268, I13009, g1948, g8809, g7142;
wire g6201, g2926, g7342, I11008, g9369, I10565, g6957, g7255, g4617, I8452, g649;
wire g8672, g3316, g9059, I11476, I11485, I7800, g6449, g2273, g1814, g6865, I7554;
wire g7097, g7726, I13454, g7497, I10292, g2044, g7354, g5163, g6604, g5810, I13570;
wire I6021, g6498, g2269, g1773, I8486, I10409, g4547, g5053, g6833, I8730, g3533;
wire g5453, g2862, I15631, I12463, g4892, I11239, g2712, I14136, g9227, g1769, I9126;
wire I7902, g2543, g6896, I13238, I9760, g3013, g1918, g1967, g7112, g7267, I5966;
wire g5157, g2961, g4738, g8754, I5471, g6019, g6362, I13185, I6723, I13092, g7293;
wire g2927, I12514, I5948, g3936, I13518, g7129, I15571, I15308, g1822, g7329, g7761;
wire g4907, g2885, g4035, g2660, g2946, I12421, I14109, g7727, I15495, g4482, I7964;
wire g2903, g5626, g7592, I8766, I9588, g6486, I8105, I10283, g4656, g7746, g6730;
wire g9188, g7221, I15687, g9388, g3922, I15985, I14492, g9216, g6385, g6881, I12541;
wire I8748, g4915, I11215, g9028, g6070, I11729, g1895, g6897, g1837, I13577, g9030;
wire g6025, I6673, g6425, I14381, I13728, g5683, I12325, I9633, g2288, I7118, I7167;
wire I14091, g2382, g7068, I12829, I12535, I15669, g3784, I10796, g8014, I9103, I12358;
wire I13438, g3739, I6669, g4663, I6368, g2916, I15842, I8373, g5735, g1788, g3995;
wire g3937, g8903, g3079, g5782, g4002, I10390, I13906, I11284, I13284, g6131, g7576;
wire g6331, g5075, g3840, g2947, g7716, g7149, g2798, I11622, g1842, g7349, g6635;
wire I13622, g9108, g3390, g9308, I8868, g5627, g6682, g6766, g6087, I12173, g8178;
wire g6305, g6801, I6856, g4590, I10522, I15830, I8718, g3501, I9443, g5526, g7198;
wire g4657, g7747, g7855, g9217, g2873, g1854, g2632, I9116, I8261, g4556, g9066;
wire I13653, g5084, g5603, g1941, I6474, g2495, I8793, I9034, g2653, g7241, g6755;
wire g2208, g3942, I12760, g5439, g4928, I10862, g6226, g4930, g8916, g2869, I15610;
wire I15705, I10949, g9048, g4899, g4464, I9347, g1708, I9681, g7524, g6173, g2752;
wire g3954, g6373, I10702, I15678, g9133, g2917, g9333, g7119, g1812, g7319, I14904;
wire I8721, g1958, g2265, g6369, g7352, g7577, g6007, I12927, g9196, g7717, g6059;
wire g6868, g5616, g3568, g8873, I13484, g1829, g8632, I5842, I15065, g6767, g2364;
wire I12649, g2233, I10183, g1911, I10397, g7211, I5392, g3912, I14397, g4089, I12903;
wire g2454, I11200, g8869, g4489, g2770, g6793, I10509, g9018, g4557, g5764, g7599;
wire g9067, g1974, I10933, g7274, I15218, g6015, g4071, I6000, I7341, g2532, g8752;
wire g6227, g3929, I13921, I6326, I14851, g8917, g1796, g4242, g7125, g9093, I8428;
wire g6246, I7691, I15160, I13813, g8042, g5224, g7280, g8442, g6721, g8786, g5120;
wire I12262, g2389, g9181, g2706, g7544, I8826, g9381, I5812, g7483, I15915, I9460;
wire I9597, I6183, g4350, g2888, I6608, g9197, I6220, I10574, g2371, I8910, g2787;
wire g4438, g7106, I11732, g5617, g8770, g6502, I14205, g7306, g5789, g4009, g2956;
wire I16119, I14311, g7790, g5516, I15595, g6940, I5911, I8308, g7061, g7187, I7311;
wire g5987, g1849, g3778, I13692, I13761, g642, I8883, g7756, g6388, I10592, g5299;
wire I9840, g3735, g4918, g6216, g1781, I6051, I7374, I10780, g8012, I6127, I6451;
wire g6028, I14780, I12247, g6671, g7904, g1797, g2639, g7046, I11329, g3075, g2963;
wire g4229, I10350, I13329, g7446, g7514, g3949, g2309, g9101, I7545, I12388, g9301;
wire g4822, g7145, g8029, I7380, g7345, I12098, g8787, I16036, I7832, g5738, g6826;
wire g7763, g3526, g8956, g3998, g8675, g5709, I8333, g6741, I15589, g3084, g3603;
wire I5377, g785, g5478, I13241, I14413, g1694, g7107, g4921, g7307, g3850, I15836;
wire g2957, I8196, g7159, I7931, g1852, g1923, I6072, g6108, g7359, I9250, g5435;
wire g6308, g5517, g5690, I9363, g7223, g5482, g1701, g6883, I9053, g8684, g3583;
wire g4895, g8639, I6443, g7757, I7905, I11683, g4620, g8791, g4462, g2498, g6217;
wire g3919, g6758, g6589, g1886, I7204, I16009, I15616, I5781, g2833, g7522, g7115;
wire g7251, g8808, I6434, g3952, g7315, g7811, g7047, g9368, I8994, I10046, g6861;
wire g6365, g2584, I14046, g4788, g6048, I11515, I11991, g2539, g2896, g3561, g9058;
wire I13515, g8759, I13882, g6711, g1870, I11407, I13407, g1825, g6827, g3527, g8957;
wire g6133, g6333, I14282, g3647, I9929, g2162, I7973, g2268, g6774, g2362, I12629;
wire g3764, g4085, I12451, g6846, I12472, I12220, g8865, g3546, g5002, I14743, I8847;
wire g2052, g5402, g5824, g7595, g6803, g2452, g8604, g3503, g3970, g1768, g9074;
wire g6538, I13441, I5852, I5923, I11206, I7323, g6780, g6509, g1806, g1943, I6820;
wire g7243, I6936, I11725, I12776, I13725, g2728, g2486, g6662, g6018, I6317, g1887;
wire I16176, I13758, I15693, I12355, I13435, g1934, g2185, g6290, g4640, g2881, I7648;
wire I16154, I7875, I12370, g4031, g7130, I7655, g3617, g6093, I11744, g7542, g2470;
wire g7330, g2897, g6493, g6256, I12151, g6816, g5785, I12996, g4005, I13940, I8101;
wire I8817, I14662, g3987, g3771, I11848, I9782, I11398, I12367, I12394, I6060, g6381;
wire g4286, I11652, g6847, I6460, I6597, I10482, g3547, g6700, g6397, I10552, I8751;
wire g3892, I11263, I10204, I9627, g2131, I6784, g2006, g2331, I12319, g4733, I11332;
wire g5844, I13332, g6263, g4270, I5972, g2635, g1807, g6950, g8881, g9126, g4610;
wire g2105, I7667, g3945, I12059, I10786, I12025, g2487, I9084, g5731, I9603, I13962;
wire I14786, g7512, I9484, g3991, g7090, I6294, I9850, g594, I10356, I15382, I11500;
wire g6562, g7366, g4069, I15519, g5071, g3078, g3340, I10826, I15675, I10380, g5705;
wire g5471, g7056, g6631, g4540, g2226, I7548, I10998, I12044, g6723, g7456, I13048;
wire g7529, g6257, g3959, g1815, g6101, g7148, g6817, g9183, g6301, g7348, g3517;
wire I11004, g3082, g9383, I8772, I7804, g9220, I11221, g7155, g7355, g6605, I7792;
wire I12301, g8678, g1726, g3876, g8131, I12120, g2373, g2091, g8406, I13613, g1960;
wire g5814, g7260, g6751, g5150, I8011, I9561, g8682, g8766, g5038, I5395, I8856;
wire g2283, g7063, I12699, g9161, I16138, I13106, g9361, g2007, I13605, I10448, g7463;
wire g5009, g2407, I6163, I14448, g2920, g2868, I6363, I15501, g9051, I15729, g2459;
wire I15577, g4898, g6441, I13463, g9127, g2767, g4900, g1783, I7908, g5769, I11951;
wire I11371, g8755, g636, g7279, g8226, g5836, g4510, I13234, g4245, I12427, g7720;
wire g7118, g5918, g2793, g7367, I12632, g9103, g9303, g1676, g2015, I8480, g6368;
wire g7057, g8173, g4344, g6772, I6157, I12403, I12547, g1828, g2664, g2246, g4259;
wire g5822, g6890, g7549, g1830, g4694, I15622, g1727, g3590, g3877, I10433, I5692;
wire g8602, I10387, I12226, I14433, g7686, g8407, g4088, I12481, g9072, g3657, g4923;
wire g2721, g6505, g8868, I14148, g6011, I5960, g1746, I14097, g6856, g4701, I10646;
wire g8767, g9043, g3556, I13012, I10343, I14646, g3928, I16052, g8582, g9116, g6074;
wire g3930, g2502, g9316, I11473, I13541, g4886, I10369, g9034, I12490, g8015, g2940;
wire g8227, g4114, g7253, I11359, I12376, I12385, I13359, I9892, g5462, g2689, g6573;
wire g6863, I11920, I12980, I7878, g8664, I8760, I11434, g3563, I10412, g2216, g6713;
wire g1677, g7519, g7740, g4650, I7658, I5401, I12888, I13828, I5676, I14133, g2671;
wire g9210, g1576, g6569, g1866, I7882, g5788, g4008, I10896, I6894, I11344, g3844;
wire I13344, I15484, g1848, I10716, I13682, g4594, g5842, g2826, g1747, g1855, I6075;
wire g6857, g7586, I9907, I13173, g5192, I10582, g3557, g5085, g4806, I7981, I6949;
wire I12190, g3966, I8977, g2910, g3071, g3705, g9117, I12520, g2638, g4065, g9317;
wire I8161, g8689, g4122, I15921, g4465, g7141, I14925, g3948, g4934, g7341, g8216;
wire I6646, g2308, I7132, I13134, I7332, I8665, I12211, I14112, g6326, g7525, g7710;
wire g3955, I7680, I11506, I14378, g2883, I6084, I7353, g8671, I11028, I13506, I12088;
wire I6039, g4033, I13028, g6760, I14603, g5520, I15184, g4096, g8564, g3038, g1818;
wire g1577, g1867, g9060, I9310, I7558, I10681, g5812, g6183, g7158, g2365, I12659;
wire g6383, g7358, g5176, g4195, I9663, g6220, g7506, I15732, g4891, I13927, g4913;
wire I12250, g658, g8910, I16100, g6779, I14857, g3769, I6952, g8638, g3836, g5829;
wire g7587, I13649, g5286, g1975, I5747, g4807, g6977, g7111, I5855, I5398, g3918;
wire g2774, g7275, g7311, g3967, I6561, I11648, I10690, g6588, I11491, I11903, g9079;
wire I13903, g8883, g6161, I7492, g6361, g4266, g2396, I7864, I10548, I13755, g5733;
wire g7174, g6051, g3993, g8217, I13770, I11981, I9657, I12968, g1821, I15329, g6327;
wire g2780, I6764, g3822, g5610, g2509, I15539, g5073, g5796, I8565, g5473, g7284;
wire g6146, g4081, g7239, g6346, g7545, I6970, g2662, g5124, g7180, g6103, g4692;
wire g7591, g6303, g2467, I9064, I13767, I13794, I11395, g5469, g2290, I7262, I10128;
wire g6696, g3921, I9785, I5577, g4960, g7420, I11633, g5177, I12894, g7507, g8774;
wire g5206, I7623, g2256, I11191, g2816, I13719, g6508, g6944, g3837, g6072, I11718;
wire g3062, I14298, g9032, I5386, g3462, g1756, g2381, I5975, I11832, g8780, g9053;
wire I12202, g4112, g7905, g4267, g2700, I7651, I16107, I8820, I11440, g2397, I12496;
wire g5199, g1904, I12111, g6316, g7515, I11861, g8662, g5781, g4001, g6034, g8018;
wire I13861, I9089, g8067, g2263, g7100, I13247, I6299, g7300, I11389, I11926, I12986;
wire g5797, I15414, I13045, g6147, I5984, g9157, g6347, I5939, I13099, g3842, I13388;
wire g8093, g6681, I11701, g8493, I13701, I10512, g3085, I8775, I7838, I8922, I11251;
wire I11272, g7750, g3485, g2562, g1695, g6697, g1637, g5144, g4592, g5344, g6210;
wire I5636, g2631, g4746, I12877, g8181, g6596, g5207, g8381, g3854, g2817, g3941;
wire I7672, I16135, g4703, g5819, g8685, g7440, I10445, I7523, I14445, I12196, I6078;
wire g2605, I13140, I9350, g7123, g8421, g5088, I8784, I13997, I8739, g1757, g5488;
wire g4932, I12526, I15759, g5701, g6820, g4624, I9009, I6959, g3520, g6936, g3219;
wire I6517, g3640, I16049, g6117, g1811, g6317, I7551, I7104, g3812, I12457, g7528;
wire I14722, g7151, g3958, g7351, g4677, g6601, g7530, I12866, I8190, g8562, I9918;
wire I10271, g5114, g4576, I15940, I13447, g8631, g2673, g6775, g3829, g6922, I5763;
wire g3911, I6214, g6581, g5825, I14342, g8605, I14145, I12256, I14031, g4198, I7044;
wire g6597, g9075, I13451, I13472, I14199, I12280, g3974, I6663, I13628, g8751, g2458;
wire I5359, g6784, g2743, g3610, g2890, g5768, I10528, I16033, g8585, g1612, I10393;
wire g7172, g1017, I7712, I14330, g2505, g8041, I15962, g2011, g3124, g5806, I5416;
wire g1935, g3980, g6937, g7143, I11591, g2734, g7343, I13776, g9039, g4524, g6294;
wire g6840, g4644, I6590, I13147, g8673, g3540, I15833, g4119, I9837, g6190, g2074;
wire I6657, g6390, g7134, I12885, g7334, I13825, g2992, g4258, I11858, g4577, g6501;
wire g7548, g8669, g4867, I13858, I14709, I10259, g6156, I12511, g6356, g5433, I10708;
wire g7555, g1800, I12763, g3287, g8772, I7885, I5654, I8357, I6930, g2573, g2863;
wire g7792, g2480, I15613, I9788, g8743, g3849, g6704, I15947, g5845, g4599, g5137;
wire g5395, g8856, g7113, g3898, g8734, g4026, g7313, g4274, g4426, I7036, g6250;
wire g6810, g4614, g6363, g4370, I5978, g3510, I10810, g6032, I11446, g4125, I14810;
wire I11227, g6432, g5807, I14657, g7094, I12307, I11025, I12085, g2976, I7335, g1823;
wire g7494, g7518, g5266, g6568, g4544, I11203, I5542, I13203, g7776, g1649, I7749;
wire g7593, g3819, g4636, g3694, g2326, I14792, I9520, g6357, g4106, I15507, I12942;
wire g3852, I6471, g3923, g4306, I8778, I11281, I12268, g9320, g5481, g3488, I7947;
wire I13281, g1698, I6242, I16173, I12655, I11377, g7264, g5726, g5154, I10919, I9005;
wire g7160, g7360, I11562, I11645, I13562, g7521, g4622, g4027, g2183, g3951, g7050;
wire I6254, g2383, g2924, I12839, I12930, I8949, I7632, I7095, I12993, I10545, g6626;
wire I11290, I13290, I7495, I14079, g4904, g4200, I13698, I7302, I12965, I12131, g9299;
wire I6009, g3870, I8998, I5512, g4003, I9974, g5112, g3825, g3650, g5267, I12487;
wire g4841, g2161, I8084, g1652, g2361, I7752, I12502, g4191, g1843, g8760, g3008;
wire I8850, g2665, g7289, g7777, g6683, g5401, I10125, g4695, I10532, g4637, I5649;
wire g7835, g2327, g5129, g6778, g5761, g3768, I10783, g6894, I13403, I13547, g4307;
wire g4536, g2999, I14783, g3972, g1686, g5828, g2346, g2633, I12469, g9244, I10561;
wire I6229, g8608, g8220, I10353, I12286, g6782, I7164, I10295, I8919, g3943, g9140;
wire I9177, g9078, g9340, I13481, g5592, I14680, g6661, g6075, g4016, I8952, g699;
wire I12038, g5746, g6475, g9035, g1670, g3465, g8977, I7296, g3934, g9082, g3230;
wire g4522, g4115, g4251, g6292, I12187, g4811, g4642, g7541, g2944, g2240, g1938;
wire g1813, g6646, g7132, I8986, g8665, g7332, I13490, g1909, g7353, g6603, g3096;
wire I5872, I13956, g5468, g6850, g3496, g7744, g4654, I13103, g3845, g2316, g9214;
wire I5989, I7389, I11824, g5677, I7706, I13888, g3891, I8925, g3913, I10289, g9110;
wire g9310, g6702, g7558, I7888, g4595, g4537, I15927, I7029, g1687, I7371, g2347;
wire I12666, g5149, I14288, I14224, I9344, I12217, I7956, g1586, I6788, I12478, g2533;
wire g8753, g3859, g4612, g7511, g4017, I15648, g2914, I8277, g5198, I9819, g8072;
wire g9236, g2210, g6616, g4935, g7092, I5670, I15604, g7492, I14816, g1570, g1860;
wire g8443, I6192, g7574, g6004, I15770, I10687, g4629, I10976, g6404, I12223, g4328;
wire I14687, g7714, g6647, g4130, g4542, I10752, g3815, I7338, g6764, I14374, I10643;
wire g3692, I13088, g9222, I14643, g2936, g3497, g5524, g7580, g4800, g5644, I15845;
wire g3960, I8892, g1879, g4554, I11497, g9064, I15990, I5552, g7262, g5152, g5258;
wire I14260, g7736, g5818, I10842, g6224, g5577, I14668, I11659, g5717, I13126, I13659;
wire I8945, I11987, g6320, I12373, I6431, I13250, I14489, g2922, g1587, g3783, g8013;
wire I10525, I10488, I16061, I10424, g7476, I8709, g3979, I14424, I6376, g5186, I10558;
wire I8140, I12936, g9237, I9136, I11296, I9336, g6617, g6789, I13296, g4512, g2460;
wire I7098, I8907, I11338, g7722, I12334, I13338, I9594, I7498, g5026, I6286, g3676;
wire g9194, g5426, I6911, I8517, g7285, g2784, g5170, g3761, g4056, g7500, I11060;
wire g9089, I13060, g6299, g5821, I11197, g3828, g4649, I7584, I11855, I6733, g3830;
wire I6974, I15388, I15324, I6270, g2937, I11870, g7139, g9071, g5939, I10705, g6892;
wire g1832, g2479, g7339, I13527, g2668, I14042, g1853, g2840, g4698, g8775, g3746;
wire g5083, g7838, I5879, g7024, g7424, I7362, I12909, I14270, g7737, I10678, I6124;
wire g8581, I14124, g6945, I12117, g1794, I11503, g2501, I11867, I11894, I10460, I13894;
wire g4463, I14460, g6244, g7077, I9496, g7231, g3932, g5790, g7523, I9845, g6140;
wire g3953, g6340, I11714, g9350, g5187, g5061, I14267, I14294, g6478, g8784, g2942;
wire g5461, g4279, I11707, g7205, I13707, I13819, g5756, g6035, g6959, I7728, I11257;
wire g5622, g4619, g5027, g6517, I11818, g3677, g5427, I15871, I11055, I13979, I5374;
wire I13496, g7742, g4652, g7551, g7104, g6876, g7099, g4057, g7304, g8668, I11978;
wire I6849, g3866, g2954, g4457, g7499, I8877, g2810, g2363, g6656, g9212, I12639;
wire I16151, g3716, g5514, I5545, g5403, g5145, g2453, I5380, g5841, g3848, g1750;
wire I6900, I12265, g7754, I10160, g5763, I9142, g5191, g8156, g3855, I14160, g3398;
wire I8928, g7273, I6245, I9081, I12391, g4598, g6110, g6310, I6291, g7044, I10617;
wire I15628, g4121, I5559, g2157, g7269, g6663, g4670, g5159, g4625, g7983, I10277;
wire I11018, I13196, I7635, I13695, g6824, g7712, g1666, g3524, g4253, g2929, g4938;
wire g6236, g4813, I12586, g7543, g5016, g5757, g8810, g3644, I7305, g8363, I15776;
wire I16058, I10494, g4909, I12442, I5515, I14623, I8844, g5522, g5115, g6877, g5811;
wire g5642, g2626, g3577, g7534, g7729, g3867, I15950, I13457, g1655, g6657, I7755;
wire g4552, g9062, I11917, g4606, g6556, I10418, g6222, I12041, g5874, I9001, I14822;
wire g7014, g4687, I8966, I12430, I11001, g5654, I12493, g7414, I9129, I15394, g3975;
wire g6064, g4586, g6899, g2683, g6785, I11689, I11923, I12340, I12983, g7513, I5969;
wire I12806, I12684, I7602, g2894, I15420, g4570, g4341, g9298, g9085, I8814, g1667;
wire g4525, g4710, g7178, g2782, g6295, g1235, g5612, I12517, g6237, g4645, I13157;
wire g2661, g5417, g1566, g7135, g6844, g7335, I11066, I13066, I13231, g7288, g6194;
wire I5528, g2627, I14118, g5128, I9624, g2292, I14022, g6089, I12193, g6731, g4607;
wire I8769, I13876, I13885, g5542, g7022, g2646, g7422, g4659, g7749, g1555, I12523;
wire g4358, g1804, I6887, g8683, I13854, g6071, g9219, g1792, g2039, g3061, g3187;
wire g6471, g8778, I14276, I14285, g2484, g9031, g5800, I5410, g3461, g6242, I14305;
wire g9252, g4587, I12475, I6033, I9576, I10466, g6948, g4111, I5839, g7560, g4275;
wire g4311, g9376, I15738, I15562, I15645, g6955, g4615, g3904, g8661, I10177, I15699;
wire I6096, g6254, g6814, g7095, g3514, g2919, g7037, g6150, g7495, g1908, g7437;
wire g6350, g7102, g7208, I6195, g7302, I13550, g6038, I5667, I11314, I6337, g3841;
wire I13314, I11287, g2276, I12253, g6773, I13287, g1567, I16103, g7579, I14064, g6009;
wire g3191, g4545, g2616, g7719, g2561, g5490, g691, g5823, g534, g5166, I11596;
wire g4591, g8603, I13054, g8039, g1776, g6769, g7752, I11431, g9073, g6836, g4020;
wire g6212, g2404, I5548, I8895, g2647, g5529, g3159, I10166, g5148, g3359, g5649;
wire g6918, g6967, I5555, I11269, I14166, I14009, g2764, g7265, g9324, g7042, g2546;
wire I11773, g5155, g4559, g9069, I11942, I11341, I13773, g3858, g7442, g8583, I13341;
wire g4931, I6248, I7564, I9258, g3757, g2970, g6229, I15481, I10485, g6993, g1933;
wire g7164, g7364, I6081, g2925, g9177, g7233, g9206, I10555, I10454, g6822, g3522;
wire I14454, g7054, g2224, g3642, I13734, g3047, I10914, I11335, g7454, g4628, I14712;
wire I13335, g7770, g5463, I6154, g7296, I6354, g4630, I13930, g7725, I11838, I5908;
wire g4300, g7532, g1724, I7308, g3874, I12208, I13131, g3654, g9199, I15784, g8647;
wire I15956, g2617, g2906, I15385, g1878, g5167, I14238, g5367, g5872, I13487, g7412;
wire g6462, g8925, g4969, g7429, g9144, g9344, g4123, g8320, I8431, g9259, g8277;
wire I8005, g4351, g8299, g6941, g4410, g8892, I7994, g5552, g8945, g8738, g6431;
wire g4172, g7449, g8709, g6176, g6005, g4343, g8078, g8340, g6405, g4282, g7604;
wire g1714, g5570, g8690, g7833, g4334, g8876, g6733, g6974, g4804, g8915, g7419;
wire g8310, g4494, g8824, g8877, g6399, I9330, g9142, g8928, g5020, g4933, g8930;
wire I8114, g8064, g7678, g4724, g7087, g4379, g8295, g8237, g6923, g4878, g8844;
wire I8594, I9166, g8089, g8731, g4271, g6951, g8071, g8705, g4799, I8033, g8948;
wire g5969, g7602, g7007, g5123, g4132, I8496, g4238, g8814, g6408, g8150, g4744;
wire g8438, g6972, g7415, g8836, g4901, g6433, g8229, g9349, g8822, g6395, g8921;
wire g7689, g5334, g5548, g4968, g6266, g8837, g7030, g8062, g8620, g8462, g9119;
wire I8001, g7564, g9258, I8401, g4175, g4375, g5313, g6726, g6154, g8842, g7609;
wire g8298, g5094, g9274, g4139, g4384, g4838, g8854, g7217, g8941, g4424, g6979;
wire g5593, g6112, g4077, g6001, g6401, g8708, g7827, g5050, g1725, g6727, g8405;
wire g4099, g4304, g8829, g8286, g8911, g8733, g8270, g8610, g9345, g4269, I8524;
wire g2781, g8069, g4712, g7181, g9159, g9359, g8377, g7197, g7700, g7021, g4729;
wire g4961, g9016, g8287, I8186, g5132, g8849, I7995, g9251, g4414, g3313, g7631;
wire g8291, g3094, g4436, g6577, g7605, g4378, g4135, g5092, g4182, g4288, g9272;
wire g8259, g5714, g8088, g8852, g8923, I8461, g7041, g4422, g8701, g2768, g9328;
wire g4798, g9130, g6125, g2972, I8046, g8951, g8314, g4437, g8825, g8650, g4302;
wire g1728, g8336, g6061, g8943, g6046, I8115, I8642, g8322, g6003, g8934, g9348;
wire g7713, g6145, g4054, g4454, g5077, g4532, g6107, g8845, I9202, g8337, g4412;
wire g5104, g6757, g9279, g4389, I8612, g6416, I8417, g9118, g4787, g6047, g8266;
wire g6447, g4956, g2979, g5044, g8081, g8815, g7183, g7608, g8692, g8726, g4138;
wire g4109, g4791, g4707, g6417, I8090, I8490, g4201, g8267, g8312, g6629, g4957;
wire g4049, I8456, I8529, g8293, g8329, g7696, g5513, g4098, g6554, g8828, g8830;
wire g8727, g5436, g7240, I8063, g8703, g4268, g8932, g6166, g8624, g8953, g4052;
wire g8068, g4452, g6056, g6456, I8057, g7681, g9158, g5560, g4086, g4728, g4486;
wire g8716, g7596, g4504, g4185, g9275, g4385, g8848, g5579, g4425, g2386, g5442;
wire g6057, g4131, g8319, I8552, g8258, g6971, g8717, g7597, g7079, g8274, g4445;
wire g4091, g4491, g8325, g8821, g4169, g5029, g4369, g8280, g8939, g4407, g4059;
wire g4868, g8306, g4793, g8461, g8622, g4246, g8403, g8841, g5049, I8020, g8695;
wire g8307, g9278, g4388, g8359, g4216, g9143, g9343, g7626, g8858, g4430, I9534;
wire g9334, g8315, g4826, g6239, g5019, g2935, g7683, g5452, g8654, g6420, g4108;
wire g4883, I8040, g4066, g8272, g4466, g8978, g8612, g3429, g6204, g4365, g4048;
wire g8935, g5425, g4448, g4711, I8528, g8328, g4133, g4333, g8542, g8330, g4396;
wire g9160, g6040, g5105, g7616, g7561, g4067, I8618, I8143, g3049, g8090, g6151;
wire g8823, g5045, g5091, g4181, g8456, g9271, g4397, g8851, g4421, g8698, g8260;
wire g5767, g6172, g9238, g8720, g4101, g8318, g8652, g8843, I8593, g8457, I10597;
wire g1753, g8686, g7709, g8321, g6908, g4168, g6567, g4368, g8938, g5428, g8813;
wire g5030, g4058, g4743, g8740, g6965, g4411, g8687, g6160, g3226, g4074, g5108;
wire g6641, g7002, g6996, g5066, g8860, g8341, g8710, g9384, g8645, I8209, g7657;
wire g8691, g5048, g9024, g8879, g8607, g8962, g6611, g1739, g8275, g8311, g4400;
wire g6541, I8574, g5018, g5067, g5093, g9273, g7557, g4383, g4220, g8380, g8832;
wire g7071, g4779, g7705, g8853, g7242, g4423, g3188, g5700, g4361, g8931, g4127;
wire g4451, g4327, g6574, g7038, g8628, g8300, g9014, g7212, g5817, g4472, g3466;
wire g8440, I8523, g5585, I8643, I9535, g6175, g8323, g9335, g5441, g4434, I9261;
wire g4147, I8551, g9022, g4681, g8151, g8648, g7837, g5458, g3509, I8613, g8839;
wire g9037, g6643, g4936, g4117, g4317, g8278, g7192, g8282, g5080, g5573, g8693;
wire g8334, I8014, g1919, g6044, g7031, g6444, g7252, g8621, g4937, g8313, g4840;
wire I8436, g4190, g4390, g5126, g9012, I8288, g4356, g9371, g6414, g8264, g4163;
wire g8933, g7177, g4053, g5588, g4453, I8495, I8437, g6182, g8724, g8379, g7199;
wire g6916, g6022, g8878, g6422, g8289, g8835, g8271, g8611, g5043, I8296, g6437;
wire g5443, g7694, g5116, g8238, g5034, g8332, g7701, g8153, g4778, g8744, g7215;
wire I8412, g4782, g6042, I8029, g8901, g6054, g4526, g7008, g2889, g7136, g5117;
wire g8714, g9025, I8109, g4702, g6412, g7228, g6990, g8262, g6171, g8736, g4276;
wire g6429, g7033, g9131, g8623, g8076, g7096, g8722, g7195, g1844, g5937, g5079;
wire g4546, g5479, g6745, g8285, g9226, g6109, g4224, g8384, g8339, g4320, g8838;
wire I8019, g8737, I8052, g4906, g4789, g6049, g8077, g7692, g8643, g6715, g6098;
wire g5032, g5432, g4299, g9015, g8742, g8304, g8926, g6162, g6268, g7001, g8273;
wire g6419, g7676, g6052, g4078, g8269, g4959, I8006, g4435, g4517, g4690, g4082;
wire g8712, g8543, g7703, g8729, g8961, g9247, g8927, I8045, g5894, g8660, g8946;
wire g7677, I8491, g6006, g4236, g8513, g6406, g5475, g3190, g6105, g4877, g8378;
wire g6487, g7699, g8335, g8831, g8288, g8382, g5484, I8015, g8749, g4785, g6045;
wire g5583, g6091, g8947, g6407, g6578, g4194, g8653, g4394, g8302, g7186, g6582;
wire g1733, g8719, g4705, g6415, g7614, g5970, I8028, g8265, g4955, g4254, g4814;
wire g4150, g4038, g9021, g8296, g4409, g8725, I8108, g6689, g7027, g5547, g7427;
wire g1898, I8589, g6428, g6430, g7003, I8455, g7695, g8281, g5078, g6638, g7536;
wire g8297, g5082, g8745, g4837, g8338, g8963, g4062, g7416, g8309, I8418, g6448;
wire g6055, g7654, g4192, g4392, g6196, g6396, g8715, g7537, g8833, g7017, g7417;
wire g8584, g9080, g6418, g6994, g7128, g8268, g5064, g8362, g4958, g4176, g4376;
wire g7554, g5563, g1913, g6021, g6421, g8728, g8730, g4225, g8385, I8041, g4073;
wire g4796, g8070, g5089, g4473, g5489, g4124, g4469, g4377, I8058, g8331, g9023;
wire g4287, g7698, g8087, g8305, g4199, g5438, g4781, g6041, g8748, g9327, g4797;
wire g9146, g9346, g3002, I8573, g6168, g7652, g6058, g7193, I8569, g6743, g4819;
wire g8283, g9240, g8059, g8920, g8459, g6411, g8718, g7598, g3222, g8261, g6474;
wire g7625, g8793, g6992, g7232, I8000, g4314, I8400, g9147, g5062, g9347, g4825;
wire g8721, g7552, g7606, g4408, g9013, g5298, g6976, g8940, I8588, g4230, g6400;
wire I8127, g4433, g7691, g5031, g7607, g8826, g4395, g8741, g5005, g2827, g6423;
wire g5765, I8240, I8072, g8609, g8308, g7615, g3229, g8066, I8034, g4142, g4342;
wire I9222, g6999, g4255, g6633, g8711, g5069, g4097, g7832, g4497, g8455, g4154;
wire g8827, g8333, g6732, g8846, g6753, g7559, I8413, g5287, g4783, g6043, g4312;
wire g7628, g6434, g8290, g4129, g8256, g4830, g8816, g6914, I8460, g6013, g6413;
wire g8700, g7323, g8263, g8950, g4068, I8079, g5314, g8723, g8257, g8817, g8301;
wire g7010, g6060, g4699, g6460, g4398, g5008, g7278, g6995, g8441, g7235, I8432;
wire g9084, I8053, g7282, g5065, g5122, g4319, g7693, I8568, g4352, g5033, I8157;
wire g8458, g5096, g4186, g9276, g4386, g6954, g8074, g6053, g4083, g8080, g4483;
wire g3259, g8713, g5142, g6157, g5081, g9120, g4187, g9277, g4387, g8688, g8857;
wire g8976, g4427, g4514, g5783, g7724, g7179, g4403, g8326, g4145, g4391, g5001;
wire g7658, g4107, g1834, g7271, g4159, g8383, g8924, g7611, g8779, g6949, g4315;
wire g4047, g8361, g6998, g7238, g5624, g7680, g8327, g6039, g5068, g6439, I8546;
wire g8303, g8696, g8732, g4272, g8944, g5699, g4417, I8617, g7600, g4128, g3081;
wire g8316, I8299, I8547, g6970, g8147, g5119, g8697, g8914, g4902, I8078, g7175;
wire g5599, g4490, g4823, g4166, g8820, g4366, g8936, g6771, g8317, g4529, g5125;
wire g7184, g4155, g5984, g4355, g8922, g6738, g8060, g5106, g6991, g8460, g9038;
wire g8739, g4720, g4118, g4167, g4367, g4872, g7634, g8937, g8079, g8294, g5046;
wire g8840, g4193, g4393, g4549, g6915, I8064, g8942, g2912, g5107, g8704, g6002;
wire g6402, g8954, I8237, g6762, g4740, g3258, g5047, I8089, g8912, I8071, g6464;
wire g8929, g3614, g7036, g7679, g8626, g3984, g5017, g4691, g2949, g7182, g6394;
wire g4962, g4158, g6966, g8735, g8075, g8949, g7632, g7653, g8292, g2952, g6438;
wire g4284, g4239, g5090, g8646, g6409, g4180, g9270, g4380, g4832, g8439, g2986;
wire g4420, g4507, g4794, g8702, g8919, g8952, g8276, g5063, g4100, g7553, g8404;
wire g5118, g8764, g5057, I14941, g5193, g9291, g5549, g7029, g7787, g6249, g8906;
wire g5232, g8987, g5253, g7791, I8225, I15250, g8991, I9107, g9008, g2214, g7575;
wire g9136, g8907, g8082, g5710, I9047, g9122, g6270, g6610, g6124, g6980, I14484;
wire g9137, g9337, g7086, I15055, I15111, g5545, g7025, g4264, g8899, g8785, I15019;
wire g6144, g9154, g9354, I15018, g4179, g7682, g6694, g5204, g9267, g9001, g8966;
wire g7445, g5040, g5440, I15102, g2229, I14771, I15231, g8773, g8009, g8769, g7227;
wire g6934, g8993, g6913, g5235, g5343, I15085, g5566, I14759, I15054, I15243, I14758;
wire g4736, g8895, g7428, g9352, g7826, g8788, g5202, g5518, g4737, g7165, g5264;
wire g8176, g9387, g2206, I14951, g9046, g6932, I15169, g9003, g8796, g8980, g6716;
wire g7421, g6699, g5238, g4927, g5209, I15084, I15110, g8900, g5511, g6717, g3160;
wire g8886, g2230, I15242, g5722, g2845, I15230, I15265, g4786, I13553, g8887, g7080;
wire g4364, g9148, I14767, g9355, g3541, I14990, g5231, g5205, g8891, I15041, g6115;
wire I15275, g4297, g7220, g5572, g8154, I14766, g6935, I15165, g8979, g5036, g3339;
wire I15253, g7443, I14754, I15175, I15264, g9358, g7697, g6698, g6964, g5208, g9174;
wire I15021, g9239, g5265, I15073, I15274, g6457, g5233, g6686, I15292, g8893, g7784;
wire g6121, I14366, g5706, g6740, g4283, g8984, I15109, g9123, I15283, g5138, g7810;
wire g7363, I9099, g9151, g6525, g6710, I6209, g8904, g5707, I14980, g9010, g5201;
wire g8763, I9044, g8637, g5715, g9282, I15040, g5052, I15252, g7782, g6931, I14969;
wire g5070, g2213, g8982, g4055, g8128, I11603, g9264, g6440, g6123, I15051, I15072;
wire I14496, g8902, I15152, g8155, g8964, g5227, I15020, g5203, I9029, g8989, I15113;
wire g8834, g5188, g7435, g7690, g5216, g3131, g8909, g4734, g6933, I14480, g9285;
wire I6208, g5217, g9139, g9339, g5711, g7222, I14942, g4688, g5196, g6132, g8985;
wire g7089, g5256, I14468, g8794, g5021, g7254, g6600, g8905, g7438, g6580, g6262;
wire I15229, I14479, I15228, g4072, g9135, g9288, I15112, g5673, g7062, g4413, g8884;
wire g7788, g8988, g6926, g8804, g9054, I15298, g6543, g8908, I14772, I15232, I15261;
wire g6927, g9171, g8965, g5220, g6436, g8996, g9138, g9338, g8777, g9049, I15031;
wire g8981, g1690, g8997, g6579, g7088, g6719, g6917, g9162, g4735, g9052, g5210;
wire g2262, I15043, g7825, g3760, I9041, g5317, I14952, g6706, g7230, g9006, g8889;
wire I14834, g7337, g6138, I15086, g6707, g8795, g7248, g1955, g5704, g9007, g7081;
wire g9261, g8634, I15017, g7783, g8613, g8983, g4876, g6728, g6470, g8885, I7232;
wire g9165, I15042, g9055, g6445, g7258, g6602, g4295, I15030, g6920, g5561, g6459;
wire g6718, g7026, I14933, g7426, g7170, g7083, I15075, g8990, g8888, g7191, g5244;
wire g5140, g7016, g9168, I15276, I15285, g5214, I15053, I15254, g4249, g3986, I14302;
wire g9011, I15101, g5236, g7272, g8896, g5222, g4812, g4829, g6685, g5237, I15074;
wire I15239, g5194, g9000, g8897, g7166, g5242, g5254, I14932, g6585, g6673, g5212;
wire g7167, g8091, I15083, g5229, I15284, g6458, g7834, g6734, g4870, g7687, g6688;
wire I15052, I14959, g5708, g5219, g6924, I15400, g9294, g8758, g9356, g7020, I15241;
wire I15100, g9363, g6116, g6565, g8994, g5245, g9357, g3192, g4727, g7040, g5259;
wire I14831, I9038, I15082, g5215, I14753, g2368, g4747, I13220, I15263, g6739, I5757;
wire I8363, I14960, g5228, g5230, g8890, I15273, g5195, g9004, g7202, I15033, g8992;
wire I14970, g4280, g6912, g5255, g4790, g6929, g7450, g1872, g5218, g6735, g5830;
wire I15291, I7233, g5221, I15029, g2043, g8999, g8146, I8224, g5716, g6919, g9002;
wire g6952, I15240, I14495, g5241, I14985, g3097, I15262, g6925, g6120, g5211, g6906;
wire I15099, I15098, I15251, I15272, g5483, I15032, g6907, g9009, g8995, I14219, g5200;
wire g5345, g5223, I15071, I14467, I15147, g6590, I15172, g6928, g6930, g5537, g7436;
wire g5243, g5234, I15044, g6705, g8894, g8782, g9005, g5213, I15290, g4374, g8998;
wire g9124, g5698, I14485, g5260, g9377, g6921, g8986, I15297, I15888, I7466, I10092;
wire g5686, I5521, g4528, g5625, I7538, I11143, I7467, g4839, I10906, I12575, I7181;
wire g4235, g6286, I7421, g5141, g6911, g4548, I15855, I11110, I11179, g6473, I6524;
wire I11178, I8510, I8245, g4313, I11186, g6469, I13685, I6258, g6177, I13800, I15819;
wire I15818, I5600, g6287, I9978, I9243, I6274, g5284, I10745, g5239, I9234, I6170;
wire I13587, g6510, I6939, I11117, g5559, g3232, I7531, g3938, I7505, I7011, I11123;
wire I11751, g6701, g4835, I13639, I10329, g6215, I6904, I13638, I10328, g5750, I7480;
wire I11841, I7569, I9964, g3525, g4332, g7535, I6757, I12051, g3358, I11116, I11615;
wire I6522, I9057, I10991, I9549, I8255, g4492, g4714, I11142, I7423, I11165, I6234;
wire I10744, g5555, I10849, g4889, g4476, g6142, I10848, g4871, g6497, I7240, g5567;
wire I10361, I7443, I13600, I9691, g6218, g4231, I11137, I7533, I11873, I12552, I9985;
wire I11614, g7093, g9191, I6843, I8119, I11122, I8152, I7460, I14473, I10789, I7937;
wire I11136, I6232, I7479, I10359, I6813, g1759, g5558, I6740, g4513, I11164, I8939;
wire g6119, g7257, I7156, g4679, I11575, g3518, I8636, g4831, I11109, g6893, I11108;
wire g6274, I9151, I7453, g6170, I11750, I7568, g6280, I7157, I8637, g4869, I8536;
wire I9278, g3658, g6187, I6275, I9235, I10981, g2395, I9693, I9548, g7480, I10899;
wire g1678, I11757, g5672, g6695, g3680, g1682, g6159, I8537, I13397, I6905, I8243;
wire I8328, g2783, I9965, I6750, I13213, g5712, g4745, I11574, g4309, I10061, I7616;
wire I8512, g3889, I10360, I8166, I7503, g3722, g4575, I15863, I13396, I14472, I14246;
wire I7277, I10071, I6172, I7617, g6902, I9153, g7316, g3231, I6134, I12080, I7892;
wire I8393, g1910, I13787, I12031, g5632, g5095, g4881, g2352, I7140, g6463, I7478;
wire I8121, I6202, I13640, g3613, g5752, I12869, I8253, I8938, I6776, I8606, I7214;
wire g4305, I9476, I13003, I6996, g5189, I13786, I6878, g3679, I8607, I8659, I9477;
wire g4227, I6997, I12079, g6570, I12078, I12598, I10889, I10980, I10888, g2315, g4502;
wire g6158, g5575, I11149, I8559, g6275, g6615, I7150, g5539, I7438, I7009, I15862;
wire I12017, g6284, g6180, g4741, I9946, g4910, I10625, g2330, g6559, g3012, g9202;
wire g3706, I9182, I9382, I10060, I10197, I6500, I10855, I8151, I13378, I9947, I11096;
wire I10867, I5505, I13802, I10315, g5305, I6523, I10819, I12016, I10818, g5748, I11549;
wire g9179, I7085, I7485, I6104, I6499, g4256, I8134, g7503, I10094, I6273, g2367;
wire g4700, I13002, I9233, I10019, g4263, I10196, I10018, g6282, I10866, I7270, I10001;
wire I7610, I9171, I10923, I7069, I10300, g7244, I7540, g7140, g5689, I9745, I9963;
wire g7082, I6135, g3678, I15881, I11080, I10854, I6916, g5564, I8658, I5696, I7510;
wire I12853, g4474, I10314, I6102, I11843, I10307, g5589, I8132, I8680, g3602, I6752;
wire I6917, g1775, I7215, g3767, I5697, I8558, I12053, I6233, I10335, g9205, I8511;
wire I10993, I14839, g5538, I15897, I14838, g7237, I9070, g6153, g6680, g8239, I11171;
wire I6171, I10039, I10306, I10038, g3028, I11079, I7891, I10143, I13599, I11078, I13598;
wire g5562, I10791, I15850, I8339, g5257, I6759, g5605, g3883, I11158, I6201, I9169;
wire g5751, I9059, g6476, I11144, I9767, g6722, I10223, g6285, I12577, I6539, I10321;
wire I13017, g6424, I10953, I15857, g6477, g4820, I10334, I13687, I11752, I7068, I12852;
wire I7468, g6273, I9826, I8660, I10000, I10908, I11842, I7576, I7149, I12576, I13016;
wire g4294, I8679, I7241, I12052, I15856, I15880, I10992, I9827, g7069, I11124, I8560;
wire g4954, g4810, g7540, g4363, I13686, I9196, I10835, g6178, I7893, I7186, I11875;
wire g4912, g3890, I9994, g3011, I7939, I6203, I9181, g5753, I8164, I9381, I15887;
wire g7144, I10142, I6940, I7187, I7461, g5565, g5681, g6265, g5697, I11170, g6164;
wire I8956, I6741, g6770, I13589, I13588, I8338, g3924, I10952, I6758, I6066, g7065;
wire I11616, I10790, I9058, I10873, I8957, g3665, I6133, g6281, I6774, I11101, I11177;
wire I10834, I6538, I9992, I11874, I15817, I12833, I10320, I10073, g8231, g5363, g3681;
wire I8504, g3914, I12951, g5568, I12033, I8470, I7512, g9203, I11185, g4244, I6257;
wire I7148, I9183, I9383, I14474, I8678, I10327, g7828, I8635, I6751, g6504, I13215;
wire g2378, I10982, I7279, I9999, g4110, g4310, g4824, g5661, I8582, I7938, I5620;
wire I10040, g8798, g4563, g6169, g6283, g4237, I11576, I8502, I10847, I8940, I10062;
wire I11115, g5546, g7325, I5520, g6203, I11184, I7158, I6924, I12832, I10072, g4836;
wire g3894, g6188, I7174, I13214, I10820, I7239, I8165, I7180, I6103, I8133, g1819;
wire I12032, g5035, I9954, I8538, I15864, I12871, g6466, g7447, g6165, g6571, g5310;
wire g4298, I10743, g5762, g3925, g5590, I11759, g5657, I11758, g6467, g5556, g4219;
wire g2385, g7234, g4252, g3906, I6775, I7010, I10890, I8605, g6181, g4911, I9475;
wire I6739, I7172, I7278, I11135, I7618, g2801, g5557, g3907, I6501, I13004, I9276;
wire g3656, g3915, g4399, I9986, I7567, I9277, I11163, I12551, g7121, I9987, g3899;
wire I9547, I7179, I8326, I12181, I10011, I7611, I10627, g4887, g4228, I10925, I6998;
wire I8327, g6023, I7511, g2333, I8472, I7574, g9190, I12870, I6925, I13395, g5540;
wire I10626, I14245, I10299, g3895, I10298, g6472, I6906, I5599, I9194, I10856, I15882;
wire I7139, I9071, I9242, g5291, I9948, I8581, I9955, g2751, I6876, I9769, I10080;
wire I10924, I15849, g3286, I15848, I9993, I12597, I5695, I7444, I7269, I10198, g5594;
wire I13785, I6877, I10868, g2474, I12854, I10225, I11151, I11172, I6064, g4893, g5550;
wire I14244, g3900, g6163, I7436, I12550, g4821, I6844, I12596, I7422, I13377, I12180;
wire I10010, g3886, I6814, I10079, I7437, g3314, I10078, g5312, I10322, g2051, I10901;
wire I6918, I9980, I9069, I8583, g4359, I10144, I11551, g3887, I7454, I10336, g6627;
wire I7532, I10017, I5619, I13376, I11103, I11095, g8633, I8503, g4880, g5576, I10224;
wire I7429, I8120, I12015, I5598, g6276, g4243, g5747, I6842, I7138, I10954, I6941;
wire g6503, I5519, I12179, g8681, I15899, I15898, I12953, I8244, g6277, I7575, I8340;
wire g4090, I9768, g6516, g3129, g4456, I7539, g2995, g2294, g3221, I7268, I5506;
wire I7452, g6709, I6540, I10093, I9195, I7086, I7486, g6435, g6482, I7504, I10875;
wire I7070, I14837, g4686, I11094, I5507, I11150, I13801, I9692, g7444, I13018, I6259;
wire I7087, I7487, I6923, g3818, I8394, I9979, g3893, I7445, I7173, I8471, I9828;
wire g5595, I8955, g9192, I8254, I10836, I9746, I7459, I11102, I11157, g3939, I8150;
wire g3083, I9953, g4879, I10313, I6065, I10305, I10900, I9747, g8627, I11550, I9241;
wire g5512, I7188, I10874, I7216, I12952, I7428, I10009, I7430, I11156, I9152, I5621;
wire I6815, g4905, g3811, g3315, I10907, I7609, I12834, I8392, I9170, I15889, g4884;
wire g8656, g3260, g5615, g8236, g4160, g7406, g6259, g6465, g3515, g8812, g3528;
wire g8073, g3555, g8819, g8694, g8806, g8230, g8807, g4888, g8859, g7326, g8699;
wire g8855, g8644, g6193, g8818, g3885, g6174, g3233, g8811, g8629, g8279, g3504;
wire g8625, g8232, g8659, g6209, g8630, g6184, g8655, g5772, g2521, g7324, g5023;
wire g8360, g8641, g3505, g8658, g8680, g4894, g7314, g8092, g7322, g8523, g7312;
wire g6452, g2014, g8862, g6185, g8679, g5039, g8805, g7152, g6664, g1980, g8233;
wire g8706, g6910, g8707, g7328, g3516, g6197, g8635, g8801, g3310, g7318, g7321;
wire g3237, g8861, g4354, g8803, g4676, g8847, g4349, g3225, g7566, g8863, g1964;
wire g7209, g5614, g4318, g6214, g4232, g6489, g3790, g5056, g8850;
wire line1, line2, line3, line4, line5, line6, line7, line8, line9, line10, line11;
wire line12, line13, line14, line15, line16, line17, line18, line19, line20, line21, line22;
wire line23, line24, line25, line26, line27, line28, line29, line30, line31, line32, line33;
wire line34, line35, line36, line37, line38, line39, line40, line41, line42, line43, line44;
wire line45, line46, line47, line48, line49, line50, line51, line52, line53, line54, line55;
wire line56, line57, line58, line59, line60, line61, line62, line63, line64, line65, line66;
wire line67, line68, line69, line70, line71, line72, line73, line74, line75, line76, line77;
wire line78, line79, line80, line81, line82, line83, line84, line85, line86, line87, line88;
wire line89, line90, line91, line92, line93, line94, line95, line96, line97, line98, line99;
wire line100, line101, line102, line103, line104, line105, line106, line107, line108, line109, line110;
wire line111, line112, line113, line114, line115, line116, line117, line118, line119, line120, line121;
wire line122, line123, line124, line125, line126, line127, line128, line129, line130, line131, line132;
wire line133, line134, line135, line136, line137, line138, line139, line140, line141, line142, line143;
wire line144, line145, line146, line147, line148, line149, line150, line151, line152, line153, line154;
wire line155, line156, line157, line158, line159, line160, line161, line162, line163, line164, line165;
wire line166, line167, line168, line169, line170, line171, line172, line173, line174, line175, line176;
wire line177, line178, line179, line180, line181, line182, line183, line184, line185, line186, line187;
wire line188, line189, line190, line191, line192, line193, line194, line195, line196, line197, line198;
wire line199, line200, line201, line202, line203, line204, line205, line206, line207, line208, line209;
wire line210, line211, line212, line213, line214, line215, line216, line217, line218, line219, line220;
wire line221, line222, line223, line224, line225, line226, line227, line228, line229, line230, line231;
wire line232, line233, line234, line235, line236, line237, line238, line239, line240, line241, line242;
wire line243, line244, line245, line246, line247, line248, line249, line250, line251, line252, line253;
wire line254, line255, line256, line257, line258, line259, line260, line261, line262, line263, line264;
wire line265, line266, line267, line268, line269, line270, line271, line272, line273, line274, line275;
wire line276, line277, line278, line279, line280, line281, line282, line283, line284, line285, line286;
wire line287, line288, line289, line290, line291, line292, line293, line294, line295, line296, line297;
wire line298, line299, line300, line301, line302, line303, line304, line305, line306, line307, line308;
wire line309, line310, line311, line312, line313, line314, line315, line316, line317, line318, line319;
wire line320, line321, line322, line323, line324, line325, line326, line327, line328, line329, line330;
wire line331, line332, line333, line334, line335, line336, line337, line338, line339, line340, line341;
wire line342, line343, line344, line345, line346, line347, line348, line349, line350, line351, line352;
wire line353, line354, line355, line356, line357, line358, line359, line360, line361, line362, line363;
wire line364, line365, line366, line367, line368, line369, line370, line371, line372, line373, line374;
wire line375, line376, line377, line378, line379, line380, line381, line382, line383, line384, line385;
wire line386, line387, line388, line389, line390, line391, line392, line393, line394, line395, line396;
wire line397, line398, line399, line400, line401, line402, line403, line404, line405, line406, line407;
wire line408, line409, line410, line411, line412, line413, line414, line415, line416, line417, line418;
wire line419, line420, line421, line422, line423, line424, line425, line426, line427, line428, line429;
wire line430, line431, line432, line433, line434, line435, line436, line437, line438, line439, line440;
wire line441, line442, line443, line444, line445, line446, line447, line448, line449, line450, line451;
wire line452, line453, line454, line455, line456, line457, line458, line459, line460, line461, line462;
wire line463, line464, line465, line466, line467, line468, line469, line470, line471, line472, line473;
wire line474, line475, line476, line477, line478, line479, line480, line481, line482, line483, line484;
wire line485, line486, line487, line488, line489, line490, line491, line492, line493, line494, line495;
wire line496, line497, line498, line499, line500, line501, line502, line503, line504, line505, line506;
wire line507, line508, line509, line510, line511, line512, line513, line514, line515, line516, line517;
wire line518, line519, line520, line521, line522, line523, line524, line525, line526, line527, line528;
wire line529, line530, line531, line532, line533, line534, line535, line536, line537, line538, line539;
wire line540, line541, line542, line543, line544, line545, line546, line547, line548, line549, line550;
wire line551, line552, line553, line554, line555, line556, line557, line558, line559, line560, line561;
wire line562, line563, line564, line565, line566, line567, line568, line569, line570, line571, line572;
wire line573, line574, line575, line576, line577, line578, line579, line580, line581, line582, line583;
wire line584, line585, line586, line587, line588, line589, line590, line591, line592, line593, line594;
wire line595, line596, line597, line598, line599, line600, line601, line602, line603, line604, line605;
wire line606, line607, line608, line609, line610, line611, line612, line613, line614, line615, line616;
wire line617, line618, line619, line620, line621, line622, line623, line624, line625, line626, line627;
wire line628, line629, line630, line631, line632, line633, line634, line635, line636, line637, line638;
DFFX1 gate1(.Q (g397), .QB (line1), .D(g4635), .CK(clk));
DFFX1 gate2(.Q (g1271), .QB (line2), .D(g5176), .CK(clk));
DFFX1 gate3(.Q (g312), .QB (line3), .D(g4618), .CK(clk));
DFFX1 gate4(.Q (g273), .QB (line4), .D(g4611), .CK(clk));
DFFX1 gate5(.Q (g452), .QB (line5), .D(g449), .CK(clk));
DFFX1 gate6(.Q (g948), .QB (line6), .D(g8664), .CK(clk));
DFFX1 gate7(.Q (g629), .QB (line7), .D(g6827), .CK(clk));
DFFX1 gate8(.Q (g207), .QB (line8), .D(g5733), .CK(clk));
DFFX1 gate9(.Q (g1541), .QB (line9), .D(g7778), .CK(clk));
DFFX1 gate10(.Q (g1153), .QB (line10), .D(g6856), .CK(clk));
DFFX1 gate11(.Q (g940), .QB (line11), .D(g5735), .CK(clk));
DFFX1 gate12(.Q (g976), .QB (line12), .D(g8864), .CK(clk));
DFFX1 gate13(.Q (g498), .QB (line13), .D(g9111), .CK(clk));
DFFX1 gate14(.Q (g314), .QB (line14), .D(g4620), .CK(clk));
DFFX1 gate15(.Q (g1092), .QB (line15), .D(g7520), .CK(clk));
DFFX1 gate16(.Q (g454), .QB (line16), .D(g4639), .CK(clk));
DFFX1 gate17(.Q (g196), .QB (line17), .D(g5731), .CK(clk));
DFFX1 gate18(.Q (g535), .QB (line18), .D(g3844), .CK(clk));
DFFX1 gate19(.Q (g292), .QB (line19), .D(g4613), .CK(clk));
DFFX1 gate20(.Q (g772), .QB (line20), .D(g6846), .CK(clk));
DFFX1 gate21(.Q (g1375), .QB (line21), .D(g6869), .CK(clk));
DFFX1 gate22(.Q (g689), .QB (line22), .D(g6371), .CK(clk));
DFFX1 gate23(.Q (g183), .QB (line23), .D(g6309), .CK(clk));
DFFX1 gate24(.Q (g359), .QB (line24), .D(g6336), .CK(clk));
DFFX1 gate25(.Q (g1384), .QB (line25), .D(g6881), .CK(clk));
DFFX1 gate26(.Q (g1339), .QB (line26), .D(g6865), .CK(clk));
DFFX1 gate27(.Q (g20), .QB (line27), .D(g6386), .CK(clk));
DFFX1 gate28(.Q (g1424), .QB (line28), .D(g3862), .CK(clk));
DFFX1 gate29(.Q (g767), .QB (line29), .D(g6841), .CK(clk));
DFFX1 gate30(.Q (g393), .QB (line30), .D(g4631), .CK(clk));
DFFX1 gate31(.Q (g1077), .QB (line31), .D(g7767), .CK(clk));
DFFX1 gate32(.Q (g1231), .QB (line32), .D(g1236), .CK(clk));
DFFX1 gate33(.Q (g294), .QB (line33), .D(g4615), .CK(clk));
DFFX1 gate34(.Q (g1477), .QB (line34), .D(g9036), .CK(clk));
DFFX1 gate35(.Q (g4), .QB (line35), .D(g9372), .CK(clk));
DFFX1 gate36(.Q (g608), .QB (line36), .D(g6806), .CK(clk));
DFFX1 gate37(.Q (g1205), .QB (line37), .D(g1204), .CK(clk));
DFFX1 gate38(.Q (g465), .QB (line38), .D(g6352), .CK(clk));
DFFX1 gate39(.Q (g774), .QB (line39), .D(g6848), .CK(clk));
DFFX1 gate40(.Q (g921), .QB (line40), .D(g916), .CK(clk));
DFFX1 gate41(.Q (g1304), .QB (line41), .D(g1312), .CK(clk));
DFFX1 gate42(.Q (g243), .QB (line42), .D(g6318), .CK(clk));
DFFX1 gate43(.Q (g1499), .QB (line43), .D(g7772), .CK(clk));
DFFX1 gate44(.Q (g80), .QB (line44), .D(g6778), .CK(clk));
DFFX1 gate45(.Q (g1444), .QB (line45), .D(g5185), .CK(clk));
DFFX1 gate46(.Q (g1269), .QB (line46), .D(g5740), .CK(clk));
DFFX1 gate47(.Q (g600), .QB (line47), .D(g6807), .CK(clk));
DFFX1 gate48(.Q (g423), .QB (line48), .D(g9105), .CK(clk));
DFFX1 gate49(.Q (g771), .QB (line49), .D(g6845), .CK(clk));
DFFX1 gate50(.Q (g803), .QB (line50), .D(g7757), .CK(clk));
DFFX1 gate51(.Q (g843), .QB (line51), .D(g2647), .CK(clk));
DFFX1 gate52(.Q (g315), .QB (line52), .D(g4621), .CK(clk));
DFFX1 gate53(.Q (g455), .QB (line53), .D(g4640), .CK(clk));
DFFX1 gate54(.Q (g906), .QB (line54), .D(g901), .CK(clk));
DFFX1 gate55(.Q (g622), .QB (line55), .D(g6821), .CK(clk));
DFFX1 gate56(.Q (g891), .QB (line56), .D(g3855), .CK(clk));
DFFX1 gate57(.Q (g1014), .QB (line57), .D(g1012), .CK(clk));
DFFX1 gate58(.Q (g984), .QB (line58), .D(g9133), .CK(clk));
DFFX1 gate59(.Q (g117), .QB (line59), .D(g5153), .CK(clk));
DFFX1 gate60(.Q (g137), .QB (line60), .D(g5150), .CK(clk));
DFFX1 gate61(.Q (g527), .QB (line61), .D(g9110), .CK(clk));
DFFX1 gate62(.Q (g1513), .QB (line62), .D(g1524), .CK(clk));
DFFX1 gate63(.Q (g278), .QB (line63), .D(g6323), .CK(clk));
DFFX1 gate64(.Q (g1378), .QB (line64), .D(g6880), .CK(clk));
DFFX1 gate65(.Q (g718), .QB (line65), .D(g7753), .CK(clk));
DFFX1 gate66(.Q (g598), .QB (line66), .D(g6797), .CK(clk));
DFFX1 gate67(.Q (g1182), .QB (line67), .D(g1160), .CK(clk));
DFFX1 gate68(.Q (g1288), .QB (line68), .D(g7527), .CK(clk));
DFFX1 gate69(.Q (g1382), .QB (line69), .D(g6888), .CK(clk));
DFFX1 gate70(.Q (g179), .QB (line70), .D(g5159), .CK(clk));
DFFX1 gate71(.Q (g624), .QB (line71), .D(g6831), .CK(clk));
DFFX1 gate72(.Q (g48), .QB (line72), .D(g9362), .CK(clk));
DFFX1 gate73(.Q (g362), .QB (line73), .D(g9093), .CK(clk));
DFFX1 gate74(.Q (g878), .QB (line74), .D(g890), .CK(clk));
DFFX1 gate75(.Q (g270), .QB (line75), .D(g9092), .CK(clk));
DFFX1 gate76(.Q (g763), .QB (line76), .D(g6836), .CK(clk));
DFFX1 gate77(.Q (g710), .QB (line77), .D(g7751), .CK(clk));
DFFX1 gate78(.Q (g730), .QB (line78), .D(g7754), .CK(clk));
DFFX1 gate79(.Q (g295), .QB (line79), .D(g4616), .CK(clk));
DFFX1 gate80(.Q (g1037), .QB (line80), .D(g7519), .CK(clk));
DFFX1 gate81(.Q (g1102), .QB (line81), .D(g6855), .CK(clk));
DFFX1 gate82(.Q (g483), .QB (line82), .D(g6356), .CK(clk));
DFFX1 gate83(.Q (g775), .QB (line83), .D(g7759), .CK(clk));
DFFX1 gate84(.Q (g621), .QB (line84), .D(g6819), .CK(clk));
DFFX1 gate85(.Q (g1364), .QB (line85), .D(g6878), .CK(clk));
DFFX1 gate86(.Q (g1454), .QB (line86), .D(g5187), .CK(clk));
DFFX1 gate87(.Q (g1296), .QB (line87), .D(g7304), .CK(clk));
DFFX1 gate88(.Q (g5), .QB (line88), .D(g9373), .CK(clk));
DFFX1 gate89(.Q (g1532), .QB (line89), .D(g7781), .CK(clk));
DFFX1 gate90(.Q (g587), .QB (line90), .D(g3852), .CK(clk));
DFFX1 gate91(.Q (g741), .QB (line91), .D(g9386), .CK(clk));
DFFX1 gate92(.Q (g13), .QB (line92), .D(g7308), .CK(clk));
DFFX1 gate93(.Q (g606), .QB (line93), .D(g6804), .CK(clk));
DFFX1 gate94(.Q (g1012), .QB (line94), .D(g6851), .CK(clk));
DFFX1 gate95(.Q (g52), .QB (line95), .D(g6781), .CK(clk));
DFFX1 gate96(.Q (g646), .QB (line96), .D(g4652), .CK(clk));
DFFX1 gate97(.Q (g1412), .QB (line97), .D(g5745), .CK(clk));
DFFX1 gate98(.Q (g327), .QB (line98), .D(g6332), .CK(clk));
DFFX1 gate99(.Q (g1189), .QB (line99), .D(g6392), .CK(clk));
DFFX1 gate100(.Q (g1389), .QB (line100), .D(g4658), .CK(clk));
DFFX1 gate101(.Q (g1029), .QB (line101), .D(g2654), .CK(clk));
DFFX1 gate102(.Q (g1371), .QB (line102), .D(g6868), .CK(clk));
DFFX1 gate103(.Q (g1429), .QB (line103), .D(g2671), .CK(clk));
DFFX1 gate104(.Q (g398), .QB (line104), .D(g4636), .CK(clk));
DFFX1 gate105(.Q (g985), .QB (line105), .D(g7515), .CK(clk));
DFFX1 gate106(.Q (g354), .QB (line106), .D(g4624), .CK(clk));
DFFX1 gate107(.Q (g619), .QB (line107), .D(g6817), .CK(clk));
DFFX1 gate108(.Q (g113), .QB (line108), .D(g5148), .CK(clk));
DFFX1 gate109(.Q (g133), .QB (line109), .D(g5149), .CK(clk));
DFFX1 gate110(.Q (g180), .QB (line110), .D(g5158), .CK(clk));
DFFX1 gate111(.Q (g1138), .QB (line111), .D(g7524), .CK(clk));
DFFX1 gate112(.Q (g1309), .QB (line112), .D(g1308), .CK(clk));
DFFX1 gate113(.Q (g889), .QB (line113), .D(g7101), .CK(clk));
DFFX1 gate114(.Q (g390), .QB (line114), .D(g6341), .CK(clk));
DFFX1 gate115(.Q (g625), .QB (line115), .D(g6823), .CK(clk));
DFFX1 gate116(.Q (g417), .QB (line116), .D(g9103), .CK(clk));
DFFX1 gate117(.Q (g681), .QB (line117), .D(g7748), .CK(clk));
DFFX1 gate118(.Q (g437), .QB (line118), .D(g6348), .CK(clk));
DFFX1 gate119(.Q (g351), .QB (line119), .D(g9100), .CK(clk));
DFFX1 gate120(.Q (g1201), .QB (line120), .D(g1200), .CK(clk));
DFFX1 gate121(.Q (g109), .QB (line121), .D(g6785), .CK(clk));
DFFX1 gate122(.Q (g1049), .QB (line122), .D(g8673), .CK(clk));
DFFX1 gate123(.Q (g1098), .QB (line123), .D(g6854), .CK(clk));
DFFX1 gate124(.Q (g200), .QB (line124), .D(g199), .CK(clk));
DFFX1 gate125(.Q (g240), .QB (line125), .D(g6317), .CK(clk));
DFFX1 gate126(.Q (g479), .QB (line126), .D(g4649), .CK(clk));
DFFX1 gate127(.Q (g126), .QB (line127), .D(g6789), .CK(clk));
DFFX1 gate128(.Q (g596), .QB (line128), .D(g6795), .CK(clk));
DFFX1 gate129(.Q (g1268), .QB (line129), .D(g5175), .CK(clk));
DFFX1 gate130(.Q (g222), .QB (line130), .D(g6313), .CK(clk));
DFFX1 gate131(.Q (g420), .QB (line131), .D(g9104), .CK(clk));
DFFX1 gate132(.Q (g3), .QB (line132), .D(g9360), .CK(clk));
DFFX1 gate133(.Q (g58), .QB (line133), .D(g7734), .CK(clk));
DFFX1 gate134(.Q (g172), .QB (line134), .D(g1270), .CK(clk));
DFFX1 gate135(.Q (g387), .QB (line135), .D(g6340), .CK(clk));
DFFX1 gate136(.Q (g840), .QB (line136), .D(g2648), .CK(clk));
DFFX1 gate137(.Q (g365), .QB (line137), .D(g9094), .CK(clk));
DFFX1 gate138(.Q (g1486), .QB (line138), .D(g8226), .CK(clk));
DFFX1 gate139(.Q (g1504), .QB (line139), .D(g7773), .CK(clk));
DFFX1 gate140(.Q (g1185), .QB (line140), .D(g1155), .CK(clk));
DFFX1 gate141(.Q (g1385), .QB (line141), .D(g6883), .CK(clk));
DFFX1 gate142(.Q (g583), .QB (line142), .D(g3851), .CK(clk));
DFFX1 gate143(.Q (g822), .QB (line143), .D(g7512), .CK(clk));
DFFX1 gate144(.Q (g1025), .QB (line144), .D(g8871), .CK(clk));
DFFX1 gate145(.Q (g969), .QB (line145), .D(g966), .CK(clk));
DFFX1 gate146(.Q (g768), .QB (line146), .D(g6842), .CK(clk));
DFFX1 gate147(.Q (g174), .QB (line147), .D(g7737), .CK(clk));
DFFX1 gate148(.Q (g685), .QB (line148), .D(g7749), .CK(clk));
DFFX1 gate149(.Q (g1087), .QB (line149), .D(g6853), .CK(clk));
DFFX1 gate150(.Q (g355), .QB (line150), .D(g4625), .CK(clk));
DFFX1 gate151(.Q (g911), .QB (line151), .D(g906), .CK(clk));
DFFX1 gate152(.Q (g1226), .QB (line152), .D(g6859), .CK(clk));
DFFX1 gate153(.Q (g99), .QB (line153), .D(g6783), .CK(clk));
DFFX1 gate154(.Q (g1045), .QB (line154), .D(g8224), .CK(clk));
DFFX1 gate155(.Q (g1173), .QB (line155), .D(g7526), .CK(clk));
DFFX1 gate156(.Q (g1373), .QB (line156), .D(g6871), .CK(clk));
DFFX1 gate157(.Q (g186), .QB (line157), .D(g3830), .CK(clk));
DFFX1 gate158(.Q (g760), .QB (line158), .D(g6833), .CK(clk));
DFFX1 gate159(.Q (g959), .QB (line159), .D(g5169), .CK(clk));
DFFX1 gate160(.Q (g1369), .QB (line160), .D(g6875), .CK(clk));
DFFX1 gate161(.Q (g1007), .QB (line161), .D(g8867), .CK(clk));
DFFX1 gate162(.Q (g1459), .QB (line162), .D(g3863), .CK(clk));
DFFX1 gate163(.Q (g758), .QB (line163), .D(g6840), .CK(clk));
DFFX1 gate164(.Q (g480), .QB (line164), .D(g6355), .CK(clk));
DFFX1 gate165(.Q (g396), .QB (line165), .D(g4634), .CK(clk));
DFFX1 gate166(.Q (g612), .QB (line166), .D(g6811), .CK(clk));
DFFX1 gate167(.Q (g38), .QB (line167), .D(g5746), .CK(clk));
DFFX1 gate168(.Q (g632), .QB (line168), .D(g6830), .CK(clk));
DFFX1 gate169(.Q (g1415), .QB (line169), .D(g5180), .CK(clk));
DFFX1 gate170(.Q (g1227), .QB (line170), .D(g7108), .CK(clk));
DFFX1 gate171(.Q (g246), .QB (line171), .D(g6319), .CK(clk));
DFFX1 gate172(.Q (g449), .QB (line172), .D(g3840), .CK(clk));
DFFX1 gate173(.Q (g517), .QB (line173), .D(g4651), .CK(clk));
DFFX1 gate174(.Q (g118), .QB (line174), .D(g6787), .CK(clk));
DFFX1 gate175(.Q (g138), .QB (line175), .D(g6792), .CK(clk));
DFFX1 gate176(.Q (g16), .QB (line176), .D(g1404), .CK(clk));
DFFX1 gate177(.Q (g284), .QB (line177), .D(g9086), .CK(clk));
DFFX1 gate178(.Q (g142), .QB (line178), .D(g6793), .CK(clk));
DFFX1 gate179(.Q (g219), .QB (line179), .D(g6312), .CK(clk));
DFFX1 gate180(.Q (g426), .QB (line180), .D(g9106), .CK(clk));
DFFX1 gate181(.Q (g1388), .QB (line181), .D(g6882), .CK(clk));
DFFX1 gate182(.Q (g806), .QB (line182), .D(g7510), .CK(clk));
DFFX1 gate183(.Q (g846), .QB (line183), .D(g2646), .CK(clk));
DFFX1 gate184(.Q (g1428), .QB (line184), .D(g2672), .CK(clk));
DFFX1 gate185(.Q (g579), .QB (line185), .D(g3850), .CK(clk));
DFFX1 gate186(.Q (g1030), .QB (line186), .D(g7518), .CK(clk));
DFFX1 gate187(.Q (g614), .QB (line187), .D(g6812), .CK(clk));
DFFX1 gate188(.Q (g1430), .QB (line188), .D(g4666), .CK(clk));
DFFX1 gate189(.Q (g1247), .QB (line189), .D(g6380), .CK(clk));
DFFX1 gate190(.Q (g669), .QB (line190), .D(g7745), .CK(clk));
DFFX1 gate191(.Q (g110), .QB (line191), .D(g109), .CK(clk));
DFFX1 gate192(.Q (g130), .QB (line192), .D(g6790), .CK(clk));
DFFX1 gate193(.Q (g225), .QB (line193), .D(g6314), .CK(clk));
DFFX1 gate194(.Q (g281), .QB (line194), .D(g9085), .CK(clk));
DFFX1 gate195(.Q (g819), .QB (line195), .D(g7761), .CK(clk));
DFFX1 gate196(.Q (g1308), .QB (line196), .D(g6385), .CK(clk));
DFFX1 gate197(.Q (g611), .QB (line197), .D(g6810), .CK(clk));
DFFX1 gate198(.Q (g631), .QB (line198), .D(g6829), .CK(clk));
DFFX1 gate199(.Q (g1217), .QB (line199), .D(g6377), .CK(clk));
DFFX1 gate200(.Q (g104), .QB (line200), .D(g6784), .CK(clk));
DFFX1 gate201(.Q (g1365), .QB (line201), .D(g6867), .CK(clk));
DFFX1 gate202(.Q (g825), .QB (line202), .D(g7513), .CK(clk));
DFFX1 gate203(.Q (g1333), .QB (line203), .D(g6863), .CK(clk));
DFFX1 gate204(.Q (g474), .QB (line204), .D(g4644), .CK(clk));
DFFX1 gate205(.Q (g1396), .QB (line205), .D(g4662), .CK(clk));
DFFX1 gate206(.Q (g141), .QB (line206), .D(g5151), .CK(clk));
DFFX1 gate207(.Q (g1509), .QB (line207), .D(g7774), .CK(clk));
DFFX1 gate208(.Q (g766), .QB (line208), .D(g6839), .CK(clk));
DFFX1 gate209(.Q (g1018), .QB (line209), .D(g8869), .CK(clk));
DFFX1 gate210(.Q (g588), .QB (line210), .D(g9031), .CK(clk));
DFFX1 gate211(.Q (g1467), .QB (line211), .D(g8875), .CK(clk));
DFFX1 gate212(.Q (g317), .QB (line212), .D(g4623), .CK(clk));
DFFX1 gate213(.Q (g457), .QB (line213), .D(g4642), .CK(clk));
DFFX1 gate214(.Q (g486), .QB (line214), .D(g6357), .CK(clk));
DFFX1 gate215(.Q (g471), .QB (line215), .D(g6354), .CK(clk));
DFFX1 gate216(.Q (g1381), .QB (line216), .D(g6887), .CK(clk));
DFFX1 gate217(.Q (g1197), .QB (line217), .D(g1196), .CK(clk));
DFFX1 gate218(.Q (g513), .QB (line218), .D(g9116), .CK(clk));
DFFX1 gate219(.Q (g1397), .QB (line219), .D(g6389), .CK(clk));
DFFX1 gate220(.Q (g533), .QB (line220), .D(g530), .CK(clk));
DFFX1 gate221(.Q (g1021), .QB (line221), .D(g8870), .CK(clk));
DFFX1 gate222(.Q (g1421), .QB (line222), .D(g5179), .CK(clk));
DFFX1 gate223(.Q (g952), .QB (line223), .D(g8668), .CK(clk));
DFFX1 gate224(.Q (g1263), .QB (line224), .D(g5737), .CK(clk));
DFFX1 gate225(.Q (g580), .QB (line225), .D(g6368), .CK(clk));
DFFX1 gate226(.Q (g615), .QB (line226), .D(g6813), .CK(clk));
DFFX1 gate227(.Q (g1257), .QB (line227), .D(g5738), .CK(clk));
DFFX1 gate228(.Q (g46), .QB (line228), .D(g8955), .CK(clk));
DFFX1 gate229(.Q (g402), .QB (line229), .D(g6343), .CK(clk));
DFFX1 gate230(.Q (g998), .QB (line230), .D(g1005), .CK(clk));
DFFX1 gate231(.Q (g1041), .QB (line231), .D(g7765), .CK(clk));
DFFX1 gate232(.Q (g297), .QB (line232), .D(g6324), .CK(clk));
DFFX1 gate233(.Q (g954), .QB (line233), .D(g8670), .CK(clk));
DFFX1 gate234(.Q (g105), .QB (line234), .D(g104), .CK(clk));
DFFX1 gate235(.Q (g145), .QB (line235), .D(g5152), .CK(clk));
DFFX1 gate236(.Q (g212), .QB (line236), .D(g4601), .CK(clk));
DFFX1 gate237(.Q (g1368), .QB (line237), .D(g6874), .CK(clk));
DFFX1 gate238(.Q (g232), .QB (line238), .D(g4606), .CK(clk));
DFFX1 gate239(.Q (g990), .QB (line239), .D(g7516), .CK(clk));
DFFX1 gate240(.Q (g475), .QB (line240), .D(g4645), .CK(clk));
DFFX1 gate241(.Q (g33), .QB (line241), .D(g5184), .CK(clk));
DFFX1 gate242(.Q (g951), .QB (line242), .D(g8667), .CK(clk));
DFFX1 gate243(.Q (g799), .QB (line243), .D(g7756), .CK(clk));
DFFX1 gate244(.Q (g812), .QB (line244), .D(g7758), .CK(clk));
DFFX1 gate245(.Q (g567), .QB (line245), .D(g6367), .CK(clk));
DFFX1 gate246(.Q (g313), .QB (line246), .D(g4619), .CK(clk));
DFFX1 gate247(.Q (g333), .QB (line247), .D(g6334), .CK(clk));
DFFX1 gate248(.Q (g168), .QB (line248), .D(g7742), .CK(clk));
DFFX1 gate249(.Q (g214), .QB (line249), .D(g4603), .CK(clk));
DFFX1 gate250(.Q (g234), .QB (line250), .D(g4608), .CK(clk));
DFFX1 gate251(.Q (g652), .QB (line251), .D(g646), .CK(clk));
DFFX1 gate252(.Q (g1126), .QB (line252), .D(g8674), .CK(clk));
DFFX1 gate253(.Q (g1400), .QB (line253), .D(g6390), .CK(clk));
DFFX1 gate254(.Q (g1326), .QB (line254), .D(g7306), .CK(clk));
DFFX1 gate255(.Q (g92), .QB (line255), .D(g6794), .CK(clk));
DFFX1 gate256(.Q (g309), .QB (line256), .D(g6328), .CK(clk));
DFFX1 gate257(.Q (g211), .QB (line257), .D(g4600), .CK(clk));
DFFX1 gate258(.Q (g834), .QB (line258), .D(g2650), .CK(clk));
DFFX1 gate259(.Q (g231), .QB (line259), .D(g4605), .CK(clk));
DFFX1 gate260(.Q (g557), .QB (line260), .D(g6366), .CK(clk));
DFFX1 gate261(.Q (g1383), .QB (line261), .D(g6889), .CK(clk));
DFFX1 gate262(.Q (g1220), .QB (line262), .D(g6378), .CK(clk));
DFFX1 gate263(.Q (g158), .QB (line263), .D(g7740), .CK(clk));
DFFX1 gate264(.Q (g627), .QB (line264), .D(g6825), .CK(clk));
DFFX1 gate265(.Q (g661), .QB (line265), .D(g7743), .CK(clk));
DFFX1 gate266(.Q (g77), .QB (line266), .D(g6777), .CK(clk));
DFFX1 gate267(.Q (g831), .QB (line267), .D(g2651), .CK(clk));
DFFX1 gate268(.Q (g1327), .QB (line268), .D(g7307), .CK(clk));
DFFX1 gate269(.Q (g293), .QB (line269), .D(g4614), .CK(clk));
DFFX1 gate270(.Q (g1146), .QB (line270), .D(g1612), .CK(clk));
DFFX1 gate271(.Q (g89), .QB (line271), .D(g92), .CK(clk));
DFFX1 gate272(.Q (g150), .QB (line272), .D(g7738), .CK(clk));
DFFX1 gate273(.Q (g773), .QB (line273), .D(g6847), .CK(clk));
DFFX1 gate274(.Q (g859), .QB (line274), .D(g8221), .CK(clk));
DFFX1 gate275(.Q (g1240), .QB (line275), .D(g1235), .CK(clk));
DFFX1 gate276(.Q (g518), .QB (line276), .D(g6361), .CK(clk));
DFFX1 gate277(.Q (g1472), .QB (line277), .D(g8960), .CK(clk));
DFFX1 gate278(.Q (g1443), .QB (line278), .D(g4667), .CK(clk));
DFFX1 gate279(.Q (g436), .QB (line279), .D(g4638), .CK(clk));
DFFX1 gate280(.Q (g405), .QB (line280), .D(g6344), .CK(clk));
DFFX1 gate281(.Q (g1034), .QB (line281), .D(g8957), .CK(clk));
DFFX1 gate282(.Q (g1147), .QB (line282), .D(g1146), .CK(clk));
DFFX1 gate283(.Q (g374), .QB (line283), .D(g4627), .CK(clk));
DFFX1 gate284(.Q (g98), .QB (line284), .D(g5146), .CK(clk));
DFFX1 gate285(.Q (g563), .QB (line285), .D(g9029), .CK(clk));
DFFX1 gate286(.Q (g510), .QB (line286), .D(g9115), .CK(clk));
DFFX1 gate287(.Q (g530), .QB (line287), .D(g3842), .CK(clk));
DFFX1 gate288(.Q (g215), .QB (line288), .D(g4604), .CK(clk));
DFFX1 gate289(.Q (g235), .QB (line289), .D(g4609), .CK(clk));
DFFX1 gate290(.Q (g1013), .QB (line290), .D(g1014), .CK(clk));
DFFX1 gate291(.Q (g6), .QB (line291), .D(g9374), .CK(clk));
DFFX1 gate292(.Q (g55), .QB (line292), .D(g7733), .CK(clk));
DFFX1 gate293(.Q (g1317), .QB (line293), .D(g5743), .CK(clk));
DFFX1 gate294(.Q (g504), .QB (line294), .D(g9113), .CK(clk));
DFFX1 gate295(.Q (g665), .QB (line295), .D(g7744), .CK(clk));
DFFX1 gate296(.Q (g544), .QB (line296), .D(g6365), .CK(clk));
DFFX1 gate297(.Q (g371), .QB (line297), .D(g368), .CK(clk));
DFFX1 gate298(.Q (g62), .QB (line298), .D(g7509), .CK(clk));
DFFX1 gate299(.Q (g792), .QB (line299), .D(g5162), .CK(clk));
DFFX1 gate300(.Q (g468), .QB (line300), .D(g6353), .CK(clk));
DFFX1 gate301(.Q (g815), .QB (line301), .D(g7760), .CK(clk));
DFFX1 gate302(.Q (g1460), .QB (line302), .D(g4668), .CK(clk));
DFFX1 gate303(.Q (g553), .QB (line303), .D(g9028), .CK(clk));
DFFX1 gate304(.Q (g623), .QB (line304), .D(g6822), .CK(clk));
DFFX1 gate305(.Q (g501), .QB (line305), .D(g9112), .CK(clk));
DFFX1 gate306(.Q (g1190), .QB (line306), .D(g8677), .CK(clk));
DFFX1 gate307(.Q (g1390), .QB (line307), .D(g4659), .CK(clk));
DFFX1 gate308(.Q (g74), .QB (line308), .D(g6776), .CK(clk));
DFFX1 gate309(.Q (g1156), .QB (line309), .D(g1081), .CK(clk));
DFFX1 gate310(.Q (g318), .QB (line310), .D(g6329), .CK(clk));
DFFX1 gate311(.Q (g458), .QB (line311), .D(g4643), .CK(clk));
DFFX1 gate312(.Q (g342), .QB (line312), .D(g9097), .CK(clk));
DFFX1 gate313(.Q (g1250), .QB (line313), .D(g7111), .CK(clk));
DFFX1 gate314(.Q (g1163), .QB (line314), .D(g2655), .CK(clk));
DFFX1 gate315(.Q (g1363), .QB (line315), .D(g6877), .CK(clk));
DFFX1 gate316(.Q (g1432), .QB (line316), .D(g5183), .CK(clk));
DFFX1 gate317(.Q (g1053), .QB (line317), .D(g8873), .CK(clk));
DFFX1 gate318(.Q (g252), .QB (line318), .D(g6321), .CK(clk));
DFFX1 gate319(.Q (g330), .QB (line319), .D(g6333), .CK(clk));
DFFX1 gate320(.Q (g264), .QB (line320), .D(g9090), .CK(clk));
DFFX1 gate321(.Q (g1157), .QB (line321), .D(g1156), .CK(clk));
DFFX1 gate322(.Q (g1357), .QB (line322), .D(g8675), .CK(clk));
DFFX1 gate323(.Q (g375), .QB (line323), .D(g4628), .CK(clk));
DFFX1 gate324(.Q (g68), .QB (line324), .D(g6774), .CK(clk));
DFFX1 gate325(.Q (g852), .QB (line325), .D(g2644), .CK(clk));
DFFX1 gate326(.Q (g261), .QB (line326), .D(g9089), .CK(clk));
DFFX1 gate327(.Q (g516), .QB (line327), .D(g4650), .CK(clk));
DFFX1 gate328(.Q (g536), .QB (line328), .D(g6363), .CK(clk));
DFFX1 gate329(.Q (g979), .QB (line329), .D(g7104), .CK(clk));
DFFX1 gate330(.Q (g778), .QB (line330), .D(g7296), .CK(clk));
DFFX1 gate331(.Q (g199), .QB (line331), .D(g3832), .CK(clk));
DFFX1 gate332(.Q (g1292), .QB (line332), .D(g7302), .CK(clk));
DFFX1 gate333(.Q (g290), .QB (line333), .D(g287), .CK(clk));
DFFX1 gate334(.Q (g1084), .QB (line334), .D(g7106), .CK(clk));
DFFX1 gate335(.Q (g1439), .QB (line335), .D(g5182), .CK(clk));
DFFX1 gate336(.Q (g770), .QB (line336), .D(g6844), .CK(clk));
DFFX1 gate337(.Q (g1276), .QB (line337), .D(g6384), .CK(clk));
DFFX1 gate338(.Q (g890), .QB (line338), .D(g7102), .CK(clk));
DFFX1 gate339(.Q (g1004), .QB (line339), .D(g7105), .CK(clk));
DFFX1 gate340(.Q (g1404), .QB (line340), .D(g1403), .CK(clk));
DFFX1 gate341(.Q (g93), .QB (line341), .D(g5145), .CK(clk));
DFFX1 gate342(.Q (g2), .QB (line342), .D(g9361), .CK(clk));
DFFX1 gate343(.Q (g287), .QB (line343), .D(g3836), .CK(clk));
DFFX1 gate344(.Q (g560), .QB (line344), .D(g6370), .CK(clk));
DFFX1 gate345(.Q (g1224), .QB (line345), .D(g6857), .CK(clk));
DFFX1 gate346(.Q (g1320), .QB (line346), .D(g7114), .CK(clk));
DFFX1 gate347(.Q (g617), .QB (line347), .D(g6815), .CK(clk));
DFFX1 gate348(.Q (g316), .QB (line348), .D(g4622), .CK(clk));
DFFX1 gate349(.Q (g336), .QB (line349), .D(g9095), .CK(clk));
DFFX1 gate350(.Q (g933), .QB (line350), .D(g5166), .CK(clk));
DFFX1 gate351(.Q (g456), .QB (line351), .D(g4641), .CK(clk));
DFFX1 gate352(.Q (g345), .QB (line352), .D(g9098), .CK(clk));
DFFX1 gate353(.Q (g628), .QB (line353), .D(g6826), .CK(clk));
DFFX1 gate354(.Q (g8), .QB (line354), .D(g9376), .CK(clk));
DFFX1 gate355(.Q (g887), .QB (line355), .D(g7099), .CK(clk));
DFFX1 gate356(.Q (g789), .QB (line356), .D(g7297), .CK(clk));
DFFX1 gate357(.Q (g173), .QB (line357), .D(g7736), .CK(clk));
DFFX1 gate358(.Q (g550), .QB (line358), .D(g9027), .CK(clk));
DFFX1 gate359(.Q (g255), .QB (line359), .D(g9087), .CK(clk));
DFFX1 gate360(.Q (g949), .QB (line360), .D(g8665), .CK(clk));
DFFX1 gate361(.Q (g1244), .QB (line361), .D(g2659), .CK(clk));
DFFX1 gate362(.Q (g620), .QB (line362), .D(g6818), .CK(clk));
DFFX1 gate363(.Q (g1435), .QB (line363), .D(g5181), .CK(clk));
DFFX1 gate364(.Q (g477), .QB (line364), .D(g4647), .CK(clk));
DFFX1 gate365(.Q (g926), .QB (line365), .D(g878), .CK(clk));
DFFX1 gate366(.Q (g368), .QB (line366), .D(g3838), .CK(clk));
DFFX1 gate367(.Q (g855), .QB (line367), .D(g8220), .CK(clk));
DFFX1 gate368(.Q (g1214), .QB (line368), .D(g5736), .CK(clk));
DFFX1 gate369(.Q (g1110), .QB (line369), .D(g7299), .CK(clk));
DFFX1 gate370(.Q (g1310), .QB (line370), .D(g1309), .CK(clk));
DFFX1 gate371(.Q (g296), .QB (line371), .D(g4617), .CK(clk));
DFFX1 gate372(.Q (g972), .QB (line372), .D(g2653), .CK(clk));
DFFX1 gate373(.Q (g1402), .QB (line373), .D(g6391), .CK(clk));
DFFX1 gate374(.Q (g1236), .QB (line374), .D(g1240), .CK(clk));
DFFX1 gate375(.Q (g896), .QB (line375), .D(g891), .CK(clk));
DFFX1 gate376(.Q (g613), .QB (line376), .D(g6820), .CK(clk));
DFFX1 gate377(.Q (g566), .QB (line377), .D(g3848), .CK(clk));
DFFX1 gate378(.Q (g1394), .QB (line378), .D(g6388), .CK(clk));
DFFX1 gate379(.Q (g1489), .QB (line379), .D(g7770), .CK(clk));
DFFX1 gate380(.Q (g883), .QB (line380), .D(g921), .CK(clk));
DFFX1 gate381(.Q (g47), .QB (line381), .D(g9389), .CK(clk));
DFFX1 gate382(.Q (g971), .QB (line382), .D(g5171), .CK(clk));
DFFX1 gate383(.Q (g609), .QB (line383), .D(g6808), .CK(clk));
DFFX1 gate384(.Q (g103), .QB (line384), .D(g5157), .CK(clk));
DFFX1 gate385(.Q (g1254), .QB (line385), .D(g6381), .CK(clk));
DFFX1 gate386(.Q (g556), .QB (line386), .D(g3847), .CK(clk));
DFFX1 gate387(.Q (g1409), .QB (line387), .D(g5178), .CK(clk));
DFFX1 gate388(.Q (g626), .QB (line388), .D(g6824), .CK(clk));
DFFX1 gate389(.Q (g1229), .QB (line389), .D(g7110), .CK(clk));
DFFX1 gate390(.Q (g782), .QB (line390), .D(g5734), .CK(clk));
DFFX1 gate391(.Q (g237), .QB (line391), .D(g6316), .CK(clk));
DFFX1 gate392(.Q (g942), .QB (line392), .D(g2652), .CK(clk));
DFFX1 gate393(.Q (g228), .QB (line393), .D(g6315), .CK(clk));
DFFX1 gate394(.Q (g706), .QB (line394), .D(g7750), .CK(clk));
DFFX1 gate395(.Q (g746), .QB (line395), .D(g8956), .CK(clk));
DFFX1 gate396(.Q (g1462), .QB (line396), .D(g8678), .CK(clk));
DFFX1 gate397(.Q (g963), .QB (line397), .D(g7764), .CK(clk));
DFFX1 gate398(.Q (g129), .QB (line398), .D(g5156), .CK(clk));
DFFX1 gate399(.Q (g837), .QB (line399), .D(g2649), .CK(clk));
DFFX1 gate400(.Q (g599), .QB (line400), .D(g6798), .CK(clk));
DFFX1 gate401(.Q (g1192), .QB (line401), .D(g1191), .CK(clk));
DFFX1 gate402(.Q (g828), .QB (line402), .D(g7762), .CK(clk));
DFFX1 gate403(.Q (g1392), .QB (line403), .D(g6387), .CK(clk));
DFFX1 gate404(.Q (g492), .QB (line404), .D(g6359), .CK(clk));
DFFX1 gate405(.Q (g95), .QB (line405), .D(g94), .CK(clk));
DFFX1 gate406(.Q (g944), .QB (line406), .D(g6372), .CK(clk));
DFFX1 gate407(.Q (g195), .QB (line407), .D(g3831), .CK(clk));
DFFX1 gate408(.Q (g1431), .QB (line408), .D(g2673), .CK(clk));
DFFX1 gate409(.Q (g1252), .QB (line409), .D(g2661), .CK(clk));
DFFX1 gate410(.Q (g356), .QB (line410), .D(g6335), .CK(clk));
DFFX1 gate411(.Q (g953), .QB (line411), .D(g8669), .CK(clk));
DFFX1 gate412(.Q (g1176), .QB (line412), .D(g5172), .CK(clk));
DFFX1 gate413(.Q (g1376), .QB (line413), .D(g6890), .CK(clk));
DFFX1 gate414(.Q (g1005), .QB (line414), .D(g1004), .CK(clk));
DFFX1 gate415(.Q (g1405), .QB (line415), .D(g5744), .CK(clk));
DFFX1 gate416(.Q (g901), .QB (line416), .D(g896), .CK(clk));
DFFX1 gate417(.Q (g1270), .QB (line417), .D(g1271), .CK(clk));
DFFX1 gate418(.Q (g1225), .QB (line418), .D(g6858), .CK(clk));
DFFX1 gate419(.Q (g1073), .QB (line419), .D(g9145), .CK(clk));
DFFX1 gate420(.Q (g1324), .QB (line420), .D(g7118), .CK(clk));
DFFX1 gate421(.Q (g1069), .QB (line421), .D(g9134), .CK(clk));
DFFX1 gate422(.Q (g443), .QB (line422), .D(g9101), .CK(clk));
DFFX1 gate423(.Q (g1377), .QB (line423), .D(g6891), .CK(clk));
DFFX1 gate424(.Q (g377), .QB (line424), .D(g4630), .CK(clk));
DFFX1 gate425(.Q (g618), .QB (line425), .D(g6816), .CK(clk));
DFFX1 gate426(.Q (g602), .QB (line426), .D(g6800), .CK(clk));
DFFX1 gate427(.Q (g213), .QB (line427), .D(g4602), .CK(clk));
DFFX1 gate428(.Q (g233), .QB (line428), .D(g4607), .CK(clk));
DFFX1 gate429(.Q (g1199), .QB (line429), .D(g6375), .CK(clk));
DFFX1 gate430(.Q (g1399), .QB (line430), .D(g3861), .CK(clk));
DFFX1 gate431(.Q (g83), .QB (line431), .D(g6779), .CK(clk));
DFFX1 gate432(.Q (g888), .QB (line432), .D(g7100), .CK(clk));
DFFX1 gate433(.Q (g573), .QB (line433), .D(g9033), .CK(clk));
DFFX1 gate434(.Q (g399), .QB (line434), .D(g6342), .CK(clk));
DFFX1 gate435(.Q (g1245), .QB (line435), .D(g1244), .CK(clk));
DFFX1 gate436(.Q (g507), .QB (line436), .D(g9114), .CK(clk));
DFFX1 gate437(.Q (g547), .QB (line437), .D(g9026), .CK(clk));
DFFX1 gate438(.Q (g108), .QB (line438), .D(g5147), .CK(clk));
DFFX1 gate439(.Q (g610), .QB (line439), .D(g6809), .CK(clk));
DFFX1 gate440(.Q (g630), .QB (line440), .D(g6828), .CK(clk));
DFFX1 gate441(.Q (g1207), .QB (line441), .D(g5173), .CK(clk));
DFFX1 gate442(.Q (g249), .QB (line442), .D(g6320), .CK(clk));
DFFX1 gate443(.Q (g65), .QB (line443), .D(g4598), .CK(clk));
DFFX1 gate444(.Q (g916), .QB (line444), .D(g911), .CK(clk));
DFFX1 gate445(.Q (g936), .QB (line445), .D(g5168), .CK(clk));
DFFX1 gate446(.Q (g478), .QB (line446), .D(g4648), .CK(clk));
DFFX1 gate447(.Q (g604), .QB (line447), .D(g6802), .CK(clk));
DFFX1 gate448(.Q (g945), .QB (line448), .D(g5170), .CK(clk));
DFFX1 gate449(.Q (g1114), .QB (line449), .D(g7521), .CK(clk));
DFFX1 gate450(.Q (g100), .QB (line450), .D(g99), .CK(clk));
DFFX1 gate451(.Q (g429), .QB (line451), .D(g9107), .CK(clk));
DFFX1 gate452(.Q (g809), .QB (line452), .D(g7511), .CK(clk));
DFFX1 gate453(.Q (g849), .QB (line453), .D(g2645), .CK(clk));
DFFX1 gate454(.Q (g1408), .QB (line454), .D(g5177), .CK(clk));
DFFX1 gate455(.Q (g1336), .QB (line455), .D(g6864), .CK(clk));
DFFX1 gate456(.Q (g601), .QB (line456), .D(g6799), .CK(clk));
DFFX1 gate457(.Q (g122), .QB (line457), .D(g6788), .CK(clk));
DFFX1 gate458(.Q (g1065), .QB (line458), .D(g9117), .CK(clk));
DFFX1 gate459(.Q (g1122), .QB (line459), .D(g8225), .CK(clk));
DFFX1 gate460(.Q (g1228), .QB (line460), .D(g7109), .CK(clk));
DFFX1 gate461(.Q (g495), .QB (line461), .D(g6360), .CK(clk));
DFFX1 gate462(.Q (g1322), .QB (line462), .D(g7116), .CK(clk));
DFFX1 gate463(.Q (g1230), .QB (line463), .D(g7300), .CK(clk));
DFFX1 gate464(.Q (g1033), .QB (line464), .D(g9034), .CK(clk));
DFFX1 gate465(.Q (g267), .QB (line465), .D(g9091), .CK(clk));
DFFX1 gate466(.Q (g1195), .QB (line466), .D(g6374), .CK(clk));
DFFX1 gate467(.Q (g1395), .QB (line467), .D(g1393), .CK(clk));
DFFX1 gate468(.Q (g373), .QB (line468), .D(g4626), .CK(clk));
DFFX1 gate469(.Q (g274), .QB (line469), .D(g4612), .CK(clk));
DFFX1 gate470(.Q (g1266), .QB (line470), .D(g5739), .CK(clk));
DFFX1 gate471(.Q (g714), .QB (line471), .D(g7752), .CK(clk));
DFFX1 gate472(.Q (g734), .QB (line472), .D(g7755), .CK(clk));
DFFX1 gate473(.Q (g1142), .QB (line473), .D(g8874), .CK(clk));
DFFX1 gate474(.Q (g1342), .QB (line474), .D(g7119), .CK(clk));
DFFX1 gate475(.Q (g769), .QB (line475), .D(g6843), .CK(clk));
DFFX1 gate476(.Q (g1081), .QB (line476), .D(g6852), .CK(clk));
DFFX1 gate477(.Q (g1481), .QB (line477), .D(g7769), .CK(clk));
DFFX1 gate478(.Q (g1097), .QB (line478), .D(g1185), .CK(clk));
DFFX1 gate479(.Q (g543), .QB (line479), .D(g3846), .CK(clk));
DFFX1 gate480(.Q (g1154), .QB (line480), .D(g1153), .CK(clk));
DFFX1 gate481(.Q (g1354), .QB (line481), .D(g7768), .CK(clk));
DFFX1 gate482(.Q (g489), .QB (line482), .D(g6358), .CK(clk));
DFFX1 gate483(.Q (g874), .QB (line483), .D(g4654), .CK(clk));
DFFX1 gate484(.Q (g121), .QB (line484), .D(g5154), .CK(clk));
DFFX1 gate485(.Q (g591), .QB (line485), .D(g9032), .CK(clk));
DFFX1 gate486(.Q (g616), .QB (line486), .D(g6814), .CK(clk));
DFFX1 gate487(.Q (g1267), .QB (line487), .D(g4656), .CK(clk));
DFFX1 gate488(.Q (g1312), .QB (line488), .D(g1311), .CK(clk));
DFFX1 gate489(.Q (g605), .QB (line489), .D(g6803), .CK(clk));
DFFX1 gate490(.Q (g182), .QB (line490), .D(g5161), .CK(clk));
DFFX1 gate491(.Q (g1401), .QB (line491), .D(g1399), .CK(clk));
DFFX1 gate492(.Q (g950), .QB (line492), .D(g8666), .CK(clk));
DFFX1 gate493(.Q (g1329), .QB (line493), .D(g2663), .CK(clk));
DFFX1 gate494(.Q (g408), .QB (line494), .D(g6345), .CK(clk));
DFFX1 gate495(.Q (g871), .QB (line495), .D(g5167), .CK(clk));
DFFX1 gate496(.Q (g759), .QB (line496), .D(g6832), .CK(clk));
DFFX1 gate497(.Q (g146), .QB (line497), .D(g7735), .CK(clk));
DFFX1 gate498(.Q (g202), .QB (line498), .D(g5732), .CK(clk));
DFFX1 gate499(.Q (g440), .QB (line499), .D(g6349), .CK(clk));
DFFX1 gate500(.Q (g476), .QB (line500), .D(g4646), .CK(clk));
DFFX1 gate501(.Q (g184), .QB (line501), .D(g6310), .CK(clk));
DFFX1 gate502(.Q (g1149), .QB (line502), .D(g7525), .CK(clk));
DFFX1 gate503(.Q (g1398), .QB (line503), .D(g1396), .CK(clk));
DFFX1 gate504(.Q (g210), .QB (line504), .D(g3834), .CK(clk));
DFFX1 gate505(.Q (g394), .QB (line505), .D(g4632), .CK(clk));
DFFX1 gate506(.Q (g86), .QB (line506), .D(g6780), .CK(clk));
DFFX1 gate507(.Q (g570), .QB (line507), .D(g9030), .CK(clk));
DFFX1 gate508(.Q (g275), .QB (line508), .D(g6322), .CK(clk));
DFFX1 gate509(.Q (g303), .QB (line509), .D(g6326), .CK(clk));
DFFX1 gate510(.Q (g125), .QB (line510), .D(g5155), .CK(clk));
DFFX1 gate511(.Q (g181), .QB (line511), .D(g5160), .CK(clk));
DFFX1 gate512(.Q (g1524), .QB (line512), .D(g6393), .CK(clk));
DFFX1 gate513(.Q (g595), .QB (line513), .D(g576), .CK(clk));
DFFX1 gate514(.Q (g1319), .QB (line514), .D(g7113), .CK(clk));
DFFX1 gate515(.Q (g863), .QB (line515), .D(g8222), .CK(clk));
DFFX1 gate516(.Q (g1211), .QB (line516), .D(g5174), .CK(clk));
DFFX1 gate517(.Q (g966), .QB (line517), .D(g8223), .CK(clk));
DFFX1 gate518(.Q (g1186), .QB (line518), .D(g1182), .CK(clk));
DFFX1 gate519(.Q (g1386), .QB (line519), .D(g6884), .CK(clk));
DFFX1 gate520(.Q (g875), .QB (line520), .D(g5165), .CK(clk));
DFFX1 gate521(.Q (g1170), .QB (line521), .D(g1173), .CK(clk));
DFFX1 gate522(.Q (g1370), .QB (line522), .D(g6876), .CK(clk));
DFFX1 gate523(.Q (g201), .QB (line523), .D(g200), .CK(clk));
DFFX1 gate524(.Q (g1325), .QB (line524), .D(g7305), .CK(clk));
DFFX1 gate525(.Q (g1280), .QB (line525), .D(g7112), .CK(clk));
DFFX1 gate526(.Q (g1106), .QB (line526), .D(g7107), .CK(clk));
DFFX1 gate527(.Q (g1061), .QB (line527), .D(g9035), .CK(clk));
DFFX1 gate528(.Q (g1387), .QB (line528), .D(g6885), .CK(clk));
DFFX1 gate529(.Q (g762), .QB (line529), .D(g6835), .CK(clk));
DFFX1 gate530(.Q (g1461), .QB (line530), .D(g4669), .CK(clk));
DFFX1 gate531(.Q (g378), .QB (line531), .D(g6337), .CK(clk));
DFFX1 gate532(.Q (g1200), .QB (line532), .D(g1199), .CK(clk));
DFFX1 gate533(.Q (g1514), .QB (line533), .D(g7775), .CK(clk));
DFFX1 gate534(.Q (g1403), .QB (line534), .D(g1402), .CK(clk));
DFFX1 gate535(.Q (g1345), .QB (line535), .D(g7528), .CK(clk));
DFFX1 gate536(.Q (g1191), .QB (line536), .D(g6373), .CK(clk));
DFFX1 gate537(.Q (g1391), .QB (line537), .D(g1390), .CK(clk));
DFFX1 gate538(.Q (g185), .QB (line538), .D(g4599), .CK(clk));
DFFX1 gate539(.Q (g1307), .QB (line539), .D(g3858), .CK(clk));
DFFX1 gate540(.Q (g1159), .QB (line540), .D(g1157), .CK(clk));
DFFX1 gate541(.Q (g1223), .QB (line541), .D(g6379), .CK(clk));
DFFX1 gate542(.Q (g446), .QB (line542), .D(g9102), .CK(clk));
DFFX1 gate543(.Q (g1416), .QB (line543), .D(g4665), .CK(clk));
DFFX1 gate544(.Q (g395), .QB (line544), .D(g4633), .CK(clk));
DFFX1 gate545(.Q (g764), .QB (line545), .D(g6837), .CK(clk));
DFFX1 gate546(.Q (g1251), .QB (line546), .D(g6860), .CK(clk));
DFFX1 gate547(.Q (g216), .QB (line547), .D(g6311), .CK(clk));
DFFX1 gate548(.Q (g236), .QB (line548), .D(g4610), .CK(clk));
DFFX1 gate549(.Q (g205), .QB (line549), .D(g3835), .CK(clk));
DFFX1 gate550(.Q (g540), .QB (line550), .D(g6364), .CK(clk));
DFFX1 gate551(.Q (g576), .QB (line551), .D(g3849), .CK(clk));
DFFX1 gate552(.Q (g1537), .QB (line552), .D(g7777), .CK(clk));
DFFX1 gate553(.Q (g727), .QB (line553), .D(g8228), .CK(clk));
DFFX1 gate554(.Q (g999), .QB (line554), .D(g8865), .CK(clk));
DFFX1 gate555(.Q (g761), .QB (line555), .D(g6834), .CK(clk));
DFFX1 gate556(.Q (g1272), .QB (line556), .D(g6383), .CK(clk));
DFFX1 gate557(.Q (g1243), .QB (line557), .D(g2660), .CK(clk));
DFFX1 gate558(.Q (g1328), .QB (line558), .D(g7309), .CK(clk));
DFFX1 gate559(.Q (g1130), .QB (line559), .D(g7522), .CK(clk));
DFFX1 gate560(.Q (g1330), .QB (line560), .D(g6862), .CK(clk));
DFFX1 gate561(.Q (g114), .QB (line561), .D(g6786), .CK(clk));
DFFX1 gate562(.Q (g134), .QB (line562), .D(g6791), .CK(clk));
DFFX1 gate563(.Q (g1166), .QB (line563), .D(g1167), .CK(clk));
DFFX1 gate564(.Q (g524), .QB (line564), .D(g9109), .CK(clk));
DFFX1 gate565(.Q (g1366), .QB (line565), .D(g6866), .CK(clk));
DFFX1 gate566(.Q (g348), .QB (line566), .D(g9099), .CK(clk));
DFFX1 gate567(.Q (g1148), .QB (line567), .D(g1147), .CK(clk));
DFFX1 gate568(.Q (g1348), .QB (line568), .D(g7529), .CK(clk));
DFFX1 gate569(.Q (g1155), .QB (line569), .D(g1154), .CK(clk));
DFFX1 gate570(.Q (g1260), .QB (line570), .D(g6382), .CK(clk));
DFFX1 gate571(.Q (g7), .QB (line571), .D(g9375), .CK(clk));
DFFX1 gate572(.Q (g258), .QB (line572), .D(g9088), .CK(clk));
DFFX1 gate573(.Q (g521), .QB (line573), .D(g6362), .CK(clk));
DFFX1 gate574(.Q (g300), .QB (line574), .D(g6325), .CK(clk));
DFFX1 gate575(.Q (g765), .QB (line575), .D(g6838), .CK(clk));
DFFX1 gate576(.Q (g1118), .QB (line576), .D(g7766), .CK(clk));
DFFX1 gate577(.Q (g1167), .QB (line577), .D(g1170), .CK(clk));
DFFX1 gate578(.Q (g1318), .QB (line578), .D(g6861), .CK(clk));
DFFX1 gate579(.Q (g1367), .QB (line579), .D(g6873), .CK(clk));
DFFX1 gate580(.Q (g677), .QB (line580), .D(g7747), .CK(clk));
DFFX1 gate581(.Q (g376), .QB (line581), .D(g4629), .CK(clk));
DFFX1 gate582(.Q (g1057), .QB (line582), .D(g8959), .CK(clk));
DFFX1 gate583(.Q (g973), .QB (line583), .D(g8672), .CK(clk));
DFFX1 gate584(.Q (g1193), .QB (line584), .D(g1192), .CK(clk));
DFFX1 gate585(.Q (g1393), .QB (line585), .D(g2664), .CK(clk));
DFFX1 gate586(.Q (g1549), .QB (line586), .D(g7780), .CK(clk));
DFFX1 gate587(.Q (g1321), .QB (line587), .D(g7115), .CK(clk));
DFFX1 gate588(.Q (g1253), .QB (line588), .D(g5741), .CK(clk));
DFFX1 gate589(.Q (g1519), .QB (line589), .D(g8227), .CK(clk));
DFFX1 gate590(.Q (g584), .QB (line590), .D(g6369), .CK(clk));
DFFX1 gate591(.Q (g539), .QB (line591), .D(g3845), .CK(clk));
DFFX1 gate592(.Q (g324), .QB (line592), .D(g6331), .CK(clk));
DFFX1 gate593(.Q (g432), .QB (line593), .D(g9108), .CK(clk));
DFFX1 gate594(.Q (g1158), .QB (line594), .D(g1159), .CK(clk));
DFFX1 gate595(.Q (g321), .QB (line595), .D(g6330), .CK(clk));
DFFX1 gate596(.Q (g1311), .QB (line596), .D(g1310), .CK(clk));
DFFX1 gate597(.Q (g414), .QB (line597), .D(g6347), .CK(clk));
DFFX1 gate598(.Q (g1374), .QB (line598), .D(g6872), .CK(clk));
DFFX1 gate599(.Q (g94), .QB (line599), .D(g6782), .CK(clk));
DFFX1 gate600(.Q (g1284), .QB (line600), .D(g7301), .CK(clk));
DFFX1 gate601(.Q (g1545), .QB (line601), .D(g7779), .CK(clk));
DFFX1 gate602(.Q (g1380), .QB (line602), .D(g6886), .CK(clk));
DFFX1 gate603(.Q (g673), .QB (line603), .D(g7746), .CK(clk));
DFFX1 gate604(.Q (g607), .QB (line604), .D(g6805), .CK(clk));
DFFX1 gate605(.Q (g306), .QB (line605), .D(g6327), .CK(clk));
DFFX1 gate606(.Q (g943), .QB (line606), .D(g8671), .CK(clk));
DFFX1 gate607(.Q (g162), .QB (line607), .D(g7741), .CK(clk));
DFFX1 gate608(.Q (g411), .QB (line608), .D(g6346), .CK(clk));
DFFX1 gate609(.Q (g866), .QB (line609), .D(g5163), .CK(clk));
DFFX1 gate610(.Q (g1204), .QB (line610), .D(g1203), .CK(clk));
DFFX1 gate611(.Q (g1300), .QB (line611), .D(g7303), .CK(clk));
DFFX1 gate612(.Q (g384), .QB (line612), .D(g6339), .CK(clk));
DFFX1 gate613(.Q (g339), .QB (line613), .D(g9096), .CK(clk));
DFFX1 gate614(.Q (g459), .QB (line614), .D(g6350), .CK(clk));
DFFX1 gate615(.Q (g1323), .QB (line615), .D(g7117), .CK(clk));
DFFX1 gate616(.Q (g381), .QB (line616), .D(g6338), .CK(clk));
DFFX1 gate617(.Q (g1528), .QB (line617), .D(g7776), .CK(clk));
DFFX1 gate618(.Q (g1351), .QB (line618), .D(g7530), .CK(clk));
DFFX1 gate619(.Q (g597), .QB (line619), .D(g6796), .CK(clk));
DFFX1 gate620(.Q (g1372), .QB (line620), .D(g6870), .CK(clk));
DFFX1 gate621(.Q (g154), .QB (line621), .D(g7739), .CK(clk));
DFFX1 gate622(.Q (g435), .QB (line622), .D(g4637), .CK(clk));
DFFX1 gate623(.Q (g970), .QB (line623), .D(g963), .CK(clk));
DFFX1 gate624(.Q (g1134), .QB (line624), .D(g7523), .CK(clk));
DFFX1 gate625(.Q (g995), .QB (line625), .D(g7517), .CK(clk));
DFFX1 gate626(.Q (g190), .QB (line626), .D(g201), .CK(clk));
DFFX1 gate627(.Q (g1313), .QB (line627), .D(g5742), .CK(clk));
DFFX1 gate628(.Q (g603), .QB (line628), .D(g6801), .CK(clk));
DFFX1 gate629(.Q (g1494), .QB (line629), .D(g7771), .CK(clk));
DFFX1 gate630(.Q (g462), .QB (line630), .D(g6351), .CK(clk));
DFFX1 gate631(.Q (g1160), .QB (line631), .D(g1163), .CK(clk));
DFFX1 gate632(.Q (g1360), .QB (line632), .D(g8676), .CK(clk));
DFFX1 gate633(.Q (g1450), .QB (line633), .D(g5186), .CK(clk));
DFFX1 gate634(.Q (g187), .QB (line634), .D(g5730), .CK(clk));
DFFX1 gate635(.Q (g1179), .QB (line635), .D(g1186), .CK(clk));
DFFX1 gate636(.Q (g1379), .QB (line636), .D(g6879), .CK(clk));
DFFX1 gate637(.Q (g12), .QB (line637), .D(g8662), .CK(clk));
DFFX1 gate638(.Q (g71), .QB (line638), .D(g6775), .CK(clk));
INVX1 gate639(.O (g1658), .I (g1313));
INVX1 gate640(.O (g1777), .I (g611));
INVX1 gate641(.O (I9325), .I (g4242));
INVX1 gate642(.O (I7758), .I (g2605));
INVX1 gate643(.O (g5652), .I (I10135));
INVX1 gate644(.O (I13502), .I (g7135));
INVX1 gate645(.O (g6895), .I (I12558));
INVX1 gate646(.O (g3880), .I (g2965));
INVX1 gate647(.O (g6837), .I (I12382));
INVX1 gate648(.O (I15824), .I (g9157));
INVX1 gate649(.O (g5843), .I (g5367));
INVX1 gate650(.O (I6112), .I (g4));
INVX1 gate651(.O (g7189), .I (I13109));
INVX1 gate652(.O (g8970), .I (I15414));
INVX1 gate653(.O (I6267), .I (g100));
INVX1 gate654(.O (g6062), .I (I10675));
INVX1 gate655(.O (I16126), .I (g9354));
INVX1 gate656(.O (I10519), .I (g5242));
INVX1 gate657(.O (I15181), .I (g8734));
INVX1 gate658(.O (I11443), .I (g6038));
INVX1 gate659(.O (I12436), .I (g6635));
INVX1 gate660(.O (I10675), .I (g5662));
INVX1 gate661(.O (g2547), .I (I6371));
INVX1 gate662(.O (I7365), .I (g3061));
INVX1 gate663(.O (I10154), .I (g5109));
INVX1 gate664(.O (g1611), .I (g1073));
INVX1 gate665(.O (I11278), .I (g5780));
INVX1 gate666(.O (g7171), .I (g7071));
INVX1 gate667(.O (I14154), .I (g7558));
INVX1 gate668(.O (I12274), .I (g6672));
INVX1 gate669(.O (g8224), .I (I14451));
INVX1 gate670(.O (g5834), .I (I10525));
INVX1 gate671(.O (g5971), .I (I10587));
INVX1 gate672(.O (g3978), .I (g3160));
INVX1 gate673(.O (I6676), .I (g1603));
INVX1 gate674(.O (g3612), .I (I7082));
INVX1 gate675(.O (I8520), .I (g3652));
INVX1 gate676(.O (g2892), .I (g2266));
INVX1 gate677(.O (I13469), .I (g7123));
INVX1 gate678(.O (I12346), .I (g6737));
INVX1 gate679(.O (I9636), .I (g4802));
INVX1 gate680(.O (I14637), .I (g8012));
INVX1 gate681(.O (g6788), .I (I12235));
INVX1 gate682(.O (g1799), .I (I5657));
INVX1 gate683(.O (g3935), .I (I7602));
INVX1 gate684(.O (I5933), .I (g1158));
INVX1 gate685(.O (g9207), .I (g9197));
INVX1 gate686(.O (I13039), .I (g6961));
INVX1 gate687(.O (I15426), .I (g8895));
INVX1 gate688(.O (g5598), .I (g4938));
INVX1 gate689(.O (g1674), .I (g1514));
INVX1 gate690(.O (g7281), .I (I13277));
INVX1 gate691(.O (g3982), .I (g3192));
INVX1 gate692(.O (g4666), .I (I8913));
INVX1 gate693(.O (I15190), .I (g8685));
INVX1 gate694(.O (g2945), .I (g2364));
INVX1 gate695(.O (g5121), .I (I9515));
INVX1 gate696(.O (g3128), .I (I6839));
INVX1 gate697(.O (g3629), .I (g2424));
INVX1 gate698(.O (g7297), .I (I13323));
INVX1 gate699(.O (g5670), .I (I10157));
INVX1 gate700(.O (I11815), .I (g6169));
INVX1 gate701(.O (g6842), .I (I12397));
INVX1 gate702(.O (g3130), .I (I6849));
INVX1 gate703(.O (g9088), .I (I15654));
INVX1 gate704(.O (g8789), .I (g8564));
INVX1 gate705(.O (g3542), .I (g1777));
INVX1 gate706(.O (I12292), .I (g6657));
INVX1 gate707(.O (g6298), .I (I11221));
INVX1 gate708(.O (g2709), .I (g1747));
INVX1 gate709(.O (I11677), .I (g6076));
INVX1 gate710(.O (g6392), .I (I11503));
INVX1 gate711(.O (g4648), .I (I8859));
INVX1 gate712(.O (I8829), .I (g4029));
INVX1 gate713(.O (I15546), .I (g9007));
INVX1 gate714(.O (g1680), .I (I5515));
INVX1 gate715(.O (I15211), .I (g8808));
INVX1 gate716(.O (g2340), .I (g1327));
INVX1 gate717(.O (I12409), .I (g6398));
INVX1 gate718(.O (g4655), .I (I8880));
INVX1 gate719(.O (g7745), .I (I14106));
INVX1 gate720(.O (g7138), .I (I12996));
INVX1 gate721(.O (I6703), .I (g1983));
INVX1 gate722(.O (g5938), .I (g5412));
INVX1 gate723(.O (g8771), .I (g8564));
INVX1 gate724(.O (g2478), .I (g31));
INVX1 gate725(.O (g5813), .I (I10472));
INVX1 gate726(.O (g7338), .I (I13432));
INVX1 gate727(.O (g2907), .I (g2289));
INVX1 gate728(.O (g1744), .I (g600));
INVX1 gate729(.O (g9215), .I (I15921));
INVX1 gate730(.O (g7109), .I (I12915));
INVX1 gate731(.O (g6854), .I (I12433));
INVX1 gate732(.O (I12635), .I (g6509));
INVX1 gate733(.O (g7309), .I (I13359));
INVX1 gate734(.O (g1802), .I (g628));
INVX1 gate735(.O (I10439), .I (g5214));
INVX1 gate736(.O (g2959), .I (g1926));
INVX1 gate737(.O (I14728), .I (g8152));
INVX1 gate738(.O (I8733), .I (g3996));
INVX1 gate739(.O (I14439), .I (g8063));
INVX1 gate740(.O (g2517), .I (I6348));
INVX1 gate741(.O (g4010), .I (g3097));
INVX1 gate742(.O (I7662), .I (g3642));
INVX1 gate743(.O (I9446), .I (g3926));
INVX1 gate744(.O (I8974), .I (g3871));
INVX1 gate745(.O (g5740), .I (I10277));
INVX1 gate746(.O (g5519), .I (I9929));
INVX1 gate747(.O (g9114), .I (I15732));
INVX1 gate748(.O (g1558), .I (I5435));
INVX1 gate749(.O (I7290), .I (g2936));
INVX1 gate750(.O (g2876), .I (g2231));
INVX1 gate751(.O (g9314), .I (I16058));
INVX1 gate752(.O (I11884), .I (g6091));
INVX1 gate753(.O (I9145), .I (g4264));
INVX1 gate754(.O (I6468), .I (g1917));
INVX1 gate755(.O (g5606), .I (g4748));
INVX1 gate756(.O (I8796), .I (g3934));
INVX1 gate757(.O (g7759), .I (I14148));
INVX1 gate758(.O (I14349), .I (g7588));
INVX1 gate759(.O (I11410), .I (g5845));
INVX1 gate760(.O (I12164), .I (g5847));
INVX1 gate761(.O (g695), .I (I5392));
INVX1 gate762(.O (g6708), .I (g6250));
INVX1 gate763(.O (I13410), .I (g7274));
INVX1 gate764(.O (I15625), .I (g9000));
INVX1 gate765(.O (g6520), .I (I11704));
INVX1 gate766(.O (g1901), .I (I5781));
INVX1 gate767(.O (g6219), .I (I10998));
INVX1 gate768(.O (g6640), .I (I11908));
INVX1 gate769(.O (I8980), .I (g4535));
INVX1 gate770(.O (g3902), .I (I7495));
INVX1 gate771(.O (I12891), .I (g6950));
INVX1 gate772(.O (I11479), .I (g6201));
INVX1 gate773(.O (I11666), .I (g5772));
INVX1 gate774(.O (g5687), .I (I10190));
INVX1 gate775(.O (g2915), .I (I6643));
INVX1 gate776(.O (I13666), .I (g7238));
INVX1 gate777(.O (g6252), .I (g5418));
INVX1 gate778(.O (g6812), .I (I12307));
INVX1 gate779(.O (g4372), .I (I8357));
INVX1 gate780(.O (g7049), .I (I12813));
INVX1 gate781(.O (g3512), .I (g1616));
INVX1 gate782(.O (I13478), .I (g7126));
INVX1 gate783(.O (g5586), .I (g4938));
INVX1 gate784(.O (g6958), .I (I12675));
INVX1 gate785(.O (I15943), .I (g9214));
INVX1 gate786(.O (g4618), .I (I8769));
INVX1 gate787(.O (I6716), .I (g1721));
INVX1 gate788(.O (g6376), .I (I11455));
INVX1 gate789(.O (g4667), .I (I8916));
INVX1 gate790(.O (I5981), .I (g459));
INVX1 gate791(.O (I8177), .I (g2810));
INVX1 gate792(.O (I7847), .I (g3798));
INVX1 gate793(.O (I16055), .I (g9291));
INVX1 gate794(.O (g9336), .I (I16084));
INVX1 gate795(.O (g2310), .I (I6087));
INVX1 gate796(.O (g7715), .I (I14022));
INVX1 gate797(.O (g1600), .I (g976));
INVX1 gate798(.O (g1574), .I (g681));
INVX1 gate799(.O (g1864), .I (g162));
INVX1 gate800(.O (g4566), .I (g2902));
INVX1 gate801(.O (I11556), .I (g6065));
INVX1 gate802(.O (g7098), .I (g6525));
INVX1 gate803(.O (I5997), .I (g114));
INVX1 gate804(.O (g6829), .I (I12358));
INVX1 gate805(.O (g7498), .I (I13672));
INVX1 gate806(.O (g2663), .I (I6460));
INVX1 gate807(.O (I12108), .I (g5939));
INVX1 gate808(.O (g6765), .I (I12164));
INVX1 gate809(.O (g3529), .I (g2323));
INVX1 gate810(.O (g8959), .I (I15391));
INVX1 gate811(.O (I6198), .I (g483));
INVX1 gate812(.O (g4693), .I (I8974));
INVX1 gate813(.O (I13580), .I (g7208));
INVX1 gate814(.O (g4134), .I (g3676));
INVX1 gate815(.O (g3649), .I (g2424));
INVX1 gate816(.O (I14139), .I (g7548));
INVX1 gate817(.O (I9416), .I (g4273));
INVX1 gate818(.O (I12283), .I (g6692));
INVX1 gate819(.O (g8482), .I (g8094));
INVX1 gate820(.O (g5525), .I (g4934));
INVX1 gate821(.O (g3851), .I (I7356));
INVX1 gate822(.O (g5645), .I (g4748));
INVX1 gate823(.O (I5353), .I (g3833));
INVX1 gate824(.O (g2402), .I (g29));
INVX1 gate825(.O (I7950), .I (g2774));
INVX1 gate826(.O (g2824), .I (g1688));
INVX1 gate827(.O (g1580), .I (g706));
INVX1 gate828(.O (g2236), .I (I5969));
INVX1 gate829(.O (g7584), .I (I13897));
INVX1 gate830(.O (g4555), .I (g2894));
INVX1 gate831(.O (g9065), .I (I15589));
INVX1 gate832(.O (I9642), .I (g4788));
INVX1 gate833(.O (g7539), .I (I13797));
INVX1 gate834(.O (I15411), .I (g8897));
INVX1 gate835(.O (I15527), .I (g9020));
INVX1 gate836(.O (I10415), .I (g5397));
INVX1 gate837(.O (I13084), .I (g7071));
INVX1 gate838(.O (g9322), .I (g9313));
INVX1 gate839(.O (g3964), .I (g3160));
INVX1 gate840(.O (g4792), .I (I9111));
INVX1 gate841(.O (g9230), .I (I15950));
INVX1 gate842(.O (g6225), .I (I11014));
INVX1 gate843(.O (I8781), .I (g3932));
INVX1 gate844(.O (I8898), .I (g4089));
INVX1 gate845(.O (g6073), .I (g5384));
INVX1 gate846(.O (g2877), .I (g2232));
INVX1 gate847(.O (g6796), .I (I12259));
INVX1 gate848(.O (g1736), .I (I5577));
INVX1 gate849(.O (I12091), .I (g5988));
INVX1 gate850(.O (g4621), .I (I8778));
INVX1 gate851(.O (g5607), .I (g4938));
INVX1 gate852(.O (g9033), .I (I15513));
INVX1 gate853(.O (g7162), .I (I13060));
INVX1 gate854(.O (g7268), .I (I13244));
INVX1 gate855(.O (g7019), .I (I12771));
INVX1 gate856(.O (I11740), .I (g6136));
INVX1 gate857(.O (g7362), .I (I13502));
INVX1 gate858(.O (g5158), .I (I9600));
INVX1 gate859(.O (I13740), .I (g7364));
INVX1 gate860(.O (I9654), .I (g4792));
INVX1 gate861(.O (I15894), .I (g9195));
INVX1 gate862(.O (g6324), .I (I11299));
INVX1 gate863(.O (I7723), .I (g3052));
INVX1 gate864(.O (g4113), .I (I7950));
INVX1 gate865(.O (g6069), .I (I10690));
INVX1 gate866(.O (g2556), .I (g1190));
INVX1 gate867(.O (g1889), .I (g1018));
INVX1 gate868(.O (I7101), .I (g2478));
INVX1 gate869(.O (I5901), .I (g52));
INVX1 gate870(.O (g2222), .I (I5939));
INVX1 gate871(.O (I13676), .I (g7256));
INVX1 gate872(.O (g9096), .I (I15678));
INVX1 gate873(.O (I8291), .I (g878));
INVX1 gate874(.O (I13373), .I (g7270));
INVX1 gate875(.O (g2928), .I (g2326));
INVX1 gate876(.O (g4202), .I (g2810));
INVX1 gate877(.O (g8663), .I (I14783));
INVX1 gate878(.O (I7605), .I (g2752));
INVX1 gate879(.O (I15714), .I (g9077));
INVX1 gate880(.O (g5587), .I (g4938));
INVX1 gate881(.O (g2930), .I (g2328));
INVX1 gate882(.O (I15315), .I (g8738));
INVX1 gate883(.O (I11800), .I (g6164));
INVX1 gate884(.O (g1871), .I (I5754));
INVX1 gate885(.O (g4908), .I (g4088));
INVX1 gate886(.O (g6377), .I (I11458));
INVX1 gate887(.O (g6206), .I (g5639));
INVX1 gate888(.O (g5311), .I (g4938));
INVX1 gate889(.O (g2899), .I (g2272));
INVX1 gate890(.O (g9195), .I (I15871));
INVX1 gate891(.O (g4094), .I (I7905));
INVX1 gate892(.O (I11936), .I (g5918));
INVX1 gate893(.O (g3872), .I (g2954));
INVX1 gate894(.O (I15202), .I (g8797));
INVX1 gate895(.O (g3652), .I (I7132));
INVX1 gate896(.O (g4567), .I (g2903));
INVX1 gate897(.O (g7728), .I (I14055));
INVX1 gate898(.O (g7486), .I (I13646));
INVX1 gate899(.O (g3843), .I (I7332));
INVX1 gate900(.O (g3989), .I (g3131));
INVX1 gate901(.O (I6186), .I (g138));
INVX1 gate902(.O (g7730), .I (I14061));
INVX1 gate903(.O (I9612), .I (g4776));
INVX1 gate904(.O (I10608), .I (g5701));
INVX1 gate905(.O (g5174), .I (I9648));
INVX1 gate906(.O (g8762), .I (g8585));
INVX1 gate907(.O (g7504), .I (I13692));
INVX1 gate908(.O (I15978), .I (g9235));
INVX1 gate909(.O (I14115), .I (g7563));
INVX1 gate910(.O (g7185), .I (I13099));
INVX1 gate911(.O (g4776), .I (I9081));
INVX1 gate912(.O (I7041), .I (g2401));
INVX1 gate913(.O (g6849), .I (I12418));
INVX1 gate914(.O (I9935), .I (g4812));
INVX1 gate915(.O (g4593), .I (g2939));
INVX1 gate916(.O (I11964), .I (g5971));
INVX1 gate917(.O (g3549), .I (g2404));
INVX1 gate918(.O (g3834), .I (I7305));
INVX1 gate919(.O (g3971), .I (I7688));
INVX1 gate920(.O (g7070), .I (g6562));
INVX1 gate921(.O (g2295), .I (g995));
INVX1 gate922(.O (I14052), .I (g7494));
INVX1 gate923(.O (g2237), .I (I5972));
INVX1 gate924(.O (g7470), .I (g7253));
INVX1 gate925(.O (I15741), .I (g9083));
INVX1 gate926(.O (g8657), .I (I14763));
INVX1 gate927(.O (g6781), .I (I12214));
INVX1 gate928(.O (g7425), .I (I13550));
INVX1 gate929(.O (g5180), .I (I9666));
INVX1 gate930(.O (g2844), .I (I6574));
INVX1 gate931(.O (I8215), .I (g3577));
INVX1 gate932(.O (g6898), .I (I12567));
INVX1 gate933(.O (g1838), .I (g1450));
INVX1 gate934(.O (g5591), .I (g4841));
INVX1 gate935(.O (g6900), .I (I12571));
INVX1 gate936(.O (g8222), .I (I14445));
INVX1 gate937(.O (I8886), .I (g4308));
INVX1 gate938(.O (g5832), .I (I10519));
INVX1 gate939(.O (I14813), .I (g8640));
INVX1 gate940(.O (g1795), .I (I5649));
INVX1 gate941(.O (g6797), .I (I12262));
INVX1 gate942(.O (g1737), .I (g597));
INVX1 gate943(.O (g2394), .I (I6270));
INVX1 gate944(.O (g9248), .I (I15978));
INVX1 gate945(.O (g1809), .I (g759));
INVX1 gate946(.O (I10973), .I (g5726));
INVX1 gate947(.O (I14798), .I (g8605));
INVX1 gate948(.O (g6245), .I (g5690));
INVX1 gate949(.O (g4360), .I (I8333));
INVX1 gate950(.O (I7368), .I (g3018));
INVX1 gate951(.O (g9255), .I (I15985));
INVX1 gate952(.O (g9081), .I (I15635));
INVX1 gate953(.O (I12948), .I (g6919));
INVX1 gate954(.O (I13909), .I (g7339));
INVX1 gate955(.O (I15735), .I (g9078));
INVX1 gate956(.O (g4521), .I (g2866));
INVX1 gate957(.O (I14184), .I (g7726));
INVX1 gate958(.O (g1672), .I (g1499));
INVX1 gate959(.O (I14674), .I (g7788));
INVX1 gate960(.O (g8464), .I (g8039));
INVX1 gate961(.O (g6291), .I (I11200));
INVX1 gate962(.O (I12702), .I (g6497));
INVX1 gate963(.O (g2557), .I (g940));
INVX1 gate964(.O (g4050), .I (g3080));
INVX1 gate965(.O (g4641), .I (I8838));
INVX1 gate966(.O (I11908), .I (g5918));
INVX1 gate967(.O (I12757), .I (g6577));
INVX1 gate968(.O (g9097), .I (I15681));
INVX1 gate969(.O (g2966), .I (g1856));
INVX1 gate970(.O (g5794), .I (I10421));
INVX1 gate971(.O (I5889), .I (g83));
INVX1 gate972(.O (g1643), .I (g1211));
INVX1 gate973(.O (I11569), .I (g6279));
INVX1 gate974(.O (g7131), .I (g6976));
INVX1 gate975(.O (g6344), .I (I11359));
INVX1 gate976(.O (g2471), .I (I6309));
INVX1 gate977(.O (g7006), .I (I12748));
INVX1 gate978(.O (g7331), .I (I13413));
INVX1 gate979(.O (I15196), .I (g8778));
INVX1 gate980(.O (I6636), .I (g1704));
INVX1 gate981(.O (I14732), .I (g8155));
INVX1 gate982(.O (g2242), .I (g985));
INVX1 gate983(.O (g6207), .I (I10962));
INVX1 gate984(.O (g3909), .I (I7520));
INVX1 gate985(.O (I11747), .I (g6123));
INVX1 gate986(.O (I12564), .I (g6720));
INVX1 gate987(.O (g8563), .I (I14662));
INVX1 gate988(.O (g2948), .I (g2366));
INVX1 gate989(.O (I11242), .I (g6183));
INVX1 gate990(.O (g7766), .I (I14169));
INVX1 gate991(.O (g6819), .I (I12328));
INVX1 gate992(.O (g7105), .I (I12903));
INVX1 gate993(.O (g3519), .I (g2185));
INVX1 gate994(.O (I10761), .I (g5302));
INVX1 gate995(.O (g7305), .I (I13347));
INVX1 gate996(.O (I7856), .I (g3805));
INVX1 gate997(.O (I7734), .I (g2595));
INVX1 gate998(.O (g2955), .I (I6703));
INVX1 gate999(.O (g7487), .I (I13649));
INVX1 gate1000(.O (g5628), .I (g4748));
INVX1 gate1001(.O (g1742), .I (g1486));
INVX1 gate1002(.O (g6088), .I (I10708));
INVX1 gate1003(.O (g6852), .I (I12427));
INVX1 gate1004(.O (g5515), .I (g4923));
INVX1 gate1005(.O (I12397), .I (g6764));
INVX1 gate1006(.O (g6488), .I (I11652));
INVX1 gate1007(.O (g4658), .I (I8889));
INVX1 gate1008(.O (g7748), .I (I14115));
INVX1 gate1009(.O (g4777), .I (I9084));
INVX1 gate1010(.O (I10400), .I (g5201));
INVX1 gate1011(.O (g5100), .I (I9484));
INVX1 gate1012(.O (I9512), .I (g3985));
INVX1 gate1013(.O (I13807), .I (g7320));
INVX1 gate1014(.O (I11974), .I (g5956));
INVX1 gate1015(.O (I12062), .I (g5988));
INVX1 gate1016(.O (I14400), .I (g7677));
INVX1 gate1017(.O (g2350), .I (I6166));
INVX1 gate1018(.O (g9112), .I (I15726));
INVX1 gate1019(.O (g7755), .I (I14136));
INVX1 gate1020(.O (g9218), .I (I15930));
INVX1 gate1021(.O (g1926), .I (g874));
INVX1 gate1022(.O (I9823), .I (g5138));
INVX1 gate1023(.O (g9312), .I (I16052));
INVX1 gate1024(.O (g2038), .I (g809));
INVX1 gate1025(.O (g4882), .I (g4069));
INVX1 gate1026(.O (I14214), .I (g7576));
INVX1 gate1027(.O (I12933), .I (g7018));
INVX1 gate1028(.O (I9366), .I (g4350));
INVX1 gate1029(.O (g7226), .I (g6937));
INVX1 gate1030(.O (I11230), .I (g6140));
INVX1 gate1031(.O (I11293), .I (g5824));
INVX1 gate1032(.O (I10207), .I (g5075));
INVX1 gate1033(.O (I13293), .I (g7159));
INVX1 gate1034(.O (I12508), .I (g6593));
INVX1 gate1035(.O (I11638), .I (g5847));
INVX1 gate1036(.O (g6886), .I (I12529));
INVX1 gate1037(.O (I6446), .I (g1812));
INVX1 gate1038(.O (g4611), .I (I8748));
INVX1 gate1039(.O (g291), .I (I5356));
INVX1 gate1040(.O (I14005), .I (g7434));
INVX1 gate1041(.O (g7045), .I (g6490));
INVX1 gate1042(.O (I11416), .I (g5829));
INVX1 gate1043(.O (I10538), .I (g5255));
INVX1 gate1044(.O (I6003), .I (g228));
INVX1 gate1045(.O (I9148), .I (g4354));
INVX1 gate1046(.O (I13416), .I (g7165));
INVX1 gate1047(.O (I5795), .I (g1236));
INVX1 gate1048(.O (g9129), .I (I15765));
INVX1 gate1049(.O (g2769), .I (g2424));
INVX1 gate1050(.O (g7173), .I (g6980));
INVX1 gate1051(.O (g9329), .I (g9317));
INVX1 gate1052(.O (g6314), .I (I11269));
INVX1 gate1053(.O (g7091), .I (g6525));
INVX1 gate1054(.O (g7491), .I (I13653));
INVX1 gate1055(.O (g6870), .I (I12481));
INVX1 gate1056(.O (g3860), .I (I7383));
INVX1 gate1057(.O (g2918), .I (g2310));
INVX1 gate1058(.O (g3341), .I (I6936));
INVX1 gate1059(.O (g1983), .I (I5839));
INVX1 gate1060(.O (g6825), .I (I12346));
INVX1 gate1061(.O (g6650), .I (g6213));
INVX1 gate1062(.O (g7169), .I (I13075));
INVX1 gate1063(.O (g7283), .I (I13281));
INVX1 gate1064(.O (g1572), .I (g673));
INVX1 gate1065(.O (g8955), .I (I15379));
INVX1 gate1066(.O (I6695), .I (g2246));
INVX1 gate1067(.O (g4541), .I (g2883));
INVX1 gate1068(.O (g7059), .I (g6538));
INVX1 gate1069(.O (g7920), .I (I14282));
INVX1 gate1070(.O (g7578), .I (I13879));
INVX1 gate1071(.O (g6008), .I (g5367));
INVX1 gate1072(.O (I11835), .I (g6181));
INVX1 gate1073(.O (g3691), .I (I7195));
INVX1 gate1074(.O (I11014), .I (g5621));
INVX1 gate1075(.O (g7459), .I (I13617));
INVX1 gate1076(.O (g9221), .I (I15937));
INVX1 gate1077(.O (I12205), .I (g6488));
INVX1 gate1078(.O (I9463), .I (g3942));
INVX1 gate1079(.O (g7718), .I (I14031));
INVX1 gate1080(.O (g7767), .I (I14172));
INVX1 gate1081(.O (g4153), .I (I8024));
INVX1 gate1082(.O (g4680), .I (I8945));
INVX1 gate1083(.O (I7688), .I (g3650));
INVX1 gate1084(.O (g6136), .I (I10773));
INVX1 gate1085(.O (g4353), .I (g3665));
INVX1 gate1086(.O (I11586), .I (g6256));
INVX1 gate1087(.O (I12912), .I (g7006));
INVX1 gate1088(.O (g6336), .I (I11335));
INVX1 gate1089(.O (I14100), .I (g7580));
INVX1 gate1090(.O (I6223), .I (g330));
INVX1 gate1091(.O (g8038), .I (g7694));
INVX1 gate1092(.O (g6768), .I (I12173));
INVX1 gate1093(.O (I8913), .I (g4306));
INVX1 gate1094(.O (g7582), .I (I13891));
INVX1 gate1095(.O (g6594), .I (I11796));
INVX1 gate1096(.O (g1961), .I (g1345));
INVX1 gate1097(.O (g3879), .I (g2963));
INVX1 gate1098(.O (g4802), .I (I9129));
INVX1 gate1099(.O (g7261), .I (I13225));
INVX1 gate1100(.O (I14683), .I (g7825));
INVX1 gate1101(.O (g3962), .I (g3131));
INVX1 gate1102(.O (g5151), .I (I9579));
INVX1 gate1103(.O (g7793), .I (I14234));
INVX1 gate1104(.O (g3158), .I (I6853));
INVX1 gate1105(.O (g3659), .I (g2293));
INVX1 gate1106(.O (g6806), .I (I12289));
INVX1 gate1107(.O (g5648), .I (g4748));
INVX1 gate1108(.O (I6416), .I (g1794));
INVX1 gate1109(.O (g3506), .I (g1781));
INVX1 gate1110(.O (g7015), .I (I12763));
INVX1 gate1111(.O (I12592), .I (g1008));
INVX1 gate1112(.O (g4558), .I (g2897));
INVX1 gate1113(.O (g9068), .I (I15598));
INVX1 gate1114(.O (I7126), .I (g2494));
INVX1 gate1115(.O (I5926), .I (g297));
INVX1 gate1116(.O (I7400), .I (g3075));
INVX1 gate1117(.O (I8859), .I (g3968));
INVX1 gate1118(.O (I7326), .I (g2940));
INVX1 gate1119(.O (I6115), .I (g134));
INVX1 gate1120(.O (I6251), .I (g489));
INVX1 gate1121(.O (g2921), .I (g2312));
INVX1 gate1122(.O (g6065), .I (I10684));
INVX1 gate1123(.O (g6887), .I (I12532));
INVX1 gate1124(.O (g6122), .I (I10752));
INVX1 gate1125(.O (I10882), .I (g5600));
INVX1 gate1126(.O (g6228), .I (I11021));
INVX1 gate1127(.O (I5754), .I (g966));
INVX1 gate1128(.O (g3587), .I (g1964));
INVX1 gate1129(.O (g6322), .I (I11293));
INVX1 gate1130(.O (I11275), .I (g5768));
INVX1 gate1131(.O (I9457), .I (g3940));
INVX1 gate1132(.O (g8918), .I (I15340));
INVX1 gate1133(.O (I16180), .I (g9387));
INVX1 gate1134(.O (g6230), .I (I11025));
INVX1 gate1135(.O (g7246), .I (I13196));
INVX1 gate1136(.O (g8967), .I (I15405));
INVX1 gate1137(.O (I13746), .I (g7311));
INVX1 gate1138(.O (I13493), .I (g7132));
INVX1 gate1139(.O (I9393), .I (g4266));
INVX1 gate1140(.O (g4511), .I (g2841));
INVX1 gate1141(.O (I15660), .I (g9062));
INVX1 gate1142(.O (g2895), .I (g2268));
INVX1 gate1143(.O (g6033), .I (g5384));
INVX1 gate1144(.O (g2837), .I (g1780));
INVX1 gate1145(.O (g7721), .I (g7344));
INVX1 gate1146(.O (g5839), .I (I10532));
INVX1 gate1147(.O (I9834), .I (g4782));
INVX1 gate1148(.O (g4092), .I (I7899));
INVX1 gate1149(.O (I13035), .I (g6964));
INVX1 gate1150(.O (g3985), .I (I7712));
INVX1 gate1151(.O (I12731), .I (g6579));
INVX1 gate1152(.O (I11806), .I (g6275));
INVX1 gate1153(.O (g4600), .I (I8715));
INVX1 gate1154(.O (I7383), .I (g3465));
INVX1 gate1155(.O (g4574), .I (g3466));
INVX1 gate1156(.O (g6096), .I (g5317));
INVX1 gate1157(.O (g6496), .I (I11662));
INVX1 gate1158(.O (g1679), .I (I5512));
INVX1 gate1159(.O (I8097), .I (g3237));
INVX1 gate1160(.O (g5172), .I (I9642));
INVX1 gate1161(.O (g5278), .I (I9794));
INVX1 gate1162(.O (g6845), .I (I12406));
INVX1 gate1163(.O (g7502), .I (I13682));
INVX1 gate1164(.O (I15550), .I (g9008));
INVX1 gate1165(.O (g9198), .I (g9187));
INVX1 gate1166(.O (g3545), .I (g2344));
INVX1 gate1167(.O (I8354), .I (g1163));
INVX1 gate1168(.O (g738), .I (I5404));
INVX1 gate1169(.O (g6195), .I (I10940));
INVX1 gate1170(.O (g5618), .I (g5015));
INVX1 gate1171(.O (g6137), .I (I10776));
INVX1 gate1172(.O (g6891), .I (I12544));
INVX1 gate1173(.O (g5143), .I (I9555));
INVX1 gate1174(.O (g1831), .I (g689));
INVX1 gate1175(.O (g6337), .I (I11338));
INVX1 gate1176(.O (g3591), .I (g1789));
INVX1 gate1177(.O (g3832), .I (I7299));
INVX1 gate1178(.O (g4580), .I (g2919));
INVX1 gate1179(.O (g9241), .I (I15971));
INVX1 gate1180(.O (I7588), .I (g2584));
INVX1 gate1181(.O (g3853), .I (I7362));
INVX1 gate1182(.O (I14725), .I (g8145));
INVX1 gate1183(.O (g7188), .I (I13106));
INVX1 gate1184(.O (g5988), .I (I10592));
INVX1 gate1185(.O (g2842), .I (g2209));
INVX1 gate1186(.O (I9938), .I (g4878));
INVX1 gate1187(.O (I10758), .I (g5662));
INVX1 gate1188(.O (g1805), .I (I5667));
INVX1 gate1189(.O (g6807), .I (I12292));
INVX1 gate1190(.O (g1916), .I (g775));
INVX1 gate1191(.O (g5693), .I (I10204));
INVX1 gate1192(.O (g7216), .I (I13152));
INVX1 gate1193(.O (g1749), .I (g371));
INVX1 gate1194(.O (g2298), .I (I6072));
INVX1 gate1195(.O (I14082), .I (g7539));
INVX1 gate1196(.O (g6859), .I (I12448));
INVX1 gate1197(.O (g2392), .I (g11));
INVX1 gate1198(.O (I13193), .I (g7007));
INVX1 gate1199(.O (g2485), .I (g62));
INVX1 gate1200(.O (I11362), .I (g5821));
INVX1 gate1201(.O (g7028), .I (g6525));
INVX1 gate1202(.O (I13362), .I (g7265));
INVX1 gate1203(.O (g3931), .I (I7592));
INVX1 gate1204(.O (I8218), .I (g3002));
INVX1 gate1205(.O (I15773), .I (g9126));
INVX1 gate1206(.O (I6629), .I (g2052));
INVX1 gate1207(.O (g4623), .I (I8784));
INVX1 gate1208(.O (g7247), .I (I13199));
INVX1 gate1209(.O (g1798), .I (I5654));
INVX1 gate1210(.O (I6130), .I (g560));
INVX1 gate1211(.O (g4076), .I (I7859));
INVX1 gate1212(.O (g9319), .I (g9309));
INVX1 gate1213(.O (I10940), .I (g5489));
INVX1 gate1214(.O (g2941), .I (g2349));
INVX1 gate1215(.O (I9606), .I (g4687));
INVX1 gate1216(.O (g6342), .I (I11353));
INVX1 gate1217(.O (g3905), .I (g3192));
INVX1 gate1218(.O (I13475), .I (g7125));
INVX1 gate1219(.O (g5621), .I (g4748));
INVX1 gate1220(.O (I14848), .I (g8625));
INVX1 gate1221(.O (g6255), .I (I11066));
INVX1 gate1222(.O (g6815), .I (I12316));
INVX1 gate1223(.O (I10804), .I (g5526));
INVX1 gate1224(.O (I6800), .I (g2016));
INVX1 gate1225(.O (I9687), .I (g4822));
INVX1 gate1226(.O (g3630), .I (I7095));
INVX1 gate1227(.O (g6481), .I (I11641));
INVX1 gate1228(.O (I14804), .I (g8563));
INVX1 gate1229(.O (g7741), .I (I14094));
INVX1 gate1230(.O (g4651), .I (I8868));
INVX1 gate1231(.O (g5113), .I (I9499));
INVX1 gate1232(.O (g6692), .I (I12008));
INVX1 gate1233(.O (g6097), .I (g5345));
INVX1 gate1234(.O (I11437), .I (g5801));
INVX1 gate1235(.O (I15839), .I (g9168));
INVX1 gate1236(.O (g2520), .I (g41));
INVX1 gate1237(.O (I15930), .I (g9209));
INVX1 gate1238(.O (g2640), .I (g1584));
INVX1 gate1239(.O (g9211), .I (I15909));
INVX1 gate1240(.O (g6354), .I (I11389));
INVX1 gate1241(.O (g4285), .I (I8233));
INVX1 gate1242(.O (I8727), .I (g3944));
INVX1 gate1243(.O (g9186), .I (I15836));
INVX1 gate1244(.O (I5679), .I (g911));
INVX1 gate1245(.O (g4500), .I (g2832));
INVX1 gate1246(.O (g9386), .I (I16176));
INVX1 gate1247(.O (g6960), .I (I12681));
INVX1 gate1248(.O (I15965), .I (g9219));
INVX1 gate1249(.O (I7944), .I (g3774));
INVX1 gate1250(.O (g1579), .I (g703));
INVX1 gate1251(.O (g1869), .I (g74));
INVX1 gate1252(.O (g7108), .I (I12912));
INVX1 gate1253(.O (I10135), .I (g4960));
INVX1 gate1254(.O (g7308), .I (I13356));
INVX1 gate1255(.O (I11347), .I (g5761));
INVX1 gate1256(.O (g2958), .I (g2377));
INVX1 gate1257(.O (I13347), .I (g7224));
INVX1 gate1258(.O (g9026), .I (I15492));
INVX1 gate1259(.O (I5831), .I (g1194));
INVX1 gate1260(.O (g2376), .I (I6226));
INVX1 gate1261(.O (g5494), .I (I9918));
INVX1 gate1262(.O (g3750), .I (g2177));
INVX1 gate1263(.O (I9570), .I (g4696));
INVX1 gate1264(.O (I10406), .I (g5203));
INVX1 gate1265(.O (I9341), .I (g4251));
INVX1 gate1266(.O (I10962), .I (g5719));
INVX1 gate1267(.O (g1752), .I (g603));
INVX1 gate1268(.O (I14406), .I (g7681));
INVX1 gate1269(.O (g3973), .I (g3097));
INVX1 gate1270(.O (I9525), .I (g4413));
INVX1 gate1271(.O (I11781), .I (g6284));
INVX1 gate1272(.O (I12768), .I (g6718));
INVX1 gate1273(.O (I15619), .I (g8998));
INVX1 gate1274(.O (g9370), .I (I16138));
INVX1 gate1275(.O (g1917), .I (I5795));
INVX1 gate1276(.O (I9645), .I (g4900));
INVX1 gate1277(.O (I15557), .I (g9010));
INVX1 gate1278(.O (g2829), .I (g1785));
INVX1 gate1279(.O (g9125), .I (I15753));
INVX1 gate1280(.O (g4024), .I (g3160));
INVX1 gate1281(.O (I11236), .I (g6148));
INVX1 gate1282(.O (g2286), .I (I6042));
INVX1 gate1283(.O (g6783), .I (I12220));
INVX1 gate1284(.O (g7758), .I (I14145));
INVX1 gate1285(.O (g7066), .I (I12839));
INVX1 gate1286(.O (I10500), .I (g5234));
INVX1 gate1287(.O (I16168), .I (g9381));
INVX1 gate1288(.O (g7589), .I (I13912));
INVX1 gate1289(.O (I6090), .I (g390));
INVX1 gate1290(.O (g2911), .I (g2292));
INVX1 gate1291(.O (g4795), .I (I9116));
INVX1 gate1292(.O (I8932), .I (g4096));
INVX1 gate1293(.O (I5422), .I (g1234));
INVX1 gate1294(.O (g7466), .I (I13622));
INVX1 gate1295(.O (g4809), .I (I9148));
INVX1 gate1296(.O (g6267), .I (I11086));
INVX1 gate1297(.O (g6312), .I (I11263));
INVX1 gate1298(.O (g3969), .I (g3192));
INVX1 gate1299(.O (I6166), .I (g480));
INVX1 gate1300(.O (I14049), .I (g7493));
INVX1 gate1301(.O (g9280), .I (I16006));
INVX1 gate1302(.O (I11821), .I (g6170));
INVX1 gate1303(.O (I12881), .I (g6478));
INVX1 gate1304(.O (g1786), .I (g623));
INVX1 gate1305(.O (g7365), .I (I13509));
INVX1 gate1306(.O (g7048), .I (I12810));
INVX1 gate1307(.O (I7347), .I (g2985));
INVX1 gate1308(.O (g9083), .I (I15641));
INVX1 gate1309(.O (g2270), .I (I6015));
INVX1 gate1310(.O (g4477), .I (I8517));
INVX1 gate1311(.O (g7448), .I (I13605));
INVX1 gate1312(.O (I13063), .I (g6973));
INVX1 gate1313(.O (g7711), .I (I14012));
INVX1 gate1314(.O (g4523), .I (g2868));
INVX1 gate1315(.O (g6676), .I (I11984));
INVX1 gate1316(.O (I11790), .I (g6282));
INVX1 gate1317(.O (g6293), .I (I11206));
INVX1 gate1318(.O (I13264), .I (g7061));
INVX1 gate1319(.O (I6148), .I (g5));
INVX1 gate1320(.O (g7055), .I (g6517));
INVX1 gate1321(.O (g8219), .I (I14436));
INVX1 gate1322(.O (g4643), .I (I8844));
INVX1 gate1323(.O (g3666), .I (g2134));
INVX1 gate1324(.O (I9158), .I (g4256));
INVX1 gate1325(.O (I13137), .I (g7027));
INVX1 gate1326(.O (I6348), .I (g1354));
INVX1 gate1327(.O (g2225), .I (I5948));
INVX1 gate1328(.O (g6129), .I (I10758));
INVX1 gate1329(.O (g8640), .I (I14728));
INVX1 gate1330(.O (g7455), .I (I13613));
INVX1 gate1331(.O (g6329), .I (I11314));
INVX1 gate1332(.O (g6761), .I (I12154));
INVX1 gate1333(.O (g2073), .I (g1254));
INVX1 gate1334(.O (g5160), .I (I9606));
INVX1 gate1335(.O (g7133), .I (I12983));
INVX1 gate1336(.O (I7697), .I (g3052));
INVX1 gate1337(.O (g9106), .I (I15708));
INVX1 gate1338(.O (g7333), .I (I13419));
INVX1 gate1339(.O (I13873), .I (g7342));
INVX1 gate1340(.O (g9306), .I (I16036));
INVX1 gate1341(.O (g6828), .I (I12355));
INVX1 gate1342(.O (g1770), .I (g606));
INVX1 gate1343(.O (g7774), .I (I14193));
INVX1 gate1344(.O (g5521), .I (g4929));
INVX1 gate1345(.O (g8958), .I (I15388));
INVX1 gate1346(.O (g6830), .I (I12361));
INVX1 gate1347(.O (g4634), .I (I8817));
INVX1 gate1348(.O (g3648), .I (g2424));
INVX1 gate1349(.O (g3875), .I (g2958));
INVX1 gate1350(.O (g2324), .I (I6115));
INVX1 gate1351(.O (g3530), .I (g2185));
INVX1 gate1352(.O (I9111), .I (g4232));
INVX1 gate1353(.O (g7196), .I (I13122));
INVX1 gate1354(.O (g4742), .I (I9064));
INVX1 gate1355(.O (g9061), .I (I15577));
INVX1 gate1356(.O (I15601), .I (g8992));
INVX1 gate1357(.O (g9187), .I (I15839));
INVX1 gate1358(.O (g4104), .I (I7925));
INVX1 gate1359(.O (I10605), .I (g5440));
INVX1 gate1360(.O (I11422), .I (g5842));
INVX1 gate1361(.O (g6592), .I (I11790));
INVX1 gate1362(.O (g3655), .I (g1844));
INVX1 gate1363(.O (I15187), .I (g8682));
INVX1 gate1364(.O (I14273), .I (g7631));
INVX1 gate1365(.O (I11209), .I (g6139));
INVX1 gate1366(.O (I13422), .I (g7131));
INVX1 gate1367(.O (I14106), .I (g7586));
INVX1 gate1368(.O (I13209), .I (g6912));
INVX1 gate1369(.O (g2540), .I (g1339));
INVX1 gate1370(.O (I9615), .I (g4739));
INVX1 gate1371(.O (g6221), .I (I11004));
INVX1 gate1372(.O (I12003), .I (g6202));
INVX1 gate1373(.O (g8765), .I (g8524));
INVX1 gate1374(.O (g7538), .I (I13794));
INVX1 gate1375(.O (I13834), .I (g7466));
INVX1 gate1376(.O (I6463), .I (g1769));
INVX1 gate1377(.O (I10463), .I (g5220));
INVX1 gate1378(.O (I16084), .I (g9324));
INVX1 gate1379(.O (g2177), .I (g1322));
INVX1 gate1380(.O (g7780), .I (I14211));
INVX1 gate1381(.O (g9027), .I (I15495));
INVX1 gate1382(.O (g5724), .I (g4969));
INVX1 gate1383(.O (g2377), .I (I6229));
INVX1 gate1384(.O (I14463), .I (g8072));
INVX1 gate1385(.O (I12779), .I (g6740));
INVX1 gate1386(.O (g5179), .I (I9663));
INVX1 gate1387(.O (g6703), .I (I12041));
INVX1 gate1388(.O (g7509), .I (I13707));
INVX1 gate1389(.O (g4926), .I (g4202));
INVX1 gate1390(.O (I15937), .I (g9212));
INVX1 gate1391(.O (g9200), .I (g9189));
INVX1 gate1392(.O (I11021), .I (g5627));
INVX1 gate1393(.O (I14234), .I (g7614));
INVX1 gate1394(.O (g3884), .I (I7417));
INVX1 gate1395(.O (g3839), .I (I7320));
INVX1 gate1396(.O (g2287), .I (I6045));
INVX1 gate1397(.O (g7018), .I (I12768));
INVX1 gate1398(.O (g4273), .I (I8215));
INVX1 gate1399(.O (g7067), .I (g6658));
INVX1 gate1400(.O (g8974), .I (I15426));
INVX1 gate1401(.O (I7317), .I (g2893));
INVX1 gate1402(.O (g5658), .I (g4748));
INVX1 gate1403(.O (I15791), .I (g9140));
INVX1 gate1404(.O (g7418), .I (I13533));
INVX1 gate1405(.O (g6624), .I (I11864));
INVX1 gate1406(.O (g7467), .I (g7236));
INVX1 gate1407(.O (g6953), .I (g6745));
INVX1 gate1408(.O (I6118), .I (g243));
INVX1 gate1409(.O (I14795), .I (g8604));
INVX1 gate1410(.O (g8225), .I (I14454));
INVX1 gate1411(.O (g5835), .I (I10528));
INVX1 gate1412(.O (g7290), .I (I13302));
INVX1 gate1413(.O (g4613), .I (I8754));
INVX1 gate1414(.O (g6068), .I (I10687));
INVX1 gate1415(.O (g1888), .I (g781));
INVX1 gate1416(.O (I6872), .I (g2185));
INVX1 gate1417(.O (g9145), .I (I15791));
INVX1 gate1418(.O (g4044), .I (g2595));
INVX1 gate1419(.O (g6468), .I (I11622));
INVX1 gate1420(.O (I12945), .I (g7066));
INVX1 gate1421(.O (I9591), .I (g4710));
INVX1 gate1422(.O (g4444), .I (I8452));
INVX1 gate1423(.O (g1787), .I (g625));
INVX1 gate1424(.O (I6652), .I (g2016));
INVX1 gate1425(.O (I11607), .I (g5767));
INVX1 gate1426(.O (I6057), .I (g518));
INVX1 gate1427(.O (I12826), .I (g6441));
INVX1 gate1428(.O (I12999), .I (g7029));
INVX1 gate1429(.O (I11320), .I (g5797));
INVX1 gate1430(.O (I15666), .I (g9070));
INVX1 gate1431(.O (I13320), .I (g7139));
INVX1 gate1432(.O (I6457), .I (g1886));
INVX1 gate1433(.O (g7493), .I (I13659));
INVX1 gate1434(.O (g1675), .I (g1519));
INVX1 gate1435(.O (g6677), .I (I11987));
INVX1 gate1436(.O (g7256), .I (g7058));
INVX1 gate1437(.O (I13274), .I (g6917));
INVX1 gate1438(.O (I7775), .I (g3705));
INVX1 gate1439(.O (g5611), .I (g4969));
INVX1 gate1440(.O (g8324), .I (I14573));
INVX1 gate1441(.O (g4572), .I (g2909));
INVX1 gate1442(.O (I7922), .I (g3462));
INVX1 gate1443(.O (g2898), .I (g2271));
INVX1 gate1444(.O (I15478), .I (g8910));
INVX1 gate1445(.O (g2900), .I (g2273));
INVX1 gate1446(.O (g6866), .I (I12469));
INVX1 gate1447(.O (I12672), .I (g6473));
INVX1 gate1448(.O (I7581), .I (g3612));
INVX1 gate1449(.O (I13122), .I (g7070));
INVX1 gate1450(.O (g9107), .I (I15711));
INVX1 gate1451(.O (g4543), .I (g2885));
INVX1 gate1452(.O (I10421), .I (g5208));
INVX1 gate1453(.O (I11464), .I (g6088));
INVX1 gate1454(.O (g5799), .I (I10436));
INVX1 gate1455(.O (I13565), .I (g7181));
INVX1 gate1456(.O (I9794), .I (g4778));
INVX1 gate1457(.O (I6834), .I (g287));
INVX1 gate1458(.O (g9307), .I (g9300));
INVX1 gate1459(.O (g2510), .I (g58));
INVX1 gate1460(.O (g639), .I (I5374));
INVX1 gate1461(.O (g2245), .I (g999));
INVX1 gate1462(.O (g6149), .I (I10810));
INVX1 gate1463(.O (g3988), .I (g3097));
INVX1 gate1464(.O (I6686), .I (g2246));
INVX1 gate1465(.O (g6349), .I (I11374));
INVX1 gate1466(.O (g5674), .I (g5042));
INVX1 gate1467(.O (g8177), .I (I14410));
INVX1 gate1468(.O (g3693), .I (g2424));
INVX1 gate1469(.O (I11034), .I (g5644));
INVX1 gate1470(.O (g9223), .I (I15943));
INVX1 gate1471(.O (I14163), .I (g7533));
INVX1 gate1472(.O (g2291), .I (I6057));
INVX1 gate1473(.O (I14012), .I (g7438));
INVX1 gate1474(.O (I11641), .I (g5918));
INVX1 gate1475(.O (g6848), .I (I12415));
INVX1 gate1476(.O (I15580), .I (g8985));
INVX1 gate1477(.O (I13797), .I (g7502));
INVX1 gate1478(.O (I12331), .I (g6704));
INVX1 gate1479(.O (g5541), .I (g4814));
INVX1 gate1480(.O (g3548), .I (g2185));
INVX1 gate1481(.O (g1684), .I (g1));
INVX1 gate1482(.O (g1745), .I (g746));
INVX1 gate1483(.O (g6198), .I (g5335));
INVX1 gate1484(.O (g1639), .I (g1207));
INVX1 gate1485(.O (g2344), .I (I6148));
INVX1 gate1486(.O (g6855), .I (I12436));
INVX1 gate1487(.O (g6398), .I (I11515));
INVX1 gate1488(.O (I10541), .I (g5256));
INVX1 gate1489(.O (I6121), .I (g321));
INVX1 gate1490(.O (g7263), .I (I13231));
INVX1 gate1491(.O (g2207), .I (I5920));
INVX1 gate1492(.O (g5153), .I (I9585));
INVX1 gate1493(.O (g5680), .I (g5101));
INVX1 gate1494(.O (I12897), .I (g6962));
INVX1 gate1495(.O (I12448), .I (g6569));
INVX1 gate1496(.O (I12961), .I (g6921));
INVX1 gate1497(.O (I9515), .I (g4301));
INVX1 gate1498(.O (I9630), .I (g4867));
INVX1 gate1499(.O (I14789), .I (g8544));
INVX1 gate1500(.O (g2259), .I (g1325));
INVX1 gate1501(.O (g9115), .I (I15735));
INVX1 gate1502(.O (g4014), .I (I7769));
INVX1 gate1503(.O (I7079), .I (g2532));
INVX1 gate1504(.O (I12505), .I (g6612));
INVX1 gate1505(.O (g9315), .I (I16061));
INVX1 gate1506(.O (g1808), .I (g629));
INVX1 gate1507(.O (g4885), .I (g4070));
INVX1 gate1508(.O (I13635), .I (g7243));
INVX1 gate1509(.O (g5744), .I (I10289));
INVX1 gate1510(.O (g8199), .I (I14424));
INVX1 gate1511(.O (g9047), .I (I15543));
INVX1 gate1512(.O (g5802), .I (I10445));
INVX1 gate1513(.O (g4660), .I (I8895));
INVX1 gate1514(.O (g2923), .I (I6657));
INVX1 gate1515(.O (I12717), .I (g6543));
INVX1 gate1516(.O (g1707), .I (g955));
INVX1 gate1517(.O (I14325), .I (g7713));
INVX1 gate1518(.O (I10829), .I (g5224));
INVX1 gate1519(.O (g8781), .I (g8585));
INVX1 gate1520(.O (I10535), .I (g5254));
INVX1 gate1521(.O (I5389), .I (g690));
INVX1 gate1522(.O (I5706), .I (g901));
INVX1 gate1523(.O (g8898), .I (I15308));
INVX1 gate1524(.O (g4903), .I (g4084));
INVX1 gate1525(.O (g7562), .I (I13858));
INVX1 gate1526(.O (I15178), .I (g8753));
INVX1 gate1527(.O (I10946), .I (g5563));
INVX1 gate1528(.O (g8797), .I (I15003));
INVX1 gate1529(.O (g6524), .I (I11710));
INVX1 gate1530(.O (I14828), .I (g8639));
INVX1 gate1531(.O (g6644), .I (g6208));
INVX1 gate1532(.O (g8510), .I (I14643));
INVX1 gate1533(.O (I13164), .I (g7086));
INVX1 gate1534(.O (I5371), .I (g633));
INVX1 gate1535(.O (g7723), .I (I14042));
INVX1 gate1536(.O (I14121), .I (g7587));
INVX1 gate1537(.O (g2215), .I (g1416));
INVX1 gate1538(.O (I15953), .I (g9215));
INVX1 gate1539(.O (g6319), .I (I11284));
INVX1 gate1540(.O (g7101), .I (I12891));
INVX1 gate1541(.O (g2886), .I (g2240));
INVX1 gate1542(.O (g3908), .I (I7517));
INVX1 gate1543(.O (g7301), .I (I13335));
INVX1 gate1544(.O (I7356), .I (g2843));
INVX1 gate1545(.O (I13891), .I (g7336));
INVX1 gate1546(.O (I15654), .I (g9057));
INVX1 gate1547(.O (g4036), .I (g3192));
INVX1 gate1548(.O (g6152), .I (I10815));
INVX1 gate1549(.O (g6258), .I (g5427));
INVX1 gate1550(.O (g6352), .I (I11383));
INVX1 gate1551(.O (g6818), .I (I12325));
INVX1 gate1552(.O (g1575), .I (g685));
INVX1 gate1553(.O (g1865), .I (g1013));
INVX1 gate1554(.O (I8483), .I (g3641));
INVX1 gate1555(.O (g6867), .I (I12472));
INVX1 gate1556(.O (g3567), .I (g2407));
INVX1 gate1557(.O (I15417), .I (g8893));
INVX1 gate1558(.O (g1715), .I (I5559));
INVX1 gate1559(.O (g2314), .I (I6099));
INVX1 gate1560(.O (I9440), .I (g4285));
INVX1 gate1561(.O (I14291), .I (g7680));
INVX1 gate1562(.O (I12433), .I (g6632));
INVX1 gate1563(.O (g4335), .I (g3659));
INVX1 gate1564(.O (I9123), .I (g4455));
INVX1 gate1565(.O (I15334), .I (g8800));
INVX1 gate1566(.O (g7751), .I (I14124));
INVX1 gate1567(.O (g2870), .I (g2225));
INVX1 gate1568(.O (g5492), .I (g4919));
INVX1 gate1569(.O (I12148), .I (g5988));
INVX1 gate1570(.O (I13109), .I (g7059));
INVX1 gate1571(.O (g4382), .I (I8373));
INVX1 gate1572(.O (g1833), .I (g770));
INVX1 gate1573(.O (g5600), .I (g5128));
INVX1 gate1574(.O (I13537), .I (g7152));
INVX1 gate1575(.O (g5574), .I (g4969));
INVX1 gate1576(.O (I8790), .I (g4020));
INVX1 gate1577(.O (g6211), .I (g5645));
INVX1 gate1578(.O (g2825), .I (I6553));
INVX1 gate1579(.O (g2650), .I (I6434));
INVX1 gate1580(.O (g6186), .I (I10919));
INVX1 gate1581(.O (g6386), .I (I11485));
INVX1 gate1582(.O (I12646), .I (g6493));
INVX1 gate1583(.O (g7585), .I (I13900));
INVX1 gate1584(.O (g9017), .I (I15475));
INVX1 gate1585(.O (I9666), .I (g4931));
INVX1 gate1586(.O (I15762), .I (g9039));
INVX1 gate1587(.O (I12343), .I (g6731));
INVX1 gate1588(.O (g4805), .I (I9136));
INVX1 gate1589(.O (g6975), .I (I12712));
INVX1 gate1590(.O (g4916), .I (g4202));
INVX1 gate1591(.O (g4022), .I (I7785));
INVX1 gate1592(.O (g3965), .I (I7676));
INVX1 gate1593(.O (I5963), .I (g225));
INVX1 gate1594(.O (g1584), .I (g738));
INVX1 gate1595(.O (g6599), .I (I11809));
INVX1 gate1596(.O (g1896), .I (g86));
INVX1 gate1597(.O (g7441), .I (I13580));
INVX1 gate1598(.O (I15423), .I (g8894));
INVX1 gate1599(.O (g6026), .I (g5384));
INVX1 gate1600(.O (I9528), .I (g4006));
INVX1 gate1601(.O (g6426), .I (I11559));
INVX1 gate1602(.O (I6860), .I (g2185));
INVX1 gate1603(.O (g3264), .I (I6900));
INVX1 gate1604(.O (I7053), .I (g2452));
INVX1 gate1605(.O (I6341), .I (g1351));
INVX1 gate1606(.O (I10506), .I (g5236));
INVX1 gate1607(.O (g5580), .I (g4938));
INVX1 gate1608(.O (I9648), .I (g4795));
INVX1 gate1609(.O (g9234), .I (I15956));
INVX1 gate1610(.O (I10028), .I (g4825));
INVX1 gate1611(.O (g9128), .I (I15762));
INVX1 gate1612(.O (g6614), .I (I11838));
INVX1 gate1613(.O (g6370), .I (I11437));
INVX1 gate1614(.O (I14028), .I (g7501));
INVX1 gate1615(.O (g3933), .I (g3131));
INVX1 gate1616(.O (I8904), .I (g4126));
INVX1 gate1617(.O (g9330), .I (g9319));
INVX1 gate1618(.O (g6325), .I (I11302));
INVX1 gate1619(.O (g6821), .I (I12334));
INVX1 gate1620(.O (g3521), .I (g2185));
INVX1 gate1621(.O (g4560), .I (g2899));
INVX1 gate1622(.O (I8446), .I (g3014));
INVX1 gate1623(.O (g3050), .I (I6788));
INVX1 gate1624(.O (g3641), .I (I7115));
INVX1 gate1625(.O (I15909), .I (g9201));
INVX1 gate1626(.O (I15543), .I (g9006));
INVX1 gate1627(.O (g5736), .I (I10265));
INVX1 gate1628(.O (g2943), .I (g2362));
INVX1 gate1629(.O (g6984), .I (I12725));
INVX1 gate1630(.O (g7168), .I (I13072));
INVX1 gate1631(.O (g6939), .I (g6543));
INVX1 gate1632(.O (g3996), .I (I7731));
INVX1 gate1633(.O (I11796), .I (g6287));
INVX1 gate1634(.O (I12412), .I (g6404));
INVX1 gate1635(.O (I8841), .I (g3979));
INVX1 gate1636(.O (g5623), .I (g4969));
INVX1 gate1637(.O (g7772), .I (I14187));
INVX1 gate1638(.O (g6083), .I (I10702));
INVX1 gate1639(.O (g7058), .I (g6649));
INVX1 gate1640(.O (I5957), .I (g110));
INVX1 gate1641(.O (g2887), .I (g2241));
INVX1 gate1642(.O (g4873), .I (I9217));
INVX1 gate1643(.O (g4632), .I (I8811));
INVX1 gate1644(.O (g7531), .I (I13773));
INVX1 gate1645(.O (g4095), .I (I7908));
INVX1 gate1646(.O (g5076), .I (I9446));
INVX1 gate1647(.O (g8870), .I (I15196));
INVX1 gate1648(.O (I8763), .I (g3947));
INVX1 gate1649(.O (g4037), .I (g2845));
INVX1 gate1650(.O (g6483), .I (I11645));
INVX1 gate1651(.O (I12229), .I (g6659));
INVX1 gate1652(.O (I9884), .I (g4868));
INVX1 gate1653(.O (g2934), .I (I6676));
INVX1 gate1654(.O (g5476), .I (g4907));
INVX1 gate1655(.O (g7743), .I (I14100));
INVX1 gate1656(.O (g4653), .I (I8874));
INVX1 gate1657(.O (I6358), .I (g13));
INVX1 gate1658(.O (g4102), .I (I7919));
INVX1 gate1659(.O (g6636), .I (I11900));
INVX1 gate1660(.O (I15568), .I (g8981));
INVX1 gate1661(.O (I15747), .I (g9042));
INVX1 gate1662(.O (I5865), .I (g1206));
INVX1 gate1663(.O (g9213), .I (I15915));
INVX1 gate1664(.O (g6106), .I (g5345));
INVX1 gate1665(.O (g5175), .I (I9651));
INVX1 gate1666(.O (g4579), .I (g2918));
INVX1 gate1667(.O (I10649), .I (g5657));
INVX1 gate1668(.O (I12011), .I (g5939));
INVX1 gate1669(.O (g6306), .I (I11245));
INVX1 gate1670(.O (I5715), .I (g896));
INVX1 gate1671(.O (g7505), .I (I13695));
INVX1 gate1672(.O (g5871), .I (I10558));
INVX1 gate1673(.O (g3878), .I (g2962));
INVX1 gate1674(.O (g8008), .I (g7559));
INVX1 gate1675(.O (g4719), .I (I9021));
INVX1 gate1676(.O (g6790), .I (I12241));
INVX1 gate1677(.O (g7734), .I (I14073));
INVX1 gate1678(.O (I6587), .I (g1708));
INVX1 gate1679(.O (g3777), .I (g2170));
INVX1 gate1680(.O (g7411), .I (g7202));
INVX1 gate1681(.O (I9372), .I (g3902));
INVX1 gate1682(.O (I10491), .I (g5231));
INVX1 gate1683(.O (I15814), .I (g9154));
INVX1 gate1684(.O (g3835), .I (I7308));
INVX1 gate1685(.O (I16116), .I (g9350));
INVX1 gate1686(.O (g6387), .I (I11488));
INVX1 gate1687(.O (I11522), .I (g5847));
INVX1 gate1688(.O (g2096), .I (g1226));
INVX1 gate1689(.O (I9618), .I (g4742));
INVX1 gate1690(.O (I12582), .I (g6745));
INVX1 gate1691(.O (g5285), .I (g4841));
INVX1 gate1692(.O (g6461), .I (I11607));
INVX1 gate1693(.O (g8768), .I (g8585));
INVX1 gate1694(.O (I13663), .I (g7235));
INVX1 gate1695(.O (g3882), .I (g2970));
INVX1 gate1696(.O (g2496), .I (g942));
INVX1 gate1697(.O (I7626), .I (g3632));
INVX1 gate1698(.O (g4917), .I (g4102));
INVX1 gate1699(.O (I15974), .I (g9234));
INVX1 gate1700(.O (I6615), .I (g1983));
INVX1 gate1701(.O (g6756), .I (I12141));
INVX1 gate1702(.O (g8972), .I (I15420));
INVX1 gate1703(.O (I10770), .I (g5441));
INVX1 gate1704(.O (I12310), .I (g6723));
INVX1 gate1705(.O (g1897), .I (g789));
INVX1 gate1706(.O (g9090), .I (I15660));
INVX1 gate1707(.O (g6622), .I (I11858));
INVX1 gate1708(.O (g7474), .I (I13628));
INVX1 gate1709(.O (I8757), .I (g3921));
INVX1 gate1710(.O (g6027), .I (g5384));
INVX1 gate1711(.O (g7992), .I (g7557));
INVX1 gate1712(.O (g4265), .I (g3591));
INVX1 gate1713(.O (g3611), .I (I7079));
INVX1 gate1714(.O (g6427), .I (I11562));
INVX1 gate1715(.O (g2137), .I (I5889));
INVX1 gate1716(.O (g2891), .I (g2265));
INVX1 gate1717(.O (g5184), .I (I9678));
INVX1 gate1718(.O (I15638), .I (g8978));
INVX1 gate1719(.O (g9366), .I (I16126));
INVX1 gate1720(.O (g2913), .I (g2307));
INVX1 gate1721(.O (I12379), .I (g6768));
INVX1 gate1722(.O (g5139), .I (I9543));
INVX1 gate1723(.O (g5384), .I (I9837));
INVX1 gate1724(.O (g6904), .I (g6426));
INVX1 gate1725(.O (I12958), .I (g6920));
INVX1 gate1726(.O (g9056), .I (I15562));
INVX1 gate1727(.O (g8065), .I (I14338));
INVX1 gate1728(.O (I8315), .I (g3691));
INVX1 gate1729(.O (I8811), .I (g4022));
INVX1 gate1730(.O (g6446), .I (I11591));
INVX1 gate1731(.O (g8228), .I (I14463));
INVX1 gate1732(.O (g3981), .I (I7706));
INVX1 gate1733(.O (g5024), .I (I9360));
INVX1 gate1734(.O (g6514), .I (I11696));
INVX1 gate1735(.O (I6239), .I (g8));
INVX1 gate1736(.O (g3674), .I (I7164));
INVX1 gate1737(.O (g2807), .I (g1782));
INVX1 gate1738(.O (I5362), .I (g3841));
INVX1 gate1739(.O (I11326), .I (g5819));
INVX1 gate1740(.O (I9555), .I (g4892));
INVX1 gate1741(.O (g5795), .I (I10424));
INVX1 gate1742(.O (g5737), .I (I10268));
INVX1 gate1743(.O (I15391), .I (g8917));
INVX1 gate1744(.O (g6403), .I (I11522));
INVX1 gate1745(.O (I13326), .I (g7176));
INVX1 gate1746(.O (g5809), .I (I10460));
INVX1 gate1747(.O (I5419), .I (g1603));
INVX1 gate1748(.O (I9804), .I (g5113));
INVX1 gate1749(.O (I10262), .I (g5551));
INVX1 gate1750(.O (I7683), .I (g2573));
INVX1 gate1751(.O (g3997), .I (I7734));
INVX1 gate1752(.O (I12742), .I (g6590));
INVX1 gate1753(.O (g6345), .I (I11362));
INVX1 gate1754(.O (g6841), .I (I12394));
INVX1 gate1755(.O (I15510), .I (g8969));
INVX1 gate1756(.O (I11040), .I (g5299));
INVX1 gate1757(.O (I11948), .I (g5897));
INVX1 gate1758(.O (I8874), .I (g3884));
INVX1 gate1759(.O (g2266), .I (I6003));
INVX1 gate1760(.O (g6763), .I (I12158));
INVX1 gate1761(.O (I7778), .I (g3019));
INVX1 gate1762(.O (I16142), .I (g9366));
INVX1 gate1763(.O (g6391), .I (I11500));
INVX1 gate1764(.O (g1006), .I (I5410));
INVX1 gate1765(.O (g4296), .I (g3790));
INVX1 gate1766(.O (I6853), .I (g2185));
INVX1 gate1767(.O (g3238), .I (I6894));
INVX1 gate1768(.O (I9621), .I (g4732));
INVX1 gate1769(.O (g5477), .I (g4908));
INVX1 gate1770(.O (g9260), .I (I15990));
INVX1 gate1771(.O (g5523), .I (I9935));
INVX1 gate1772(.O (I12681), .I (g6469));
INVX1 gate1773(.O (I10719), .I (g5559));
INVX1 gate1774(.O (g6637), .I (I11903));
INVX1 gate1775(.O (g5643), .I (I10128));
INVX1 gate1776(.O (I15014), .I (g8607));
INVX1 gate1777(.O (g1801), .I (g618));
INVX1 gate1778(.O (g4553), .I (g2891));
INVX1 gate1779(.O (g9063), .I (I15583));
INVX1 gate1780(.O (g6307), .I (I11248));
INVX1 gate1781(.O (I15586), .I (g8987));
INVX1 gate1782(.O (I15007), .I (g8627));
INVX1 gate1783(.O (I8880), .I (g4303));
INVX1 gate1784(.O (I14718), .I (g8068));
INVX1 gate1785(.O (g3802), .I (g1832));
INVX1 gate1786(.O (g7688), .I (g7406));
INVX1 gate1787(.O (g6359), .I (I11404));
INVX1 gate1788(.O (g6223), .I (I11008));
INVX1 gate1789(.O (g2481), .I (I6317));
INVX1 gate1790(.O (g8913), .I (I15329));
INVX1 gate1791(.O (g1748), .I (g601));
INVX1 gate1792(.O (g2692), .I (g1671));
INVX1 gate1793(.O (g4012), .I (I7765));
INVX1 gate1794(.O (g6858), .I (I12445));
INVX1 gate1795(.O (g5742), .I (I10283));
INVX1 gate1796(.O (g5551), .I (I9974));
INVX1 gate1797(.O (g5099), .I (g4477));
INVX1 gate1798(.O (g2497), .I (g945));
INVX1 gate1799(.O (I12690), .I (g6467));
INVX1 gate1800(.O (g2354), .I (I6178));
INVX1 gate1801(.O (I16165), .I (g9377));
INVX1 gate1802(.O (g2960), .I (g2381));
INVX1 gate1803(.O (g4706), .I (I9005));
INVX1 gate1804(.O (I9567), .I (g4693));
INVX1 gate1805(.O (I7526), .I (g2752));
INVX1 gate1806(.O (I5897), .I (g173));
INVX1 gate1807(.O (I14573), .I (g8179));
INVX1 gate1808(.O (I10247), .I (g5266));
INVX1 gate1809(.O (g3901), .I (I7492));
INVX1 gate1810(.O (g7000), .I (I12742));
INVX1 gate1811(.O (I13509), .I (g7137));
INVX1 gate1812(.O (I15720), .I (g9053));
INVX1 gate1813(.O (g9318), .I (g9304));
INVX1 gate1814(.O (g9367), .I (I16129));
INVX1 gate1815(.O (I11933), .I (g5847));
INVX1 gate1816(.O (g7126), .I (I12968));
INVX1 gate1817(.O (I8935), .I (g4005));
INVX1 gate1818(.O (I5425), .I (g1245));
INVX1 gate1819(.O (g4029), .I (I7800));
INVX1 gate1820(.O (g6251), .I (I11060));
INVX1 gate1821(.O (g6315), .I (I11272));
INVX1 gate1822(.O (g6811), .I (I12304));
INVX1 gate1823(.O (g6642), .I (I11912));
INVX1 gate1824(.O (g4371), .I (I8354));
INVX1 gate1825(.O (I11851), .I (g6277));
INVX1 gate1826(.O (g3511), .I (g1616));
INVX1 gate1827(.O (g5754), .I (g5403));
INVX1 gate1828(.O (g9057), .I (I15565));
INVX1 gate1829(.O (I16006), .I (g9261));
INVX1 gate1830(.O (g7760), .I (I14151));
INVX1 gate1831(.O (I14388), .I (g7605));
INVX1 gate1832(.O (I7850), .I (g2795));
INVX1 gate1833(.O (g9193), .I (g9181));
INVX1 gate1834(.O (g3092), .I (I6826));
INVX1 gate1835(.O (I14777), .I (g8511));
INVX1 gate1836(.O (g3492), .I (I6970));
INVX1 gate1837(.O (g4281), .I (g2562));
INVX1 gate1838(.O (g6874), .I (I12493));
INVX1 gate1839(.O (g5613), .I (g4748));
INVX1 gate1840(.O (I14251), .I (g7541));
INVX1 gate1841(.O (g3574), .I (g1771));
INVX1 gate1842(.O (g3864), .I (g2943));
INVX1 gate1843(.O (g8342), .I (g8008));
INVX1 gate1844(.O (I15340), .I (g8856));
INVX1 gate1845(.O (g2267), .I (I6006));
INVX1 gate1846(.O (g2312), .I (I6093));
INVX1 gate1847(.O (g6654), .I (I11942));
INVX1 gate1848(.O (g5444), .I (g5074));
INVX1 gate1849(.O (g5269), .I (I9791));
INVX1 gate1850(.O (I7702), .I (g3062));
INVX1 gate1851(.O (I15684), .I (g9067));
INVX1 gate1852(.O (g8481), .I (I14637));
INVX1 gate1853(.O (I12128), .I (g5897));
INVX1 gate1854(.O (g1578), .I (g699));
INVX1 gate1855(.O (g1868), .I (I5747));
INVX1 gate1856(.O (I9360), .I (g4257));
INVX1 gate1857(.O (g2401), .I (g22));
INVX1 gate1858(.O (I7919), .I (g3761));
INVX1 gate1859(.O (I10032), .I (g1236));
INVX1 gate1860(.O (g1718), .I (I5562));
INVX1 gate1861(.O (g7779), .I (I14208));
INVX1 gate1862(.O (g2293), .I (g888));
INVX1 gate1863(.O (g6880), .I (I12511));
INVX1 gate1864(.O (g4684), .I (I8949));
INVX1 gate1865(.O (I9050), .I (g3881));
INVX1 gate1866(.O (I11452), .I (g6071));
INVX1 gate1867(.O (g6595), .I (g6083));
INVX1 gate1868(.O (g4639), .I (I8832));
INVX1 gate1869(.O (I5682), .I (g168));
INVX1 gate1870(.O (I5766), .I (g1254));
INVX1 gate1871(.O (I11047), .I (g5653));
INVX1 gate1872(.O (I13574), .I (g7205));
INVX1 gate1873(.O (g2329), .I (I6130));
INVX1 gate1874(.O (I6440), .I (g1806));
INVX1 gate1875(.O (g7023), .I (I12779));
INVX1 gate1876(.O (g9121), .I (I15747));
INVX1 gate1877(.O (g4963), .I (g4328));
INVX1 gate1878(.O (g2761), .I (g1820));
INVX1 gate1879(.O (I5801), .I (g1424));
INVX1 gate1880(.O (g9321), .I (g9311));
INVX1 gate1881(.O (g8960), .I (I15394));
INVX1 gate1882(.O (g7423), .I (I13544));
INVX1 gate1883(.O (g1582), .I (g714));
INVX1 gate1884(.O (I11912), .I (g5897));
INVX1 gate1885(.O (I11311), .I (g5760));
INVX1 gate1886(.O (I13912), .I (g7359));
INVX1 gate1887(.O (I13311), .I (g7162));
INVX1 gate1888(.O (g2828), .I (g1980));
INVX1 gate1889(.O (I12298), .I (g6697));
INVX1 gate1890(.O (I6323), .I (g1342));
INVX1 gate1891(.O (I14061), .I (g7546));
INVX1 gate1892(.O (g1793), .I (g626));
INVX1 gate1893(.O (I7561), .I (g2562));
INVX1 gate1894(.O (g7588), .I (I13909));
INVX1 gate1895(.O (I10766), .I (g5674));
INVX1 gate1896(.O (g2727), .I (g2424));
INVX1 gate1897(.O (g4808), .I (I9145));
INVX1 gate1898(.O (g6978), .I (I12717));
INVX1 gate1899(.O (g6612), .I (I11832));
INVX1 gate1900(.O (g7161), .I (I13057));
INVX1 gate1901(.O (g1015), .I (I5416));
INVX1 gate1902(.O (g5729), .I (g5144));
INVX1 gate1903(.O (g3968), .I (I7683));
INVX1 gate1904(.O (g6243), .I (I11050));
INVX1 gate1905(.O (g7361), .I (I13499));
INVX1 gate1906(.O (I15193), .I (g8774));
INVX1 gate1907(.O (I13051), .I (g6967));
INVX1 gate1908(.O (I13072), .I (g6969));
INVX1 gate1909(.O (g2746), .I (g2259));
INVX1 gate1910(.O (I12737), .I (g6460));
INVX1 gate1911(.O (g2221), .I (I5936));
INVX1 gate1912(.O (g3076), .I (g1831));
INVX1 gate1913(.O (g7127), .I (g6974));
INVX1 gate1914(.O (g8783), .I (g8524));
INVX1 gate1915(.O (g7327), .I (I13403));
INVX1 gate1916(.O (I12232), .I (g6662));
INVX1 gate1917(.O (g1664), .I (g1462));
INVX1 gate1918(.O (I6151), .I (g12));
INVX1 gate1919(.O (g1246), .I (I5425));
INVX1 gate1920(.O (g2703), .I (g1809));
INVX1 gate1921(.O (g8218), .I (I14433));
INVX1 gate1922(.O (I8823), .I (g3965));
INVX1 gate1923(.O (g5014), .I (I9344));
INVX1 gate1924(.O (g206), .I (I5353));
INVX1 gate1925(.O (g6328), .I (I11311));
INVX1 gate1926(.O (g6130), .I (I10761));
INVX1 gate1927(.O (g7146), .I (g6998));
INVX1 gate1928(.O (g6542), .I (I11718));
INVX1 gate1929(.O (g6330), .I (I11317));
INVX1 gate1930(.O (g7346), .I (I13454));
INVX1 gate1931(.O (g7633), .I (I13962));
INVX1 gate1932(.O (g1721), .I (I5565));
INVX1 gate1933(.O (I11350), .I (g5763));
INVX1 gate1934(.O (g3871), .I (g2953));
INVX1 gate1935(.O (I7970), .I (g3557));
INVX1 gate1936(.O (I13350), .I (g7223));
INVX1 gate1937(.O (I15475), .I (g8901));
INVX1 gate1938(.O (g2932), .I (g2329));
INVX1 gate1939(.O (g7103), .I (I12897));
INVX1 gate1940(.O (I9271), .I (g4263));
INVX1 gate1941(.O (g3651), .I (I7129));
INVX1 gate1942(.O (g7303), .I (I13341));
INVX1 gate1943(.O (I7925), .I (g2761));
INVX1 gate1944(.O (g8676), .I (I14822));
INVX1 gate1945(.O (g2624), .I (g1569));
INVX1 gate1946(.O (g2953), .I (g2373));
INVX1 gate1947(.O (I15222), .I (g8834));
INVX1 gate1948(.O (g6800), .I (I12271));
INVX1 gate1949(.O (g3285), .I (g1689));
INVX1 gate1950(.O (I13152), .I (g6966));
INVX1 gate1951(.O (g8761), .I (g8564));
INVX1 gate1952(.O (g4604), .I (I8727));
INVX1 gate1953(.O (I10451), .I (g5216));
INVX1 gate1954(.O (I10472), .I (g5223));
INVX1 gate1955(.O (I13846), .I (g7487));
INVX1 gate1956(.O (g3500), .I (g1616));
INVX1 gate1957(.O (I14451), .I (g8172));
INVX1 gate1958(.O (g7732), .I (I14067));
INVX1 gate1959(.O (I5407), .I (g4653));
INVX1 gate1960(.O (I13731), .I (g7441));
INVX1 gate1961(.O (I5920), .I (g219));
INVX1 gate1962(.O (I6839), .I (g2185));
INVX1 gate1963(.O (I5868), .I (g74));
INVX1 gate1964(.O (I7320), .I (g2927));
INVX1 gate1965(.O (g2677), .I (g1664));
INVX1 gate1966(.O (g7753), .I (I14130));
INVX1 gate1967(.O (g5178), .I (I9660));
INVX1 gate1968(.O (g5679), .I (I10172));
INVX1 gate1969(.O (I11413), .I (g5871));
INVX1 gate1970(.O (I5718), .I (g896));
INVX1 gate1971(.O (g7508), .I (I13704));
INVX1 gate1972(.O (I13413), .I (g7127));
INVX1 gate1973(.O (g6213), .I (I10976));
INVX1 gate1974(.O (I5535), .I (g48));
INVX1 gate1975(.O (g2866), .I (g2221));
INVX1 gate1976(.O (g4584), .I (g3466));
INVX1 gate1977(.O (I12445), .I (g6568));
INVX1 gate1978(.O (g4539), .I (g2881));
INVX1 gate1979(.O (g8746), .I (g8524));
INVX1 gate1980(.O (g8221), .I (I14442));
INVX1 gate1981(.O (g5335), .I (g4677));
INVX1 gate1982(.O (g5831), .I (I10516));
INVX1 gate1983(.O (g3838), .I (I7317));
INVX1 gate1984(.O (g1689), .I (g855));
INVX1 gate1985(.O (g2149), .I (I5894));
INVX1 gate1986(.O (g2349), .I (I6163));
INVX1 gate1987(.O (I12499), .I (g6597));
INVX1 gate1988(.O (g7043), .I (g6543));
INVX1 gate1989(.O (g9141), .I (g9129));
INVX1 gate1990(.O (g5182), .I (I9672));
INVX1 gate1991(.O (I10776), .I (g5576));
INVX1 gate1992(.O (I12316), .I (g6736));
INVX1 gate1993(.O (I9132), .I (g4284));
INVX1 gate1994(.O (I6143), .I (g1217));
INVX1 gate1995(.O (I9209), .I (g4349));
INVX1 gate1996(.O (g7116), .I (I12936));
INVX1 gate1997(.O (g1671), .I (g1494));
INVX1 gate1998(.O (I7987), .I (g3528));
INVX1 gate1999(.O (g5805), .I (I10448));
INVX1 gate2000(.O (g5916), .I (g5384));
INVX1 gate2001(.O (g5022), .I (g4438));
INVX1 gate2002(.O (g2699), .I (g1674));
INVX1 gate2003(.O (g4019), .I (I7778));
INVX1 gate2004(.O (g6090), .I (g5529));
INVX1 gate2005(.O (g4362), .I (g2810));
INVX1 gate2006(.O (I11929), .I (g6190));
INVX1 gate2007(.O (I12989), .I (g6932));
INVX1 gate2008(.O (g3077), .I (I6805));
INVX1 gate2009(.O (g7034), .I (g6525));
INVX1 gate2010(.O (g5749), .I (g5207));
INVX1 gate2011(.O (g6490), .I (I11656));
INVX1 gate2012(.O (g6823), .I (I12340));
INVX1 gate2013(.O (g7434), .I (I13565));
INVX1 gate2014(.O (I14825), .I (g8651));
INVX1 gate2015(.O (g3523), .I (g2407));
INVX1 gate2016(.O (I14370), .I (g7603));
INVX1 gate2017(.O (g6366), .I (I11425));
INVX1 gate2018(.O (I12722), .I (g6611));
INVX1 gate2019(.O (g7565), .I (I13865));
INVX1 gate2020(.O (I7299), .I (g2961));
INVX1 gate2021(.O (I5664), .I (g916));
INVX1 gate2022(.O (g3643), .I (g2453));
INVX1 gate2023(.O (I12924), .I (g6983));
INVX1 gate2024(.O (I13583), .I (g7252));
INVX1 gate2025(.O (g2241), .I (I5984));
INVX1 gate2026(.O (g1564), .I (g642));
INVX1 gate2027(.O (g7147), .I (g6904));
INVX1 gate2028(.O (I16122), .I (g9353));
INVX1 gate2029(.O (I10151), .I (g5007));
INVX1 gate2030(.O (I10172), .I (g4873));
INVX1 gate2031(.O (g7347), .I (I13457));
INVX1 gate2032(.O (I15516), .I (g8977));
INVX1 gate2033(.O (I9558), .I (g4597));
INVX1 gate2034(.O (g5798), .I (I10433));
INVX1 gate2035(.O (I14151), .I (g7555));
INVX1 gate2036(.O (g1826), .I (g632));
INVX1 gate2037(.O (I12271), .I (g6663));
INVX1 gate2038(.O (I14172), .I (g7545));
INVX1 gate2039(.O (g6148), .I (I10807));
INVX1 gate2040(.O (g6649), .I (I11929));
INVX1 gate2041(.O (I14996), .I (g8510));
INVX1 gate2042(.O (g6348), .I (I11371));
INVX1 gate2043(.O (I8989), .I (g4537));
INVX1 gate2044(.O (g8677), .I (I14825));
INVX1 gate2045(.O (g7533), .I (I13779));
INVX1 gate2046(.O (g3634), .I (I7107));
INVX1 gate2047(.O (I8193), .I (g3547));
INVX1 gate2048(.O (g6155), .I (I10826));
INVX1 gate2049(.O (I14844), .I (g8641));
INVX1 gate2050(.O (g6851), .I (I12424));
INVX1 gate2051(.O (g6355), .I (I11392));
INVX1 gate2052(.O (I11787), .I (g6273));
INVX1 gate2053(.O (I14394), .I (g7536));
INVX1 gate2054(.O (I12753), .I (g6445));
INVX1 gate2055(.O (g8866), .I (I15184));
INVX1 gate2056(.O (g7210), .I (I13144));
INVX1 gate2057(.O (g2644), .I (I6416));
INVX1 gate2058(.O (g3499), .I (g2185));
INVX1 gate2059(.O (I8971), .I (g4464));
INVX1 gate2060(.O (I12145), .I (g5971));
INVX1 gate2061(.O (g1638), .I (g1092));
INVX1 gate2062(.O (I11302), .I (g5796));
INVX1 gate2063(.O (I7738), .I (g3038));
INVX1 gate2064(.O (g5873), .I (g5367));
INVX1 gate2065(.O (I13302), .I (g7164));
INVX1 gate2066(.O (g5037), .I (g4438));
INVX1 gate2067(.O (g9111), .I (I15723));
INVX1 gate2068(.O (I12199), .I (g6475));
INVX1 gate2069(.O (g7013), .I (I12757));
INVX1 gate2070(.O (g9311), .I (I16049));
INVX1 gate2071(.O (g5437), .I (g5041));
INVX1 gate2072(.O (I11827), .I (g6231));
INVX1 gate2073(.O (g5653), .I (g4748));
INVX1 gate2074(.O (g7413), .I (I13524));
INVX1 gate2075(.O (I13743), .I (g7454));
INVX1 gate2076(.O (g3926), .I (I7581));
INVX1 gate2077(.O (g5302), .I (g5028));
INVX1 gate2078(.O (I14420), .I (g7554));
INVX1 gate2079(.O (I15208), .I (g8810));
INVX1 gate2080(.O (g2818), .I (g1792));
INVX1 gate2081(.O (g6063), .I (I10678));
INVX1 gate2082(.O (g4070), .I (I7847));
INVX1 gate2083(.O (I12529), .I (g6628));
INVX1 gate2084(.O (g2867), .I (g2222));
INVX1 gate2085(.O (g3754), .I (g2543));
INVX1 gate2086(.O (I9600), .I (g4698));
INVX1 gate2087(.O (g8198), .I (g7721));
INVX1 gate2088(.O (g8747), .I (g8545));
INVX1 gate2089(.O (g4025), .I (I7792));
INVX1 gate2090(.O (I14318), .I (g7657));
INVX1 gate2091(.O (g5719), .I (I10236));
INVX1 gate2092(.O (I12696), .I (g6503));
INVX1 gate2093(.O (g9374), .I (I16148));
INVX1 gate2094(.O (I14227), .I (g7552));
INVX1 gate2095(.O (I5689), .I (g906));
INVX1 gate2096(.O (I7959), .I (g2793));
INVX1 gate2097(.O (g1758), .I (g1084));
INVX1 gate2098(.O (g1589), .I (g746));
INVX1 gate2099(.O (I14025), .I (g7500));
INVX1 gate2100(.O (I7517), .I (g3578));
INVX1 gate2101(.O (I11803), .I (g6280));
INVX1 gate2102(.O (I7082), .I (g2470));
INVX1 gate2103(.O (g2893), .I (I6615));
INVX1 gate2104(.O (I15726), .I (g9069));
INVX1 gate2105(.O (g7117), .I (I12939));
INVX1 gate2106(.O (g6279), .I (I11132));
INVX1 gate2107(.O (g5917), .I (g5412));
INVX1 gate2108(.O (g7317), .I (I13383));
INVX1 gate2109(.O (I14058), .I (g7544));
INVX1 gate2110(.O (g6720), .I (g6254));
INVX1 gate2111(.O (I5428), .I (g49));
INVX1 gate2112(.O (g6118), .I (g5549));
INVX1 gate2113(.O (g6167), .I (I10862));
INVX1 gate2114(.O (g6318), .I (I11281));
INVX1 gate2115(.O (g1571), .I (g669));
INVX1 gate2116(.O (g3983), .I (g2845));
INVX1 gate2117(.O (g6367), .I (I11428));
INVX1 gate2118(.O (g9180), .I (I15824));
INVX1 gate2119(.O (g6872), .I (I12487));
INVX1 gate2120(.O (g7601), .I (g7450));
INVX1 gate2121(.O (I15607), .I (g8994));
INVX1 gate2122(.O (g9380), .I (g9379));
INVX1 gate2123(.O (g3862), .I (I7389));
INVX1 gate2124(.O (g5042), .I (I9396));
INVX1 gate2125(.O (g1711), .I (I5555));
INVX1 gate2126(.O (g2274), .I (g782));
INVX1 gate2127(.O (g6652), .I (I11936));
INVX1 gate2128(.O (I12161), .I (g5971));
INVX1 gate2129(.O (g4678), .I (I8935));
INVX1 gate2130(.O (g3712), .I (g1952));
INVX1 gate2131(.O (g8524), .I (g7855));
INVX1 gate2132(.O (g6843), .I (I12400));
INVX1 gate2133(.O (I15530), .I (g8972));
INVX1 gate2134(.O (g5786), .I (I10403));
INVX1 gate2135(.O (g4006), .I (I7749));
INVX1 gate2136(.O (g2170), .I (g1229));
INVX1 gate2137(.O (g1827), .I (g762));
INVX1 gate2138(.O (g2614), .I (g1562));
INVX1 gate2139(.O (g9020), .I (I15484));
INVX1 gate2140(.O (g7775), .I (I14196));
INVX1 gate2141(.O (g5164), .I (I9618));
INVX1 gate2142(.O (g6393), .I (I11506));
INVX1 gate2143(.O (g4635), .I (I8820));
INVX1 gate2144(.O (g5364), .I (g5124));
INVX1 gate2145(.O (I15565), .I (g8980));
INVX1 gate2146(.O (g2325), .I (I6118));
INVX1 gate2147(.O (g2821), .I (g1786));
INVX1 gate2148(.O (I12259), .I (g6652));
INVX1 gate2149(.O (I10377), .I (g5188));
INVX1 gate2150(.O (g1774), .I (I5616));
INVX1 gate2151(.O (I12708), .I (g6482));
INVX1 gate2152(.O (g7581), .I (I13888));
INVX1 gate2153(.O (I11662), .I (g5956));
INVX1 gate2154(.O (I10739), .I (g5572));
INVX1 gate2155(.O (g4087), .I (I7882));
INVX1 gate2156(.O (g4105), .I (I7928));
INVX1 gate2157(.O (g8152), .I (I14388));
INVX1 gate2158(.O (I9076), .I (g4353));
INVX1 gate2159(.O (g5054), .I (g4457));
INVX1 gate2160(.O (g6834), .I (I12373));
INVX1 gate2161(.O (g4801), .I (I9126));
INVX1 gate2162(.O (g8867), .I (I15187));
INVX1 gate2163(.O (I9889), .I (g4819));
INVX1 gate2164(.O (I14739), .I (g8173));
INVX1 gate2165(.O (g2939), .I (g2348));
INVX1 gate2166(.O (g3961), .I (g3131));
INVX1 gate2167(.O (g7060), .I (g6654));
INVX1 gate2168(.O (I11890), .I (g6135));
INVX1 gate2169(.O (g1803), .I (g758));
INVX1 gate2170(.O (g7460), .I (g7172));
INVX1 gate2171(.O (I15641), .I (g9017));
INVX1 gate2172(.O (I6160), .I (g324));
INVX1 gate2173(.O (g5725), .I (g4841));
INVX1 gate2174(.O (g4748), .I (g4465));
INVX1 gate2175(.O (I11482), .I (g6117));
INVX1 gate2176(.O (g6598), .I (I11806));
INVX1 gate2177(.O (g3927), .I (I7584));
INVX1 gate2178(.O (I5609), .I (g16));
INVX1 gate2179(.O (I11248), .I (g6149));
INVX1 gate2180(.O (g1780), .I (g614));
INVX1 gate2181(.O (I12244), .I (g6642));
INVX1 gate2182(.O (I11710), .I (g6098));
INVX1 gate2183(.O (I13710), .I (g7340));
INVX1 gate2184(.O (g2636), .I (g1580));
INVX1 gate2185(.O (g7739), .I (I14088));
INVX1 gate2186(.O (g3014), .I (I6767));
INVX1 gate2187(.O (I9651), .I (g4805));
INVX1 gate2188(.O (g6321), .I (I11290));
INVX1 gate2189(.O (g4226), .I (g3591));
INVX1 gate2190(.O (g8386), .I (g8014));
INVX1 gate2191(.O (I5883), .I (g80));
INVX1 gate2192(.O (g2106), .I (I5883));
INVX1 gate2193(.O (g8975), .I (I15429));
INVX1 gate2194(.O (g3946), .I (g3097));
INVX1 gate2195(.O (g2306), .I (I6075));
INVX1 gate2196(.O (I13779), .I (g7406));
INVX1 gate2197(.O (g9204), .I (I15894));
INVX1 gate2198(.O (I15408), .I (g8896));
INVX1 gate2199(.O (I15635), .I (g8976));
INVX1 gate2200(.O (g6625), .I (I11867));
INVX1 gate2201(.O (g1662), .I (g1412));
INVX1 gate2202(.O (g2790), .I (g1793));
INVX1 gate2203(.O (g7937), .I (I14285));
INVX1 gate2204(.O (I7762), .I (g3029));
INVX1 gate2205(.O (I12810), .I (g6607));
INVX1 gate2206(.O (g6232), .I (I11031));
INVX1 gate2207(.O (I11778), .I (g6180));
INVX1 gate2208(.O (g3903), .I (I7498));
INVX1 gate2209(.O (g9100), .I (I15690));
INVX1 gate2210(.O (I12068), .I (g5847));
INVX1 gate2211(.O (I10427), .I (g5210));
INVX1 gate2212(.O (g7479), .I (I13635));
INVX1 gate2213(.O (g9300), .I (I16026));
INVX1 gate2214(.O (g5412), .I (I9850));
INVX1 gate2215(.O (I10366), .I (g5715));
INVX1 gate2216(.O (g6253), .I (g5403));
INVX1 gate2217(.O (g6938), .I (I12635));
INVX1 gate2218(.O (I14427), .I (g7835));
INVX1 gate2219(.O (I5466), .I (g926));
INVX1 gate2220(.O (g6813), .I (I12310));
INVX1 gate2221(.O (g7294), .I (I13314));
INVX1 gate2222(.O (g4373), .I (I8360));
INVX1 gate2223(.O (g3513), .I (g2407));
INVX1 gate2224(.O (I9139), .I (g4364));
INVX1 gate2225(.O (g6909), .I (I12592));
INVX1 gate2226(.O (g7190), .I (I13112));
INVX1 gate2227(.O (g2622), .I (g1568));
INVX1 gate2228(.O (I11945), .I (g5874));
INVX1 gate2229(.O (I12337), .I (g6724));
INVX1 gate2230(.O (I5365), .I (g3843));
INVX1 gate2231(.O (I5861), .I (g1313));
INVX1 gate2232(.O (I11356), .I (g5799));
INVX1 gate2233(.O (I13356), .I (g7221));
INVX1 gate2234(.O (g1816), .I (g767));
INVX1 gate2235(.O (g5171), .I (I9639));
INVX1 gate2236(.O (g4602), .I (I8721));
INVX1 gate2237(.O (g7501), .I (I13679));
INVX1 gate2238(.O (I11380), .I (g5822));
INVX1 gate2239(.O (I10403), .I (g5202));
INVX1 gate2240(.O (g5787), .I (I10406));
INVX1 gate2241(.O (g4007), .I (I7752));
INVX1 gate2242(.O (g2904), .I (g2287));
INVX1 gate2243(.O (I14403), .I (g7679));
INVX1 gate2244(.O (g7156), .I (I13042));
INVX1 gate2245(.O (g5956), .I (I10582));
INVX1 gate2246(.O (g6552), .I (I11722));
INVX1 gate2247(.O (g7356), .I (I13484));
INVX1 gate2248(.O (g4920), .I (g4105));
INVX1 gate2249(.O (g6606), .I (I11824));
INVX1 gate2250(.O (g4578), .I (g2917));
INVX1 gate2251(.O (I11090), .I (g1000));
INVX1 gate2252(.O (I7928), .I (g2873));
INVX1 gate2253(.O (I11998), .I (g5918));
INVX1 gate2254(.O (g8544), .I (I14657));
INVX1 gate2255(.O (g3831), .I (I7296));
INVX1 gate2256(.O (I11233), .I (g6147));
INVX1 gate2257(.O (g2514), .I (g1330));
INVX1 gate2258(.O (g4718), .I (I9018));
INVX1 gate2259(.O (g8483), .I (g8038));
INVX1 gate2260(.O (I8962), .I (g4553));
INVX1 gate2261(.O (I7064), .I (g2458));
INVX1 gate2262(.O (I11672), .I (g5971));
INVX1 gate2263(.O (g1847), .I (g765));
INVX1 gate2264(.O (I9672), .I (g4803));
INVX1 gate2265(.O (I15711), .I (g9075));
INVX1 gate2266(.O (I13672), .I (g7242));
INVX1 gate2267(.O (I7899), .I (g3743));
INVX1 gate2268(.O (g4535), .I (g2876));
INVX1 gate2269(.O (g2403), .I (g1176));
INVX1 gate2270(.O (g8636), .I (I14718));
INVX1 gate2271(.O (g1685), .I (I5528));
INVX1 gate2272(.O (g2145), .I (g1296));
INVX1 gate2273(.O (g6687), .I (I12003));
INVX1 gate2274(.O (g2345), .I (I6151));
INVX1 gate2275(.O (g2841), .I (g2208));
INVX1 gate2276(.O (I7785), .I (g3029));
INVX1 gate2277(.O (g7704), .I (I14001));
INVX1 gate2278(.O (g4582), .I (g2922));
INVX1 gate2279(.O (g3805), .I (g1752));
INVX1 gate2280(.O (g3916), .I (I7545));
INVX1 gate2281(.O (g9323), .I (g9315));
INVX1 gate2282(.O (g6586), .I (I11778));
INVX1 gate2283(.O (g8790), .I (g8585));
INVX1 gate2284(.O (g2695), .I (g1672));
INVX1 gate2285(.O (g4015), .I (g3160));
INVX1 gate2286(.O (g2637), .I (g1581));
INVX1 gate2287(.O (I11449), .I (g6068));
INVX1 gate2288(.O (I12918), .I (g7013));
INVX1 gate2289(.O (g5684), .I (I10183));
INVX1 gate2290(.O (g8061), .I (I14330));
INVX1 gate2291(.O (g5745), .I (I10292));
INVX1 gate2292(.O (I15492), .I (g8971));
INVX1 gate2293(.O (g5639), .I (g4748));
INVX1 gate2294(.O (I14127), .I (g7594));
INVX1 gate2295(.O (g7163), .I (I13063));
INVX1 gate2296(.O (g3947), .I (I7640));
INVX1 gate2297(.O (I11897), .I (g6141));
INVX1 gate2298(.O (g2307), .I (I6078));
INVX1 gate2299(.O (I11961), .I (g5988));
INVX1 gate2300(.O (g7032), .I (g6525));
INVX1 gate2301(.O (g2536), .I (g1354));
INVX1 gate2302(.O (g5109), .I (I9493));
INVX1 gate2303(.O (I13897), .I (g7354));
INVX1 gate2304(.O (g8756), .I (g8564));
INVX1 gate2305(.O (g3798), .I (g1757));
INVX1 gate2306(.O (g5309), .I (g4969));
INVX1 gate2307(.O (g7432), .I (I13559));
INVX1 gate2308(.O (g6141), .I (I10786));
INVX1 gate2309(.O (g6860), .I (I12451));
INVX1 gate2310(.O (g2359), .I (g1397));
INVX1 gate2311(.O (g4664), .I (I8907));
INVX1 gate2312(.O (I9499), .I (g4382));
INVX1 gate2313(.O (g6341), .I (I11350));
INVX1 gate2314(.O (I11404), .I (g5834));
INVX1 gate2315(.O (g3560), .I (g2361));
INVX1 gate2316(.O (g9351), .I (I16103));
INVX1 gate2317(.O (g2223), .I (I5942));
INVX1 gate2318(.O (I7844), .I (g3784));
INVX1 gate2319(.O (I15982), .I (g9236));
INVX1 gate2320(.O (g5808), .I (I10457));
INVX1 gate2321(.O (g1562), .I (g636));
INVX1 gate2322(.O (I6680), .I (g1558));
INVX1 gate2323(.O (g6645), .I (I11917));
INVX1 gate2324(.O (I16040), .I (g9285));
INVX1 gate2325(.O (g4721), .I (I9025));
INVX1 gate2326(.O (I14103), .I (g7584));
INVX1 gate2327(.O (I11212), .I (g6146));
INVX1 gate2328(.O (g2016), .I (I5852));
INVX1 gate2329(.O (I7731), .I (g3029));
INVX1 gate2330(.O (g5759), .I (I10350));
INVX1 gate2331(.O (g8514), .I (g8040));
INVX1 gate2332(.O (g3873), .I (g2956));
INVX1 gate2333(.O (g3632), .I (I7101));
INVX1 gate2334(.O (g3095), .I (I6831));
INVX1 gate2335(.O (g1817), .I (I5689));
INVX1 gate2336(.O (g3495), .I (g1616));
INVX1 gate2337(.O (g3653), .I (g2459));
INVX1 gate2338(.O (I8180), .I (g3529));
INVX1 gate2339(.O (I12322), .I (g6751));
INVX1 gate2340(.O (g8145), .I (I14381));
INVX1 gate2341(.O (g2522), .I (g1342));
INVX1 gate2342(.O (I14181), .I (g7725));
INVX1 gate2343(.O (g7157), .I (I13045));
INVX1 gate2344(.O (g2642), .I (g1588));
INVX1 gate2345(.O (I8832), .I (g3936));
INVX1 gate2346(.O (g6879), .I (I12508));
INVX1 gate2347(.O (g7357), .I (I13487));
INVX1 gate2348(.O (g6607), .I (I11827));
INVX1 gate2349(.O (I12532), .I (g6594));
INVX1 gate2350(.O (g3579), .I (g1929));
INVX1 gate2351(.O (g3869), .I (I7400));
INVX1 gate2352(.O (g6962), .I (I12687));
INVX1 gate2353(.O (I8853), .I (g4034));
INVX1 gate2354(.O (g6659), .I (I11955));
INVX1 gate2355(.O (I12158), .I (g5956));
INVX1 gate2356(.O (g6358), .I (I11401));
INVX1 gate2357(.O (g6506), .I (I11680));
INVX1 gate2358(.O (g1751), .I (g452));
INVX1 gate2359(.O (I5847), .I (g1360));
INVX1 gate2360(.O (I12561), .I (g6449));
INVX1 gate2361(.O (I16183), .I (g9388));
INVX1 gate2362(.O (g5604), .I (g4969));
INVX1 gate2363(.O (I12295), .I (g6693));
INVX1 gate2364(.O (g3917), .I (I7548));
INVX1 gate2365(.O (g2654), .I (I6446));
INVX1 gate2366(.O (I10190), .I (g4670));
INVX1 gate2367(.O (g1585), .I (g724));
INVX1 gate2368(.O (g4689), .I (I8966));
INVX1 gate2369(.O (g6587), .I (I11781));
INVX1 gate2370(.O (g9372), .I (I16142));
INVX1 gate2371(.O (I15522), .I (g9018));
INVX1 gate2372(.O (I15663), .I (g9066));
INVX1 gate2373(.O (I14190), .I (g7531));
INVX1 gate2374(.O (I9543), .I (g4279));
INVX1 gate2375(.O (g6111), .I (g5453));
INVX1 gate2376(.O (g8223), .I (I14448));
INVX1 gate2377(.O (g6311), .I (I11260));
INVX1 gate2378(.O (g5833), .I (I10522));
INVX1 gate2379(.O (I7814), .I (g2605));
INVX1 gate2380(.O (I13646), .I (g7245));
INVX1 gate2381(.O (g9235), .I (I15959));
INVX1 gate2382(.O (g4028), .I (I7797));
INVX1 gate2383(.O (g2880), .I (g2234));
INVX1 gate2384(.O (I7350), .I (g2971));
INVX1 gate2385(.O (I6574), .I (g576));
INVX1 gate2386(.O (g2595), .I (g1643));
INVX1 gate2387(.O (I6864), .I (g2528));
INVX1 gate2388(.O (I11971), .I (g6179));
INVX1 gate2389(.O (g4030), .I (g3160));
INVX1 gate2390(.O (g8016), .I (I14311));
INVX1 gate2391(.O (g8757), .I (g8585));
INVX1 gate2392(.O (g5584), .I (g4841));
INVX1 gate2393(.O (g1673), .I (g1504));
INVX1 gate2394(.O (g6374), .I (I11449));
INVX1 gate2395(.O (I14211), .I (g7712));
INVX1 gate2396(.O (g9134), .I (I15776));
INVX1 gate2397(.O (I15553), .I (g9009));
INVX1 gate2398(.O (I13369), .I (g7268));
INVX1 gate2399(.O (g2272), .I (I6021));
INVX1 gate2400(.O (I14088), .I (g7585));
INVX1 gate2401(.O (g4564), .I (I8665));
INVX1 gate2402(.O (I11368), .I (g5833));
INVX1 gate2403(.O (g8642), .I (I14732));
INVX1 gate2404(.O (I5562), .I (g1300));
INVX1 gate2405(.O (I12364), .I (g6714));
INVX1 gate2406(.O (I7769), .I (g3038));
INVX1 gate2407(.O (g5162), .I (I9612));
INVX1 gate2408(.O (g3770), .I (g2551));
INVX1 gate2409(.O (g5268), .I (I9788));
INVX1 gate2410(.O (I9014), .I (g3864));
INVX1 gate2411(.O (g5362), .I (I9823));
INVX1 gate2412(.O (I10497), .I (g5233));
INVX1 gate2413(.O (I15536), .I (g9004));
INVX1 gate2414(.O (g1772), .I (g607));
INVX1 gate2415(.O (g6380), .I (I11467));
INVX1 gate2416(.O (I9660), .I (g4806));
INVX1 gate2417(.O (g6591), .I (I11787));
INVX1 gate2418(.O (I15702), .I (g9064));
INVX1 gate2419(.O (I13850), .I (g7328));
INVX1 gate2420(.O (g6832), .I (I12367));
INVX1 gate2421(.O (I5817), .I (g1081));
INVX1 gate2422(.O (g2982), .I (g1848));
INVX1 gate2423(.O (g8874), .I (I15208));
INVX1 gate2424(.O (g3532), .I (g2407));
INVX1 gate2425(.O (I7967), .I (g2787));
INVX1 gate2426(.O (g7778), .I (I14205));
INVX1 gate2427(.O (g1743), .I (g598));
INVX1 gate2428(.O (g2234), .I (I5963));
INVX1 gate2429(.O (g6853), .I (I12430));
INVX1 gate2430(.O (g2128), .I (g1284));
INVX1 gate2431(.O (g4638), .I (I8829));
INVX1 gate2432(.O (g2629), .I (g1574));
INVX1 gate2433(.O (g6020), .I (g5367));
INVX1 gate2434(.O (g2328), .I (I6127));
INVX1 gate2435(.O (I10987), .I (g5609));
INVX1 gate2436(.O (I12289), .I (g6702));
INVX1 gate2437(.O (I5605), .I (g58));
INVX1 gate2438(.O (I10250), .I (g5268));
INVX1 gate2439(.O (g7735), .I (I14076));
INVX1 gate2440(.O (g4609), .I (I8742));
INVX1 gate2441(.O (g6507), .I (I11683));
INVX1 gate2442(.O (g4308), .I (I8277));
INVX1 gate2443(.O (g1011), .I (I5413));
INVX1 gate2444(.O (I13228), .I (g6892));
INVX1 gate2445(.O (g9113), .I (I15729));
INVX1 gate2446(.O (g6794), .I (I12253));
INVX1 gate2447(.O (g1856), .I (g774));
INVX1 gate2448(.O (I12571), .I (g6729));
INVX1 gate2449(.O (g9313), .I (I16055));
INVX1 gate2450(.O (I11011), .I (g5693));
INVX1 gate2451(.O (I5751), .I (g963));
INVX1 gate2452(.O (g5086), .I (I9460));
INVX1 gate2453(.O (g8880), .I (I15218));
INVX1 gate2454(.O (g3189), .I (I6864));
INVX1 gate2455(.O (I13716), .I (g7331));
INVX1 gate2456(.O (g5730), .I (I10247));
INVX1 gate2457(.O (g7475), .I (I13631));
INVX1 gate2458(.O (I16072), .I (g9303));
INVX1 gate2459(.O (g3990), .I (g3160));
INVX1 gate2460(.O (g2554), .I (I6376));
INVX1 gate2461(.O (I14338), .I (g7581));
INVX1 gate2462(.O (g5185), .I (I9681));
INVX1 gate2463(.O (g4589), .I (g2930));
INVX1 gate2464(.O (I10969), .I (g5606));
INVX1 gate2465(.O (g9094), .I (I15672));
INVX1 gate2466(.O (g7627), .I (I13956));
INVX1 gate2467(.O (g3888), .I (g3097));
INVX1 gate2468(.O (I15062), .I (g8632));
INVX1 gate2469(.O (g6905), .I (I12586));
INVX1 gate2470(.O (g3029), .I (g1929));
INVX1 gate2471(.O (g7292), .I (I13308));
INVX1 gate2472(.O (g3787), .I (g1842));
INVX1 gate2473(.O (g8017), .I (g7692));
INVX1 gate2474(.O (g6628), .I (I11880));
INVX1 gate2475(.O (I15933), .I (g9210));
INVX1 gate2476(.O (g7526), .I (I13758));
INVX1 gate2477(.O (g5470), .I (g4899));
INVX1 gate2478(.O (g5897), .I (I10569));
INVX1 gate2479(.O (g3956), .I (g2845));
INVX1 gate2480(.O (g5025), .I (I9363));
INVX1 gate2481(.O (g6515), .I (g6125));
INVX1 gate2482(.O (I11627), .I (g5874));
INVX1 gate2483(.O (g6630), .I (I11884));
INVX1 gate2484(.O (g4571), .I (g2908));
INVX1 gate2485(.O (I12687), .I (g6745));
INVX1 gate2486(.O (g3675), .I (I7167));
INVX1 gate2487(.O (I12976), .I (g6928));
INVX1 gate2488(.O (g1573), .I (g677));
INVX1 gate2489(.O (g1863), .I (g68));
INVX1 gate2490(.O (g6300), .I (I11227));
INVX1 gate2491(.O (I13112), .I (g7021));
INVX1 gate2492(.O (g7603), .I (I13940));
INVX1 gate2493(.O (I11050), .I (g5335));
INVX1 gate2494(.O (I11958), .I (g5874));
INVX1 gate2495(.O (g7039), .I (g6543));
INVX1 gate2496(.O (I9422), .I (g4360));
INVX1 gate2497(.O (I8351), .I (g1160));
INVX1 gate2498(.O (g8234), .I (I14489));
INVX1 gate2499(.O (g4455), .I (g3811));
INVX1 gate2500(.O (g2902), .I (g2285));
INVX1 gate2501(.O (g7439), .I (I13574));
INVX1 gate2502(.O (I12643), .I (g6501));
INVX1 gate2503(.O (I5368), .I (g3853));
INVX1 gate2504(.O (I11386), .I (g5764));
INVX1 gate2505(.O (g1569), .I (g661));
INVX1 gate2506(.O (g453), .I (I5362));
INVX1 gate2507(.O (I5772), .I (g1240));
INVX1 gate2508(.O (g2490), .I (I6326));
INVX1 gate2509(.O (I6024), .I (g544));
INVX1 gate2510(.O (I5531), .I (g866));
INVX1 gate2511(.O (g2366), .I (I6198));
INVX1 gate2512(.O (I12669), .I (g6477));
INVX1 gate2513(.O (g7583), .I (I13894));
INVX1 gate2514(.O (g7702), .I (I13997));
INVX1 gate2515(.O (g4196), .I (I8097));
INVX1 gate2516(.O (g5678), .I (I10169));
INVX1 gate2517(.O (I6795), .I (g1683));
INVX1 gate2518(.O (I10503), .I (g5235));
INVX1 gate2519(.O (g3684), .I (g2180));
INVX1 gate2520(.O (g3639), .I (g2424));
INVX1 gate2521(.O (g4803), .I (I9132));
INVX1 gate2522(.O (g6973), .I (I12708));
INVX1 gate2523(.O (g5006), .I (I9333));
INVX1 gate2524(.O (g3338), .I (g1901));
INVX1 gate2525(.O (g8800), .I (I15010));
INVX1 gate2526(.O (g3963), .I (I7672));
INVX1 gate2527(.O (g9360), .I (I16116));
INVX1 gate2528(.O (I15574), .I (g8983));
INVX1 gate2529(.O (g4538), .I (g2880));
INVX1 gate2530(.O (g1688), .I (I5535));
INVX1 gate2531(.O (g2148), .I (g1304));
INVX1 gate2532(.O (I15205), .I (g8809));
INVX1 gate2533(.O (g2649), .I (I6431));
INVX1 gate2534(.O (g4780), .I (I9089));
INVX1 gate2535(.O (g1857), .I (g889));
INVX1 gate2536(.O (g2348), .I (I6160));
INVX1 gate2537(.O (I7788), .I (g2595));
INVX1 gate2538(.O (g9050), .I (I15550));
INVX1 gate2539(.O (g5682), .I (I10177));
INVX1 gate2540(.O (g5766), .I (I10373));
INVX1 gate2541(.O (g5087), .I (I9463));
INVX1 gate2542(.O (g1976), .I (g1269));
INVX1 gate2543(.O (g6969), .I (I12702));
INVX1 gate2544(.O (I15912), .I (g9193));
INVX1 gate2545(.O (I9095), .I (g4283));
INVX1 gate2546(.O (g5801), .I (I10442));
INVX1 gate2547(.O (g3808), .I (g1827));
INVX1 gate2548(.O (g7276), .I (I13264));
INVX1 gate2549(.O (g5487), .I (I9907));
INVX1 gate2550(.O (I14315), .I (g7676));
INVX1 gate2551(.O (I6643), .I (g1970));
INVX1 gate2552(.O (I11793), .I (g6188));
INVX1 gate2553(.O (I11428), .I (g5813));
INVX1 gate2554(.O (I12424), .I (g6446));
INVX1 gate2555(.O (I13428), .I (g7167));
INVX1 gate2556(.O (g3707), .I (g2226));
INVX1 gate2557(.O (g6323), .I (I11296));
INVX1 gate2558(.O (I14819), .I (g8647));
INVX1 gate2559(.O (g4662), .I (I8901));
INVX1 gate2560(.O (g2698), .I (g1673));
INVX1 gate2561(.O (g4018), .I (I7775));
INVX1 gate2562(.O (I12558), .I (g6449));
INVX1 gate2563(.O (I14202), .I (g7708));
INVX1 gate2564(.O (I8172), .I (g3524));
INVX1 gate2565(.O (I14257), .I (g7716));
INVX1 gate2566(.O (I9579), .I (g4713));
INVX1 gate2567(.O (g2964), .I (I6716));
INVX1 gate2568(.O (I14055), .I (g7495));
INVX1 gate2569(.O (I16020), .I (g9264));
INVX1 gate2570(.O (g9379), .I (I16161));
INVX1 gate2571(.O (I7392), .I (g3230));
INVX1 gate2572(.O (g5755), .I (g5494));
INVX1 gate2573(.O (I15592), .I (g8989));
INVX1 gate2574(.O (I15756), .I (g9081));
INVX1 gate2575(.O (g7527), .I (I13761));
INVX1 gate2576(.O (I14070), .I (g7714));
INVX1 gate2577(.O (g3957), .I (I7662));
INVX1 gate2578(.O (I12544), .I (g6617));
INVX1 gate2579(.O (I6099), .I (g584));
INVX1 gate2580(.O (I9752), .I (g4705));
INVX1 gate2581(.O (g4093), .I (I7902));
INVX1 gate2582(.O (g8512), .I (g8094));
INVX1 gate2583(.O (I8282), .I (g3515));
INVX1 gate2584(.O (I16046), .I (g9288));
INVX1 gate2585(.O (g1760), .I (I5605));
INVX1 gate2586(.O (g4493), .I (I8543));
INVX1 gate2587(.O (g7764), .I (I14163));
INVX1 gate2588(.O (g6351), .I (I11380));
INVX1 gate2589(.O (g6648), .I (I11926));
INVX1 gate2590(.O (g6875), .I (I12496));
INVX1 gate2591(.O (g7546), .I (I13822));
INVX1 gate2592(.O (g3865), .I (g2944));
INVX1 gate2593(.O (I10384), .I (g5193));
INVX1 gate2594(.O (g6655), .I (I11945));
INVX1 gate2595(.O (g5445), .I (g5059));
INVX1 gate2596(.O (g5173), .I (I9645));
INVX1 gate2597(.O (I11317), .I (g5787));
INVX1 gate2598(.O (g3604), .I (g2407));
INVX1 gate2599(.O (I13317), .I (g7211));
INVX1 gate2600(.O (g5491), .I (g4918));
INVX1 gate2601(.O (g3498), .I (g1616));
INVX1 gate2602(.O (I14067), .I (g7550));
INVX1 gate2603(.O (I14094), .I (g7593));
INVX1 gate2604(.O (g4381), .I (g3466));
INVX1 gate2605(.O (g8649), .I (I14743));
INVX1 gate2606(.O (g6010), .I (I10608));
INVX1 gate2607(.O (g3833), .I (I7302));
INVX1 gate2608(.O (I11129), .I (g5418));
INVX1 gate2609(.O (g2872), .I (I6590));
INVX1 gate2610(.O (g1924), .I (g174));
INVX1 gate2611(.O (g5169), .I (I9633));
INVX1 gate2612(.O (g4685), .I (I8952));
INVX1 gate2613(.O (g4197), .I (g3591));
INVX1 gate2614(.O (I10801), .I (g5463));
INVX1 gate2615(.O (g6410), .I (I11533));
INVX1 gate2616(.O (g7224), .I (I13164));
INVX1 gate2617(.O (I7520), .I (g2734));
INVX1 gate2618(.O (g4021), .I (g3131));
INVX1 gate2619(.O (g5007), .I (I9336));
INVX1 gate2620(.O (I13057), .I (g6968));
INVX1 gate2621(.O (I14801), .I (g8608));
INVX1 gate2622(.O (g2652), .I (I6440));
INVX1 gate2623(.O (g1779), .I (g612));
INVX1 gate2624(.O (g2057), .I (I5868));
INVX1 gate2625(.O (I7640), .I (g3062));
INVX1 gate2626(.O (I12124), .I (g5847));
INVX1 gate2627(.O (I12678), .I (g6516));
INVX1 gate2628(.O (g6884), .I (I12523));
INVX1 gate2629(.O (g2843), .I (I6571));
INVX1 gate2630(.O (g7120), .I (I12948));
INVX1 gate2631(.O (g5059), .I (I9419));
INVX1 gate2632(.O (g6839), .I (I12388));
INVX1 gate2633(.O (g2457), .I (g24));
INVX1 gate2634(.O (g5578), .I (g4841));
INVX1 gate2635(.O (g5868), .I (I10555));
INVX1 gate2636(.O (g7320), .I (I13388));
INVX1 gate2637(.O (g2989), .I (g1843));
INVX1 gate2638(.O (g3539), .I (g2424));
INVX1 gate2639(.O (g3896), .I (I7473));
INVX1 gate2640(.O (I11245), .I (g6143));
INVX1 gate2641(.O (g5459), .I (g4882));
INVX1 gate2642(.O (I14019), .I (g7480));
INVX1 gate2643(.O (g2393), .I (I6267));
INVX1 gate2644(.O (g5718), .I (g4841));
INVX1 gate2645(.O (I12460), .I (g6674));
INVX1 gate2646(.O (I12939), .I (g7022));
INVX1 gate2647(.O (I11323), .I (g5808));
INVX1 gate2648(.O (g1977), .I (g1357));
INVX1 gate2649(.O (I11299), .I (g5786));
INVX1 gate2650(.O (I13323), .I (g7145));
INVX1 gate2651(.O (I14196), .I (g7534));
INVX1 gate2652(.O (I13299), .I (g7163));
INVX1 gate2653(.O (I14695), .I (g8016));
INVX1 gate2654(.O (g7277), .I (I13267));
INVX1 gate2655(.O (g1588), .I (g741));
INVX1 gate2656(.O (I11533), .I (g5847));
INVX1 gate2657(.O (g2834), .I (I6564));
INVX1 gate2658(.O (g2971), .I (I6723));
INVX1 gate2659(.O (I13533), .I (g7220));
INVX1 gate2660(.O (g8063), .I (I14334));
INVX1 gate2661(.O (g5582), .I (g4969));
INVX1 gate2662(.O (I15405), .I (g8902));
INVX1 gate2663(.O (g6278), .I (I11129));
INVX1 gate2664(.O (g8463), .I (g8094));
INVX1 gate2665(.O (g2686), .I (g1667));
INVX1 gate2666(.O (g6372), .I (I11443));
INVX1 gate2667(.O (g7789), .I (I14224));
INVX1 gate2668(.O (g5261), .I (g4748));
INVX1 gate2669(.O (g3019), .I (g2007));
INVX1 gate2670(.O (g9132), .I (I15770));
INVX1 gate2671(.O (g5793), .I (I10418));
INVX1 gate2672(.O (I12065), .I (g5897));
INVX1 gate2673(.O (I8202), .I (g3560));
INVX1 gate2674(.O (g9332), .I (g9322));
INVX1 gate2675(.O (g6618), .I (g6003));
INVX1 gate2676(.O (g1665), .I (g1467));
INVX1 gate2677(.O (g6143), .I (I10796));
INVX1 gate2678(.O (g7516), .I (I13728));
INVX1 gate2679(.O (I7765), .I (g2595));
INVX1 gate2680(.O (g6343), .I (I11356));
INVX1 gate2681(.O (g4562), .I (g3466));
INVX1 gate2682(.O (g6235), .I (I11034));
INVX1 gate2683(.O (g5015), .I (I9347));
INVX1 gate2684(.O (g3052), .I (g2096));
INVX1 gate2685(.O (g9209), .I (g9199));
INVX1 gate2686(.O (g9353), .I (I16107));
INVX1 gate2687(.O (I7911), .I (g2767));
INVX1 gate2688(.O (I10457), .I (g5218));
INVX1 gate2689(.O (I8094), .I (g2976));
INVX1 gate2690(.O (g7771), .I (I14184));
INVX1 gate2691(.O (I14457), .I (g8093));
INVX1 gate2692(.O (g6566), .I (I11740));
INVX1 gate2693(.O (g4631), .I (I8808));
INVX1 gate2694(.O (I13737), .I (g7446));
INVX1 gate2695(.O (g372), .I (I5359));
INVX1 gate2696(.O (I15583), .I (g8986));
INVX1 gate2697(.O (g7299), .I (I13329));
INVX1 gate2698(.O (g4257), .I (I8190));
INVX1 gate2699(.O (g6693), .I (I12011));
INVX1 gate2700(.O (g6134), .I (g5428));
INVX1 gate2701(.O (g8619), .I (I14695));
INVX1 gate2702(.O (g7547), .I (I13825));
INVX1 gate2703(.O (g6334), .I (I11329));
INVX1 gate2704(.O (g4301), .I (I8264));
INVX1 gate2705(.O (g5246), .I (I9760));
INVX1 gate2706(.O (g2625), .I (g1570));
INVX1 gate2707(.O (g8872), .I (I15202));
INVX1 gate2708(.O (g2232), .I (I5957));
INVX1 gate2709(.O (g4605), .I (I8730));
INVX1 gate2710(.O (g3086), .I (g1852));
INVX1 gate2711(.O (g2253), .I (g1323));
INVX1 gate2712(.O (g2938), .I (g2347));
INVX1 gate2713(.O (g3728), .I (g2202));
INVX1 gate2714(.O (I14001), .I (g7433));
INVX1 gate2715(.O (I13261), .I (g7041));
INVX1 gate2716(.O (I11880), .I (g5748));
INVX1 gate2717(.O (g6555), .I (I11729));
INVX1 gate2718(.O (g6804), .I (I12283));
INVX1 gate2719(.O (I7473), .I (g3546));
INVX1 gate2720(.O (g2909), .I (g2291));
INVX1 gate2721(.O (I6946), .I (g1887));
INVX1 gate2722(.O (I10256), .I (g5401));
INVX1 gate2723(.O (g6792), .I (I12247));
INVX1 gate2724(.O (I11512), .I (g5874));
INVX1 gate2725(.O (g1732), .I (g1439));
INVX1 gate2726(.O (I9675), .I (g4807));
INVX1 gate2727(.O (I13512), .I (g7138));
INVX1 gate2728(.O (g3881), .I (g2969));
INVX1 gate2729(.O (I5383), .I (g647));
INVX1 gate2730(.O (I10280), .I (g5488));
INVX1 gate2731(.O (g8971), .I (I15417));
INVX1 gate2732(.O (g7738), .I (I14085));
INVX1 gate2733(.O (g4585), .I (g2925));
INVX1 gate2734(.O (I8264), .I (g3653));
INVX1 gate2735(.O (g6621), .I (I11855));
INVX1 gate2736(.O (g1944), .I (I5817));
INVX1 gate2737(.O (g3897), .I (g3131));
INVX1 gate2738(.O (g4041), .I (g2605));
INVX1 gate2739(.O (I12915), .I (g7000));
INVX1 gate2740(.O (g9092), .I (I15666));
INVX1 gate2741(.O (I8360), .I (g1186));
INVX1 gate2742(.O (g6313), .I (I11266));
INVX1 gate2743(.O (g7078), .I (g6683));
INVX1 gate2744(.O (g7340), .I (I13438));
INVX1 gate2745(.O (I7377), .I (g3189));
INVX1 gate2746(.O (I10157), .I (g5109));
INVX1 gate2747(.O (I13831), .I (g7322));
INVX1 gate2748(.O (I6036), .I (g130));
INVX1 gate2749(.O (I14157), .I (g7547));
INVX1 gate2750(.O (I12277), .I (g6681));
INVX1 gate2751(.O (I6178), .I (g1220));
INVX1 gate2752(.O (g4673), .I (I8928));
INVX1 gate2753(.O (g6202), .I (I10949));
INVX1 gate2754(.O (g8670), .I (I14804));
INVX1 gate2755(.O (I9684), .I (g4813));
INVX1 gate2756(.O (g7035), .I (g6543));
INVX1 gate2757(.O (I13499), .I (g7134));
INVX1 gate2758(.O (I15803), .I (g9148));
INVX1 gate2759(.O (I9639), .I (g4685));
INVX1 gate2760(.O (g7517), .I (I13731));
INVX1 gate2761(.O (I7287), .I (g2561));
INVX1 gate2762(.O (g6094), .I (I10716));
INVX1 gate2763(.O (I14231), .I (g7566));
INVX1 gate2764(.O (I9791), .I (g4779));
INVX1 gate2765(.O (I6831), .I (g2185));
INVX1 gate2766(.O (g5028), .I (I9372));
INVX1 gate2767(.O (g4669), .I (I8922));
INVX1 gate2768(.O (g1565), .I (g649));
INVX1 gate2769(.O (I8724), .I (g3927));
INVX1 gate2770(.O (g5671), .I (I10160));
INVX1 gate2771(.O (I11722), .I (g5772));
INVX1 gate2772(.O (I12782), .I (g6463));
INVX1 gate2773(.O (I13722), .I (g7442));
INVX1 gate2774(.O (I16090), .I (g9336));
INVX1 gate2775(.O (I6805), .I (g1603));
INVX1 gate2776(.O (g3635), .I (g1949));
INVX1 gate2777(.O (I13924), .I (g7365));
INVX1 gate2778(.O (I5633), .I (g891));
INVX1 gate2779(.O (g1681), .I (g929));
INVX1 gate2780(.O (g6776), .I (I12199));
INVX1 gate2781(.O (I7781), .I (g2605));
INVX1 gate2782(.O (I6422), .I (g1805));
INVX1 gate2783(.O (g6593), .I (I11793));
INVX1 gate2784(.O (g4890), .I (g4075));
INVX1 gate2785(.O (I12352), .I (g6752));
INVX1 gate2786(.O (I13432), .I (g7280));
INVX1 gate2787(.O (g2525), .I (I6354));
INVX1 gate2788(.O (g3801), .I (I7262));
INVX1 gate2789(.O (I14763), .I (g7834));
INVX1 gate2790(.O (I13271), .I (g7067));
INVX1 gate2791(.O (g2645), .I (I6419));
INVX1 gate2792(.O (I8835), .I (g3954));
INVX1 gate2793(.O (g5826), .I (I10503));
INVX1 gate2794(.O (I12418), .I (g6572));
INVX1 gate2795(.O (I7797), .I (g3019));
INVX1 gate2796(.O (g8606), .I (I14683));
INVX1 gate2797(.O (I12170), .I (g5956));
INVX1 gate2798(.O (g4011), .I (I7762));
INVX1 gate2799(.O (I11461), .I (g6094));
INVX1 gate2800(.O (g9076), .I (I15622));
INVX1 gate2801(.O (g5741), .I (I10280));
INVX1 gate2802(.O (g7110), .I (I12918));
INVX1 gate2803(.O (I5732), .I (g859));
INVX1 gate2804(.O (g6264), .I (g5403));
INVX1 gate2805(.O (g7310), .I (I13362));
INVX1 gate2806(.O (I11031), .I (g5335));
INVX1 gate2807(.O (I13031), .I (g6984));
INVX1 gate2808(.O (g5638), .I (g4748));
INVX1 gate2809(.O (g6360), .I (I11407));
INVX1 gate2810(.O (g2879), .I (I6597));
INVX1 gate2811(.O (I13199), .I (g7025));
INVX1 gate2812(.O (I11736), .I (g6076));
INVX1 gate2813(.O (I11887), .I (g5918));
INVX1 gate2814(.O (g9375), .I (I16151));
INVX1 gate2815(.O (I7344), .I (g2964));
INVX1 gate2816(.O (g2962), .I (g2382));
INVX1 gate2817(.O (g5609), .I (g4748));
INVX1 gate2818(.O (I15003), .I (g8633));
INVX1 gate2819(.O (I8799), .I (g3951));
INVX1 gate2820(.O (g2659), .I (g1655));
INVX1 gate2821(.O (g6050), .I (g5246));
INVX1 gate2822(.O (I12167), .I (g5939));
INVX1 gate2823(.O (g2506), .I (I6341));
INVX1 gate2824(.O (g1820), .I (g621));
INVX1 gate2825(.O (I6437), .I (g1784));
INVX1 gate2826(.O (I11696), .I (g5971));
INVX1 gate2827(.O (g7236), .I (g6944));
INVX1 gate2828(.O (I6302), .I (g1313));
INVX1 gate2829(.O (g3091), .I (g1603));
INVX1 gate2830(.O (I13843), .I (g7326));
INVX1 gate2831(.O (I16026), .I (g9267));
INVX1 gate2832(.O (g7762), .I (I14157));
INVX1 gate2833(.O (g3491), .I (g1800));
INVX1 gate2834(.O (g4080), .I (I7867));
INVX1 gate2835(.O (I14076), .I (g7577));
INVX1 gate2836(.O (I14085), .I (g7583));
INVX1 gate2837(.O (g4573), .I (g2911));
INVX1 gate2838(.O (I11764), .I (g6056));
INVX1 gate2839(.O (g5758), .I (I10347));
INVX1 gate2840(.O (I13764), .I (g7479));
INVX1 gate2841(.O (g6724), .I (I12088));
INVX1 gate2842(.O (I11365), .I (g5826));
INVX1 gate2843(.O (g2275), .I (g990));
INVX1 gate2844(.O (g2311), .I (I6090));
INVX1 gate2845(.O (I9539), .I (g4018));
INVX1 gate2846(.O (g6179), .I (I10896));
INVX1 gate2847(.O (I13365), .I (g7267));
INVX1 gate2848(.O (g5466), .I (g4890));
INVX1 gate2849(.O (g4713), .I (I9014));
INVX1 gate2850(.O (I10243), .I (g5026));
INVX1 gate2851(.O (g6379), .I (I11464));
INVX1 gate2852(.O (I11132), .I (g5624));
INVX1 gate2853(.O (g7590), .I (I13915));
INVX1 gate2854(.O (g9184), .I (I15830));
INVX1 gate2855(.O (I13869), .I (g7338));
INVX1 gate2856(.O (I5565), .I (g1296));
INVX1 gate2857(.O (g2615), .I (g1563));
INVX1 gate2858(.O (g6878), .I (I12505));
INVX1 gate2859(.O (g5165), .I (I9621));
INVX1 gate2860(.O (g4569), .I (g2906));
INVX1 gate2861(.O (g5571), .I (I10032));
INVX1 gate2862(.O (g3920), .I (g3097));
INVX1 gate2863(.O (I12022), .I (g5874));
INVX1 gate2864(.O (g3578), .I (I7053));
INVX1 gate2865(.O (g3868), .I (g2948));
INVX1 gate2866(.O (g2174), .I (g1319));
INVX1 gate2867(.O (g6289), .I (I11194));
INVX1 gate2868(.O (g6777), .I (I12202));
INVX1 gate2869(.O (I8802), .I (g3963));
INVX1 gate2870(.O (g6658), .I (g6224));
INVX1 gate2871(.O (g2374), .I (I6220));
INVX1 gate2872(.O (g5448), .I (g5137));
INVX1 gate2873(.O (g1922), .I (g1251));
INVX1 gate2874(.O (I9162), .I (g4272));
INVX1 gate2875(.O (g7556), .I (I13846));
INVX1 gate2876(.O (I13161), .I (g7080));
INVX1 gate2877(.O (I10773), .I (g5708));
INVX1 gate2878(.O (g5055), .I (g4477));
INVX1 gate2879(.O (I12313), .I (g6730));
INVX1 gate2880(.O (g6835), .I (I12376));
INVX1 gate2881(.O (g2985), .I (I6733));
INVX1 gate2882(.O (I9419), .I (g3916));
INVX1 gate2883(.O (I10268), .I (g5471));
INVX1 gate2884(.O (g1581), .I (g710));
INVX1 gate2885(.O (g5827), .I (I10506));
INVX1 gate2886(.O (I12748), .I (g6585));
INVX1 gate2887(.O (g6882), .I (I12517));
INVX1 gate2888(.O (I6042), .I (g237));
INVX1 gate2889(.O (I15651), .I (g9056));
INVX1 gate2890(.O (I15672), .I (g9047));
INVX1 gate2891(.O (g3582), .I (g2407));
INVX1 gate2892(.O (g2284), .I (I6036));
INVX1 gate2893(.O (I5914), .I (g1097));
INVX1 gate2894(.O (I13225), .I (g7095));
INVX1 gate2895(.O (g7064), .I (I12829));
INVX1 gate2896(.O (g2239), .I (I5978));
INVX1 gate2897(.O (I7314), .I (g2916));
INVX1 gate2898(.O (I10180), .I (g4721));
INVX1 gate2899(.O (I16148), .I (g9368));
INVX1 gate2900(.O (g1597), .I (g973));
INVX1 gate2901(.O (g9077), .I (I15625));
INVX1 gate2902(.O (g2180), .I (g1318));
INVX1 gate2903(.O (g5846), .I (g5367));
INVX1 gate2904(.O (g2380), .I (I6242));
INVX1 gate2905(.O (I13258), .I (g6907));
INVX1 gate2906(.O (I12900), .I (g6947));
INVX1 gate2907(.O (I7870), .I (g2827));
INVX1 gate2908(.O (I8901), .I (g4122));
INVX1 gate2909(.O (g2832), .I (g2184));
INVX1 gate2910(.O (I12466), .I (g6687));
INVX1 gate2911(.O (g5396), .I (g4692));
INVX1 gate2912(.O (I5413), .I (g1016));
INVX1 gate2913(.O (g1784), .I (I5636));
INVX1 gate2914(.O (g6799), .I (I12268));
INVX1 gate2915(.O (I6054), .I (g465));
INVX1 gate2916(.O (g2020), .I (I5855));
INVX1 gate2917(.O (I10930), .I (g5600));
INVX1 gate2918(.O (I15513), .I (g8970));
INVX1 gate2919(.O (I11043), .I (g5648));
INVX1 gate2920(.O (I6454), .I (g1868));
INVX1 gate2921(.O (I12101), .I (g5971));
INVX1 gate2922(.O (I6770), .I (g1590));
INVX1 gate2923(.O (g6674), .I (I11978));
INVX1 gate2924(.O (I13244), .I (g7033));
INVX1 gate2925(.O (g7563), .I (I13861));
INVX1 gate2926(.O (g8111), .I (I14374));
INVX1 gate2927(.O (g5780), .I (I10387));
INVX1 gate2928(.O (g4000), .I (g3131));
INVX1 gate2929(.O (I10694), .I (g5445));
INVX1 gate2930(.O (g4126), .I (I7981));
INVX1 gate2931(.O (I10965), .I (g5719));
INVX1 gate2932(.O (g6997), .I (I12737));
INVX1 gate2933(.O (g7295), .I (I13317));
INVX1 gate2934(.O (g2794), .I (g2185));
INVX1 gate2935(.O (I11069), .I (g5671));
INVX1 gate2936(.O (g9104), .I (I15702));
INVX1 gate2937(.O (I5936), .I (g222));
INVX1 gate2938(.O (g9099), .I (I15687));
INVX1 gate2939(.O (I6532), .I (g1694));
INVX1 gate2940(.O (g9304), .I (g9298));
INVX1 gate2941(.O (g2931), .I (I6669));
INVX1 gate2942(.O (g3721), .I (I7211));
INVX1 gate2943(.O (g6238), .I (I11043));
INVX1 gate2944(.O (I6553), .I (g2246));
INVX1 gate2945(.O (g5662), .I (g5027));
INVX1 gate2946(.O (I13810), .I (g7312));
INVX1 gate2947(.O (g8174), .I (I14403));
INVX1 gate2948(.O (g6332), .I (I11323));
INVX1 gate2949(.O (I15717), .I (g9051));
INVX1 gate2950(.O (I11955), .I (g5988));
INVX1 gate2951(.O (g5418), .I (g5100));
INVX1 gate2952(.O (g5467), .I (g4891));
INVX1 gate2953(.O (I9025), .I (g4462));
INVX1 gate2954(.O (g6353), .I (I11386));
INVX1 gate2955(.O (g7194), .I (I13118));
INVX1 gate2956(.O (I13879), .I (g7332));
INVX1 gate2957(.O (I9425), .I (g3917));
INVX1 gate2958(.O (g655), .I (I5383));
INVX1 gate2959(.O (g2905), .I (I6629));
INVX1 gate2960(.O (I6012), .I (g384));
INVX1 gate2961(.O (g6744), .I (I12124));
INVX1 gate2962(.O (g7731), .I (I14064));
INVX1 gate2963(.O (g6802), .I (I12277));
INVX1 gate2964(.O (g8284), .I (I14531));
INVX1 gate2965(.O (g2628), .I (g1573));
INVX1 gate2966(.O (g3502), .I (g1616));
INVX1 gate2967(.O (g8545), .I (g7905));
INVX1 gate2968(.O (I6189), .I (g249));
INVX1 gate2969(.O (g2630), .I (g1575));
INVX1 gate2970(.O (g5493), .I (g4920));
INVX1 gate2971(.O (g8180), .I (g7719));
INVX1 gate2972(.O (I14279), .I (g7700));
INVX1 gate2973(.O (g4608), .I (I8739));
INVX1 gate2974(.O (g4924), .I (g4113));
INVX1 gate2975(.O (I5775), .I (g1240));
INVX1 gate2976(.O (g7966), .I (I14291));
INVX1 gate2977(.O (g2100), .I (g1227));
INVX1 gate2978(.O (g3940), .I (I7623));
INVX1 gate2979(.O (I10469), .I (g5222));
INVX1 gate2980(.O (I11967), .I (g5971));
INVX1 gate2981(.O (I11994), .I (g6195));
INVX1 gate2982(.O (g7471), .I (g7233));
INVX1 gate2983(.O (I15723), .I (g9065));
INVX1 gate2984(.O (g9044), .I (I15536));
INVX1 gate2985(.O (g1942), .I (g828));
INVX1 gate2986(.O (I6029), .I (g1207));
INVX1 gate2987(.O (g4023), .I (I7788));
INVX1 gate2988(.O (I8736), .I (g4008));
INVX1 gate2989(.O (I10286), .I (g5519));
INVX1 gate2990(.O (I6371), .I (g33));
INVX1 gate2991(.O (g1704), .I (I5548));
INVX1 gate2992(.O (g5181), .I (I9669));
INVX1 gate2993(.O (I12008), .I (g5897));
INVX1 gate2994(.O (I9678), .I (g4808));
INVX1 gate2995(.O (I15433), .I (g8911));
INVX1 gate2996(.O (g5847), .I (I10552));
INVX1 gate2997(.O (I6956), .I (g1907));
INVX1 gate2998(.O (g6901), .I (g6525));
INVX1 gate2999(.O (I14039), .I (g7449));
INVX1 gate3000(.O (g4588), .I (g2929));
INVX1 gate3001(.O (I11425), .I (g5872));
INVX1 gate3002(.O (g5685), .I (I10186));
INVX1 gate3003(.O (g5197), .I (g4938));
INVX1 gate3004(.O (I13425), .I (g7166));
INVX1 gate3005(.O (g5397), .I (g5076));
INVX1 gate3006(.O (I8889), .I (g4311));
INVX1 gate3007(.O (g6511), .I (I11693));
INVX1 gate3008(.O (g703), .I (I5398));
INVX1 gate3009(.O (I11458), .I (g6063));
INVX1 gate3010(.O (I15811), .I (g9151));
INVX1 gate3011(.O (I10815), .I (g5418));
INVX1 gate3012(.O (I12454), .I (g6581));
INVX1 gate3013(.O (g2973), .I (g1854));
INVX1 gate3014(.O (g1810), .I (I5676));
INVX1 gate3015(.O (g3430), .I (I6956));
INVX1 gate3016(.O (g4665), .I (I8910));
INVX1 gate3017(.O (I12712), .I (g6543));
INVX1 gate3018(.O (g4051), .I (g3093));
INVX1 gate3019(.O (g6092), .I (g5317));
INVX1 gate3020(.O (I13918), .I (g7361));
INVX1 gate3021(.O (I15971), .I (g9233));
INVX1 gate3022(.O (I8871), .I (g3869));
INVX1 gate3023(.O (I14187), .I (g7728));
INVX1 gate3024(.O (g7150), .I (g6952));
INVX1 gate3025(.O (I14677), .I (g7791));
INVX1 gate3026(.O (g7350), .I (I13466));
INVX1 gate3027(.O (g6864), .I (I12463));
INVX1 gate3028(.O (I7195), .I (g1795));
INVX1 gate3029(.O (g2969), .I (g2393));
INVX1 gate3030(.O (I13444), .I (g7282));
INVX1 gate3031(.O (g6714), .I (I12068));
INVX1 gate3032(.O (g7773), .I (I14190));
INVX1 gate3033(.O (g4146), .I (I8011));
INVX1 gate3034(.O (g7009), .I (I12753));
INVX1 gate3035(.O (g4633), .I (I8814));
INVX1 gate3036(.O (g2323), .I (I6112));
INVX1 gate3037(.O (I10937), .I (g5560));
INVX1 gate3038(.O (I6963), .I (g1558));
INVX1 gate3039(.O (g1568), .I (g658));
INVX1 gate3040(.O (I6109), .I (g1214));
INVX1 gate3041(.O (I6791), .I (g1967));
INVX1 gate3042(.O (g4103), .I (I7922));
INVX1 gate3043(.O (I12567), .I (g6721));
INVX1 gate3044(.O (I6309), .I (g1336));
INVX1 gate3045(.O (g4303), .I (I8268));
INVX1 gate3046(.O (I11086), .I (g5397));
INVX1 gate3047(.O (I7807), .I (g2595));
INVX1 gate3048(.O (g3910), .I (I7523));
INVX1 gate3049(.O (I12238), .I (g6637));
INVX1 gate3050(.O (g7769), .I (I14178));
INVX1 gate3051(.O (I10169), .I (g4873));
INVX1 gate3052(.O (I7859), .I (g2804));
INVX1 gate3053(.O (g4696), .I (I8983));
INVX1 gate3054(.O (g1912), .I (g1524));
INVX1 gate3055(.O (g5631), .I (g4938));
INVX1 gate3056(.O (g7836), .I (I14260));
INVX1 gate3057(.O (I14169), .I (g7715));
INVX1 gate3058(.O (g5723), .I (g4938));
INVX1 gate3059(.O (g4732), .I (I9034));
INVX1 gate3060(.O (g5101), .I (g4259));
INVX1 gate3061(.O (I12382), .I (g6772));
INVX1 gate3062(.O (I5356), .I (g3837));
INVX1 gate3063(.O (g2528), .I (g1260));
INVX1 gate3064(.O (I14410), .I (g7697));
INVX1 gate3065(.O (g2351), .I (g792));
INVX1 gate3066(.O (g2648), .I (I6428));
INVX1 gate3067(.O (I8838), .I (g3967));
INVX1 gate3068(.O (I12176), .I (g5939));
INVX1 gate3069(.O (I8024), .I (g3076));
INVX1 gate3070(.O (I12675), .I (g6510));
INVX1 gate3071(.O (g6736), .I (I12108));
INVX1 gate3072(.O (g8750), .I (g8524));
INVX1 gate3073(.O (I10479), .I (g5227));
INVX1 gate3074(.O (g6968), .I (I12699));
INVX1 gate3075(.O (g2655), .I (g1611));
INVX1 gate3076(.O (g8973), .I (I15423));
INVX1 gate3077(.O (g1929), .I (g1224));
INVX1 gate3078(.O (I12154), .I (g5874));
INVX1 gate3079(.O (I5942), .I (g300));
INVX1 gate3080(.O (I9369), .I (g3901));
INVX1 gate3081(.O (g7229), .I (g6938));
INVX1 gate3082(.O (g6623), .I (I11861));
INVX1 gate3083(.O (g7993), .I (I14298));
INVX1 gate3084(.O (I7255), .I (g1955));
INVX1 gate3085(.O (g6076), .I (g5287));
INVX1 gate3086(.O (I14015), .I (g7440));
INVX1 gate3087(.O (I9407), .I (g4232));
INVX1 gate3088(.O (g6889), .I (I12538));
INVX1 gate3089(.O (I11656), .I (g5772));
INVX1 gate3090(.O (I13656), .I (g7228));
INVX1 gate3091(.O (g3589), .I (I7061));
INVX1 gate3092(.O (g8040), .I (g7699));
INVX1 gate3093(.O (I11353), .I (g5788));
INVX1 gate3094(.O (g9036), .I (I15522));
INVX1 gate3095(.O (g4443), .I (I8449));
INVX1 gate3096(.O (I13353), .I (g7231));
INVX1 gate3097(.O (I11680), .I (g5939));
INVX1 gate3098(.O (g8969), .I (I15411));
INVX1 gate3099(.O (I8477), .I (g3014));
INVX1 gate3100(.O (g9178), .I (I15814));
INVX1 gate3101(.O (g9378), .I (I16158));
INVX1 gate3102(.O (I13144), .I (g7031));
INVX1 gate3103(.O (g4116), .I (I7959));
INVX1 gate3104(.O (g6375), .I (I11452));
INVX1 gate3105(.O (g6871), .I (I12484));
INVX1 gate3106(.O (g4316), .I (I8291));
INVX1 gate3107(.O (I5954), .I (g89));
INVX1 gate3108(.O (g2884), .I (g2238));
INVX1 gate3109(.O (g3861), .I (I7386));
INVX1 gate3110(.O (g5041), .I (I9393));
INVX1 gate3111(.O (g3048), .I (I6784));
INVX1 gate3112(.O (g4034), .I (I7811));
INVX1 gate3113(.O (I9582), .I (g4694));
INVX1 gate3114(.O (I8205), .I (g2655));
INVX1 gate3115(.O (g6651), .I (I11933));
INVX1 gate3116(.O (g9182), .I (g9178));
INVX1 gate3117(.O (I5432), .I (g1176));
INVX1 gate3118(.O (g4565), .I (g2901));
INVX1 gate3119(.O (g8666), .I (I14792));
INVX1 gate3120(.O (g9382), .I (I16168));
INVX1 gate3121(.O (I15959), .I (g9217));
INVX1 gate3122(.O (I15379), .I (g8882));
INVX1 gate3123(.O (I8742), .I (g3919));
INVX1 gate3124(.O (g2372), .I (I6214));
INVX1 gate3125(.O (g3774), .I (g1770));
INVX1 gate3126(.O (I13631), .I (g7248));
INVX1 gate3127(.O (I5568), .I (g1409));
INVX1 gate3128(.O (g8875), .I (I15211));
INVX1 gate3129(.O (g3846), .I (I7341));
INVX1 gate3130(.O (g2618), .I (g1566));
INVX1 gate3131(.O (g1683), .I (g795));
INVX1 gate3132(.O (I16129), .I (g9355));
INVX1 gate3133(.O (g6384), .I (I11479));
INVX1 gate3134(.O (g2235), .I (I5966));
INVX1 gate3135(.O (g2343), .I (g1392));
INVX1 gate3136(.O (g6139), .I (I10780));
INVX1 gate3137(.O (g5168), .I (I9630));
INVX1 gate3138(.O (I12439), .I (g6566));
INVX1 gate3139(.O (g5669), .I (I10154));
INVX1 gate3140(.O (g4697), .I (I8986));
INVX1 gate3141(.O (g6339), .I (I11344));
INVX1 gate3142(.O (g4914), .I (g4093));
INVX1 gate3143(.O (I14531), .I (g8178));
INVX1 gate3144(.O (g2282), .I (g1400));
INVX1 gate3145(.O (I7112), .I (g2546));
INVX1 gate3146(.O (g1778), .I (g613));
INVX1 gate3147(.O (g1894), .I (I5772));
INVX1 gate3148(.O (g5058), .I (I9416));
INVX1 gate3149(.O (g6838), .I (I12385));
INVX1 gate3150(.O (g4596), .I (g3466));
INVX1 gate3151(.O (I8754), .I (g3911));
INVX1 gate3152(.O (g6024), .I (g5494));
INVX1 gate3153(.O (I14178), .I (g7562));
INVX1 gate3154(.O (g4013), .I (g3131));
INVX1 gate3155(.O (g2134), .I (g1317));
INVX1 gate3156(.O (g6795), .I (I12256));
INVX1 gate3157(.O (g3780), .I (g1847));
INVX1 gate3158(.O (I10186), .I (g5129));
INVX1 gate3159(.O (g6737), .I (I12111));
INVX1 gate3160(.O (g2334), .I (I6143));
INVX1 gate3161(.O (I15681), .I (g9063));
INVX1 gate3162(.O (g6809), .I (I12298));
INVX1 gate3163(.O (I8273), .I (g2976));
INVX1 gate3164(.O (I12349), .I (g6742));
INVX1 gate3165(.O (g5743), .I (I10286));
INVX1 gate3166(.O (I6419), .I (g1799));
INVX1 gate3167(.O (I10373), .I (g5722));
INVX1 gate3168(.O (g1782), .I (g624));
INVX1 gate3169(.O (I7676), .I (g2584));
INVX1 gate3170(.O (g2548), .I (g1351));
INVX1 gate3171(.O (I7293), .I (g2955));
INVX1 gate3172(.O (I12906), .I (g6918));
INVX1 gate3173(.O (I15429), .I (g8899));
INVX1 gate3174(.O (I7129), .I (g2495));
INVX1 gate3175(.O (I13023), .I (g7040));
INVX1 gate3176(.O (g1661), .I (g1405));
INVX1 gate3177(.O (I7329), .I (g2920));
INVX1 gate3178(.O (I11224), .I (g6255));
INVX1 gate3179(.O (g6672), .I (I11974));
INVX1 gate3180(.O (g2555), .I (g936));
INVX1 gate3181(.O (g6231), .I (I11028));
INVX1 gate3182(.O (g3018), .I (I6770));
INVX1 gate3183(.O (I11308), .I (g5759));
INVX1 gate3184(.O (g2804), .I (g1796));
INVX1 gate3185(.O (I12304), .I (g6711));
INVX1 gate3186(.O (g9095), .I (I15675));
INVX1 gate3187(.O (I13308), .I (g7169));
INVX1 gate3188(.O (g5734), .I (I10259));
INVX1 gate3189(.O (g1949), .I (g1292));
INVX1 gate3190(.O (g6523), .I (I11707));
INVX1 gate3191(.O (I9502), .I (g3972));
INVX1 gate3192(.O (g3994), .I (g3192));
INVX1 gate3193(.O (I8983), .I (g4536));
INVX1 gate3194(.O (g9102), .I (I15696));
INVX1 gate3195(.O (g9208), .I (g9198));
INVX1 gate3196(.O (I15765), .I (g9039));
INVX1 gate3197(.O (g9302), .I (g9281));
INVX1 gate3198(.O (I8862), .I (g3981));
INVX1 gate3199(.O (g6205), .I (g5628));
INVX1 gate3200(.O (I14334), .I (g7578));
INVX1 gate3201(.O (g8172), .I (I14397));
INVX1 gate3202(.O (I15690), .I (g9074));
INVX1 gate3203(.O (g2621), .I (g1567));
INVX1 gate3204(.O (I8712), .I (g4007));
INVX1 gate3205(.O (I7592), .I (g2712));
INVX1 gate3206(.O (g5074), .I (I9440));
INVX1 gate3207(.O (g3093), .I (g1686));
INVX1 gate3208(.O (I6728), .I (g1959));
INVX1 gate3209(.O (I8543), .I (g2810));
INVX1 gate3210(.O (g5474), .I (g4904));
INVX1 gate3211(.O (g1646), .I (g1214));
INVX1 gate3212(.O (g7298), .I (I13326));
INVX1 gate3213(.O (g4601), .I (I8718));
INVX1 gate3214(.O (I7746), .I (g3591));
INVX1 gate3215(.O (g6634), .I (I11894));
INVX1 gate3216(.O (g8667), .I (I14795));
INVX1 gate3217(.O (I13816), .I (g7455));
INVX1 gate3218(.O (g8235), .I (I14492));
INVX1 gate3219(.O (g2313), .I (I6096));
INVX1 gate3220(.O (g6742), .I (I12120));
INVX1 gate3221(.O (g1603), .I (I5471));
INVX1 gate3222(.O (g6104), .I (g5345));
INVX1 gate3223(.O (I14964), .I (g8406));
INVX1 gate3224(.O (g6304), .I (I11239));
INVX1 gate3225(.O (I15504), .I (g8967));
INVX1 gate3226(.O (g2202), .I (g1321));
INVX1 gate3227(.O (I12138), .I (g5874));
INVX1 gate3228(.O (g4922), .I (g4111));
INVX1 gate3229(.O (I10587), .I (g5439));
INVX1 gate3230(.O (I13752), .I (g7315));
INVX1 gate3231(.O (I11374), .I (g5844));
INVX1 gate3232(.O (g3847), .I (I7344));
INVX1 gate3233(.O (g2908), .I (g2290));
INVX1 gate3234(.O (g5480), .I (g4913));
INVX1 gate3235(.O (I6425), .I (g1811));
INVX1 gate3236(.O (g5713), .I (g4841));
INVX1 gate3237(.O (g4581), .I (g2921));
INVX1 gate3238(.O (I12415), .I (g6410));
INVX1 gate3239(.O (g3700), .I (g2514));
INVX1 gate3240(.O (g9042), .I (I15530));
INVX1 gate3241(.O (g2494), .I (g9));
INVX1 gate3242(.O (I7953), .I (g3542));
INVX1 gate3243(.O (g6754), .I (I12135));
INVX1 gate3244(.O (g1583), .I (g718));
INVX1 gate3245(.O (g5569), .I (I10028));
INVX1 gate3246(.O (g4597), .I (I8706));
INVX1 gate3247(.O (I9564), .I (g4703));
INVX1 gate3248(.O (I5894), .I (g86));
INVX1 gate3249(.O (I11669), .I (g5918));
INVX1 gate3250(.O (g7708), .I (I14005));
INVX1 gate3251(.O (I13669), .I (g7240));
INVX1 gate3252(.O (g9233), .I (I15953));
INVX1 gate3253(.O (g7520), .I (I13740));
INVX1 gate3254(.O (g8792), .I (I14996));
INVX1 gate3255(.O (I11260), .I (g5779));
INVX1 gate3256(.O (g6613), .I (I11835));
INVX1 gate3257(.O (g3950), .I (g3131));
INVX1 gate3258(.O (g4784), .I (I9095));
INVX1 gate3259(.O (I10569), .I (g5417));
INVX1 gate3260(.O (g4739), .I (I9053));
INVX1 gate3261(.O (I11392), .I (g5800));
INVX1 gate3262(.O (g1952), .I (g1333));
INVX1 gate3263(.O (I9910), .I (g4681));
INVX1 gate3264(.O (g6269), .I (I11090));
INVX1 gate3265(.O (g5688), .I (I10193));
INVX1 gate3266(.O (I6006), .I (g306));
INVX1 gate3267(.O (I15533), .I (g9002));
INVX1 gate3268(.O (g2965), .I (g2384));
INVX1 gate3269(.O (g6983), .I (I12722));
INVX1 gate3270(.O (g1616), .I (I5478));
INVX1 gate3271(.O (I14747), .I (g8175));
INVX1 gate3272(.O (g7176), .I (I13084));
INVX1 gate3273(.O (I5475), .I (g1084));
INVX1 gate3274(.O (I7716), .I (g3038));
INVX1 gate3275(.O (g6572), .I (I11764));
INVX1 gate3276(.O (g6862), .I (I12457));
INVX1 gate3277(.O (I11559), .I (g6065));
INVX1 gate3278(.O (g4079), .I (I7864));
INVX1 gate3279(.O (I11525), .I (g5874));
INVX1 gate3280(.O (I11488), .I (g6034));
INVX1 gate3281(.O (I13559), .I (g7177));
INVX1 gate3282(.O (g3562), .I (I7044));
INVX1 gate3283(.O (I12484), .I (g6621));
INVX1 gate3284(.O (I9609), .I (g4780));
INVX1 gate3285(.O (g2264), .I (I5997));
INVX1 gate3286(.O (g6712), .I (I12062));
INVX1 gate3287(.O (g7405), .I (I13518));
INVX1 gate3288(.O (g4668), .I (I8919));
INVX1 gate3289(.O (I6087), .I (g318));
INVX1 gate3290(.O (I6305), .I (g1333));
INVX1 gate3291(.O (g3631), .I (I7098));
INVX1 gate3292(.O (g7829), .I (I14251));
INVX1 gate3293(.O (g2360), .I (g1435));
INVX1 gate3294(.O (g2933), .I (I6673));
INVX1 gate3295(.O (g3723), .I (g2096));
INVX1 gate3296(.O (I12609), .I (g6571));
INVX1 gate3297(.O (g7286), .I (I13290));
INVX1 gate3298(.O (g7765), .I (I14166));
INVX1 gate3299(.O (I7198), .I (g2509));
INVX1 gate3300(.O (I10807), .I (g5294));
INVX1 gate3301(.O (g5000), .I (I9325));
INVX1 gate3302(.O (I5646), .I (g883));
INVX1 gate3303(.O (g8094), .I (g7705));
INVX1 gate3304(.O (I14807), .I (g8603));
INVX1 gate3305(.O (g2641), .I (g1587));
INVX1 gate3306(.O (I14974), .I (g8442));
INVX1 gate3307(.O (I9217), .I (g4443));
INVX1 gate3308(.O (I10639), .I (g5224));
INVX1 gate3309(.O (g4501), .I (g2801));
INVX1 gate3310(.O (g6729), .I (g6263));
INVX1 gate3311(.O (g6961), .I (I12684));
INVX1 gate3312(.O (I13544), .I (g1167));
INVX1 gate3313(.O (g3605), .I (g1938));
INVX1 gate3314(.O (I13865), .I (g7333));
INVX1 gate3315(.O (g2996), .I (g1828));
INVX1 gate3316(.O (I9466), .I (g3943));
INVX1 gate3317(.O (g5760), .I (I10353));
INVX1 gate3318(.O (g9189), .I (I15845));
INVX1 gate3319(.O (g7733), .I (I14070));
INVX1 gate3320(.O (I12921), .I (g6993));
INVX1 gate3321(.O (I13713), .I (g7341));
INVX1 gate3322(.O (g9389), .I (I16183));
INVX1 gate3323(.O (g1970), .I (I5831));
INVX1 gate3324(.O (I6226), .I (g408));
INVX1 gate3325(.O (g7270), .I (I13250));
INVX1 gate3326(.O (I8805), .I (g3976));
INVX1 gate3327(.O (I10265), .I (g5468));
INVX1 gate3328(.O (I8916), .I (g4195));
INVX1 gate3329(.O (g1925), .I (g825));
INVX1 gate3330(.O (g8776), .I (g8585));
INVX1 gate3331(.O (g2724), .I (g1814));
INVX1 gate3332(.O (g7225), .I (g6936));
INVX1 gate3333(.O (g7610), .I (g7450));
INVX1 gate3334(.O (g9029), .I (I15501));
INVX1 gate3335(.O (g6014), .I (I10614));
INVX1 gate3336(.O (I14416), .I (g7727));
INVX1 gate3337(.O (g2379), .I (I6239));
INVX1 gate3338(.O (I13610), .I (g7227));
INVX1 gate3339(.O (I12813), .I (g6607));
INVX1 gate3340(.O (I16145), .I (g9367));
INVX1 gate3341(.O (g6885), .I (I12526));
INVX1 gate3342(.O (I6045), .I (g309));
INVX1 gate3343(.O (g4704), .I (I9001));
INVX1 gate3344(.O (I13042), .I (g6963));
INVX1 gate3345(.O (g6660), .I (I11958));
INVX1 gate3346(.O (g6946), .I (I12649));
INVX1 gate3347(.O (I13255), .I (g7057));
INVX1 gate3348(.O (g2878), .I (g2233));
INVX1 gate3349(.O (I13189), .I (g7002));
INVX1 gate3350(.O (I7644), .I (g2584));
INVX1 gate3351(.O (g5183), .I (I9675));
INVX1 gate3352(.O (I13679), .I (g7259));
INVX1 gate3353(.O (g7124), .I (g6896));
INVX1 gate3354(.O (I12973), .I (g6927));
INVX1 gate3355(.O (g5608), .I (g4969));
INVX1 gate3356(.O (I9333), .I (g4245));
INVX1 gate3357(.O (g2289), .I (I6051));
INVX1 gate3358(.O (g6903), .I (I12582));
INVX1 gate3359(.O (g2777), .I (g1797));
INVX1 gate3360(.O (g9281), .I (I16009));
INVX1 gate3361(.O (g5779), .I (I10384));
INVX1 gate3362(.O (I10579), .I (g5433));
INVX1 gate3363(.O (I9774), .I (g4678));
INVX1 gate3364(.O (g4250), .I (I8177));
INVX1 gate3365(.O (g2882), .I (g2236));
INVX1 gate3366(.O (I11686), .I (g6076));
INVX1 gate3367(.O (I11939), .I (g6015));
INVX1 gate3368(.O (I7867), .I (g2818));
INVX1 gate3369(.O (g9297), .I (I16017));
INVX1 gate3370(.O (I13460), .I (g7263));
INVX1 gate3371(.O (g4032), .I (I7807));
INVX1 gate3372(.O (I11383), .I (g5827));
INVX1 gate3373(.O (g2271), .I (I6018));
INVX1 gate3374(.O (I9396), .I (g3908));
INVX1 gate3375(.O (I13383), .I (g7275));
INVX1 gate3376(.O (g1789), .I (g1034));
INVX1 gate3377(.O (g7206), .I (I13134));
INVX1 gate3378(.O (I6578), .I (g1603));
INVX1 gate3379(.O (I6868), .I (g530));
INVX1 gate3380(.O (I5616), .I (g979));
INVX1 gate3381(.O (g6036), .I (I10643));
INVX1 gate3382(.O (I13267), .I (g6913));
INVX1 gate3383(.O (g6378), .I (I11461));
INVX1 gate3384(.O (I6767), .I (g1933));
INVX1 gate3385(.O (g5161), .I (I9609));
INVX1 gate3386(.O (I16132), .I (g9356));
INVX1 gate3387(.O (I10442), .I (g5215));
INVX1 gate3388(.O (I15498), .I (g8974));
INVX1 gate3389(.O (g1987), .I (I5842));
INVX1 gate3390(.O (g1771), .I (g609));
INVX1 gate3391(.O (I7211), .I (g1742));
INVX1 gate3392(.O (g7287), .I (I13293));
INVX1 gate3393(.O (I14442), .I (g8065));
INVX1 gate3394(.O (g6135), .I (I10770));
INVX1 gate3395(.O (I5404), .I (g722));
INVX1 gate3396(.O (g4568), .I (g2904));
INVX1 gate3397(.O (I7386), .I (g3013));
INVX1 gate3398(.O (g5665), .I (g4748));
INVX1 gate3399(.O (g9109), .I (I15717));
INVX1 gate3400(.O (g5051), .I (I9407));
INVX1 gate3401(.O (g6335), .I (I11332));
INVX1 gate3402(.O (g6831), .I (I12364));
INVX1 gate3403(.O (g9309), .I (I16043));
INVX1 gate3404(.O (g3531), .I (g1616));
INVX1 gate3405(.O (g5127), .I (I9525));
INVX1 gate3406(.O (g2674), .I (g1675));
INVX1 gate3407(.O (g6288), .I (I11191));
INVX1 gate3408(.O (g6382), .I (I11473));
INVX1 gate3409(.O (I16161), .I (g9363));
INVX1 gate3410(.O (g8179), .I (I14416));
INVX1 gate3411(.O (I9018), .I (g3872));
INVX1 gate3412(.O (g3743), .I (g1776));
INVX1 gate3413(.O (I7599), .I (g2734));
INVX1 gate3414(.O (I15924), .I (g9207));
INVX1 gate3415(.O (I6015), .I (g437));
INVX1 gate3416(.O (I12400), .I (g6767));
INVX1 gate3417(.O (g4357), .I (g3679));
INVX1 gate3418(.O (g5146), .I (I9564));
INVX1 gate3419(.O (g6805), .I (I12286));
INVX1 gate3420(.O (g5633), .I (g4895));
INVX1 gate3421(.O (I11218), .I (g6161));
INVX1 gate3422(.O (I12214), .I (g6507));
INVX1 gate3423(.O (g7781), .I (I14214));
INVX1 gate3424(.O (g2238), .I (I5975));
INVX1 gate3425(.O (g2332), .I (g926));
INVX1 gate3426(.O (I10430), .I (g5211));
INVX1 gate3427(.O (I13837), .I (g7324));
INVX1 gate3428(.O (g3856), .I (I7371));
INVX1 gate3429(.O (g2680), .I (g1665));
INVX1 gate3430(.O (I14430), .I (g7836));
INVX1 gate3431(.O (g2209), .I (I5926));
INVX1 gate3432(.O (g2353), .I (g871));
INVX1 gate3433(.O (I9493), .I (g4426));
INVX1 gate3434(.O (g4929), .I (g4120));
INVX1 gate3435(.O (g9201), .I (g9183));
INVX1 gate3436(.O (I12328), .I (g6760));
INVX1 gate3437(.O (I15753), .I (g9080));
INVX1 gate3438(.O (g5696), .I (I10207));
INVX1 gate3439(.O (g8882), .I (I15222));
INVX1 gate3440(.O (g1945), .I (g1081));
INVX1 gate3441(.O (g6947), .I (I12652));
INVX1 gate3442(.O (g7510), .I (I13710));
INVX1 gate3443(.O (g7245), .I (I13193));
INVX1 gate3444(.O (g6798), .I (I12265));
INVX1 gate3445(.O (I12538), .I (g6606));
INVX1 gate3446(.O (g1738), .I (g741));
INVX1 gate3447(.O (g3074), .I (I6800));
INVX1 gate3448(.O (I16043), .I (g9285));
INVX1 gate3449(.O (g5732), .I (I10253));
INVX1 gate3450(.O (g7291), .I (I13305));
INVX1 gate3451(.O (g3992), .I (I7723));
INVX1 gate3452(.O (I14035), .I (g7310));
INVX1 gate3453(.O (I15199), .I (g8792));
INVX1 gate3454(.O (I10684), .I (g5258));
INVX1 gate3455(.O (I11455), .I (g6087));
INVX1 gate3456(.O (g4626), .I (I8793));
INVX1 gate3457(.O (I8233), .I (g3588));
INVX1 gate3458(.O (I11470), .I (g6095));
INVX1 gate3459(.O (g5240), .I (I9752));
INVX1 gate3460(.O (g7344), .I (g7150));
INVX1 gate3461(.O (I13617), .I (g7276));
INVX1 gate3462(.O (g5072), .I (g4457));
INVX1 gate3463(.O (g9098), .I (I15684));
INVX1 gate3464(.O (I13915), .I (g7360));
INVX1 gate3465(.O (g8799), .I (I15007));
INVX1 gate3466(.O (I12241), .I (g6640));
INVX1 gate3467(.O (I14142), .I (g7551));
INVX1 gate3468(.O (g1907), .I (g52));
INVX1 gate3469(.O (g5472), .I (I9892));
INVX1 gate3470(.O (I9021), .I (g4489));
INVX1 gate3471(.O (g6873), .I (I12490));
INVX1 gate3472(.O (g7207), .I (I13137));
INVX1 gate3473(.O (g6632), .I (I11890));
INVX1 gate3474(.O (g6095), .I (I10719));
INVX1 gate3475(.O (g3080), .I (g1679));
INVX1 gate3476(.O (g8674), .I (I14816));
INVX1 gate3477(.O (g6037), .I (I10646));
INVX1 gate3478(.O (g3573), .I (g2424));
INVX1 gate3479(.O (I15696), .I (g9050));
INVX1 gate3480(.O (g3863), .I (I7392));
INVX1 gate3481(.O (I5789), .I (g1524));
INVX1 gate3482(.O (g1959), .I (g1252));
INVX1 gate3483(.O (g2901), .I (g2284));
INVX1 gate3484(.O (g7259), .I (g7060));
INVX1 gate3485(.O (g6653), .I (I11939));
INVX1 gate3486(.O (I13277), .I (g7078));
INVX1 gate3487(.O (g6102), .I (g5345));
INVX1 gate3488(.O (g6208), .I (I10965));
INVX1 gate3489(.O (g6302), .I (I11233));
INVX1 gate3490(.O (g8541), .I (g8094));
INVX1 gate3491(.O (I13075), .I (g6958));
INVX1 gate3492(.O (g2511), .I (g1328));
INVX1 gate3493(.O (I7061), .I (g2457));
INVX1 gate3494(.O (g6869), .I (I12478));
INVX1 gate3495(.O (g1876), .I (g77));
INVX1 gate3496(.O (I12771), .I (g6735));
INVX1 gate3497(.O (I11467), .I (g6064));
INVX1 gate3498(.O (I11494), .I (g6037));
INVX1 gate3499(.O (I13595), .I (g7216));
INVX1 gate3500(.O (g7488), .I (g7225));
INVX1 gate3501(.O (I12235), .I (g6634));
INVX1 gate3502(.O (g2092), .I (g1225));
INVX1 gate3503(.O (g5434), .I (g5112));
INVX1 gate3504(.O (I10193), .I (g4670));
INVX1 gate3505(.O (I11037), .I (g5299));
INVX1 gate3506(.O (I14130), .I (g7592));
INVX1 gate3507(.O (I14193), .I (g7532));
INVX1 gate3508(.O (g6752), .I (I12131));
INVX1 gate3509(.O (g5147), .I (I9567));
INVX1 gate3510(.O (I13782), .I (g7498));
INVX1 gate3511(.O (I11984), .I (g6246));
INVX1 gate3512(.O (g8802), .I (I15014));
INVX1 gate3513(.O (I11419), .I (g5835));
INVX1 gate3514(.O (I6428), .I (g1818));
INVX1 gate3515(.O (g9019), .I (I15481));
INVX1 gate3516(.O (g9362), .I (I16122));
INVX1 gate3517(.O (I13419), .I (g7277));
INVX1 gate3518(.O (g3857), .I (I7374));
INVX1 gate3519(.O (g7951), .I (I14288));
INVX1 gate3520(.O (I8706), .I (g3828));
INVX1 gate3521(.O (g3976), .I (I7697));
INVX1 gate3522(.O (I15225), .I (g8689));
INVX1 gate3523(.O (I15708), .I (g9072));
INVX1 gate3524(.O (I13822), .I (g7459));
INVX1 gate3525(.O (I10475), .I (g5529));
INVX1 gate3526(.O (I9301), .I (g4295));
INVX1 gate3527(.O (g7114), .I (I12930));
INVX1 gate3528(.O (I11266), .I (g5794));
INVX1 gate3529(.O (g4661), .I (I8898));
INVX1 gate3530(.O (g6786), .I (I12229));
INVX1 gate3531(.O (I7145), .I (g2501));
INVX1 gate3532(.O (I6564), .I (g2073));
INVX1 gate3533(.O (g4075), .I (I7856));
INVX1 gate3534(.O (I5945), .I (g333));
INVX1 gate3535(.O (I8787), .I (g4012));
INVX1 gate3536(.O (g4475), .I (g3818));
INVX1 gate3537(.O (g5596), .I (g4841));
INVX1 gate3538(.O (g1663), .I (g1416));
INVX1 gate3539(.O (I6826), .I (g2185));
INVX1 gate3540(.O (g6364), .I (I11419));
INVX1 gate3541(.O (g7870), .I (I14270));
INVX1 gate3542(.O (g5013), .I (I9341));
INVX1 gate3543(.O (g4627), .I (I8796));
INVX1 gate3544(.O (I5709), .I (g901));
INVX1 gate3545(.O (g8511), .I (I14646));
INVX1 gate3546(.O (g9086), .I (I15648));
INVX1 gate3547(.O (g1824), .I (I5706));
INVX1 gate3548(.O (I5478), .I (g1148));
INVX1 gate3549(.O (g6296), .I (I11215));
INVX1 gate3550(.O (I11194), .I (g6243));
INVX1 gate3551(.O (g4646), .I (I8853));
INVX1 gate3552(.O (I7107), .I (g2480));
INVX1 gate3553(.O (g2623), .I (g1585));
INVX1 gate3554(.O (g6725), .I (I12091));
INVX1 gate3555(.O (I9585), .I (g4697));
INVX1 gate3556(.O (I10347), .I (g5706));
INVX1 gate3557(.O (I10253), .I (g5240));
INVX1 gate3558(.O (g5820), .I (I10485));
INVX1 gate3559(.O (I7359), .I (g2871));
INVX1 gate3560(.O (g9185), .I (I15833));
INVX1 gate3561(.O (g4084), .I (I7875));
INVX1 gate3562(.O (g4603), .I (I8724));
INVX1 gate3563(.O (I5435), .I (g1461));
INVX1 gate3564(.O (g7336), .I (I13428));
INVX1 gate3565(.O (I13524), .I (g7151));
INVX1 gate3566(.O (I15657), .I (g9059));
INVX1 gate3567(.O (g9385), .I (I16173));
INVX1 gate3568(.O (g8864), .I (I15178));
INVX1 gate3569(.O (I15068), .I (g8638));
INVX1 gate3570(.O (g7768), .I (I14175));
INVX1 gate3571(.O (g1590), .I (I5466));
INVX1 gate3572(.O (g1877), .I (g595));
INVX1 gate3573(.O (I11401), .I (g5828));
INVX1 gate3574(.O (g6553), .I (I11725));
INVX1 gate3575(.O (g9070), .I (I15604));
INVX1 gate3576(.O (g7594), .I (I13927));
INVX1 gate3577(.O (I8745), .I (g3929));
INVX1 gate3578(.O (I10236), .I (g5014));
INVX1 gate3579(.O (g2375), .I (I6223));
INVX1 gate3580(.O (g2871), .I (I6587));
INVX1 gate3581(.O (I12725), .I (g6565));
INVX1 gate3582(.O (g3220), .I (g1889));
INVX1 gate3583(.O (I15337), .I (g8802));
INVX1 gate3584(.O (g2651), .I (I6437));
INVX1 gate3585(.O (I6217), .I (g105));
INVX1 gate3586(.O (g6012), .I (g5367));
INVX1 gate3587(.O (g1556), .I (g65));
INVX1 gate3588(.O (I13118), .I (g7068));
INVX1 gate3589(.O (g3779), .I (g2511));
INVX1 gate3590(.O (g4583), .I (g2924));
INVX1 gate3591(.O (I11864), .I (g5753));
INVX1 gate3592(.O (I14175), .I (g7718));
INVX1 gate3593(.O (g2285), .I (I6039));
INVX1 gate3594(.O (I7115), .I (g2547));
INVX1 gate3595(.O (g6189), .I (I10930));
INVX1 gate3596(.O (I8808), .I (g4014));
INVX1 gate3597(.O (g6389), .I (I11494));
INVX1 gate3598(.O (I7811), .I (g3019));
INVX1 gate3599(.O (I16158), .I (g9363));
INVX1 gate3600(.O (I9669), .I (g4909));
INVX1 gate3601(.O (I13749), .I (g7313));
INVX1 gate3602(.O (g7887), .I (I14273));
INVX1 gate3603(.O (g7122), .I (I12958));
INVX1 gate3604(.O (g4919), .I (g4104));
INVX1 gate3605(.O (g3977), .I (g3160));
INVX1 gate3606(.O (I6571), .I (g1711));
INVX1 gate3607(.O (g6888), .I (I12535));
INVX1 gate3608(.O (I6048), .I (g387));
INVX1 gate3609(.O (I10516), .I (g5241));
INVX1 gate3610(.O (g5581), .I (g4969));
INVX1 gate3611(.O (I14264), .I (g7698));
INVX1 gate3612(.O (g3588), .I (g2379));
INVX1 gate3613(.O (I9531), .I (g4463));
INVX1 gate3614(.O (g2184), .I (I5911));
INVX1 gate3615(.O (I6711), .I (g1726));
INVX1 gate3616(.O (g6371), .I (I11440));
INVX1 gate3617(.O (g1785), .I (g615));
INVX1 gate3618(.O (g6787), .I (I12232));
INVX1 gate3619(.O (g8968), .I (I15408));
INVX1 gate3620(.O (g2384), .I (I6254));
INVX1 gate3621(.O (I11704), .I (g6076));
INVX1 gate3622(.O (g5060), .I (I9422));
INVX1 gate3623(.O (I13704), .I (g7352));
INVX1 gate3624(.O (I11305), .I (g5807));
INVX1 gate3625(.O (g9331), .I (g9321));
INVX1 gate3626(.O (g6956), .I (I12669));
INVX1 gate3627(.O (I13305), .I (g7168));
INVX1 gate3628(.O (g5460), .I (g4684));
INVX1 gate3629(.O (g5597), .I (g4969));
INVX1 gate3630(.O (I11254), .I (g5793));
INVX1 gate3631(.O (g7433), .I (I13562));
INVX1 gate3632(.O (g6675), .I (I11981));
INVX1 gate3633(.O (g4616), .I (I8763));
INVX1 gate3634(.O (I11809), .I (g6285));
INVX1 gate3635(.O (I11900), .I (g5847));
INVX1 gate3636(.O (g4561), .I (g2900));
INVX1 gate3637(.O (g3051), .I (I6791));
INVX1 gate3638(.O (I13900), .I (g7356));
INVX1 gate3639(.O (I6333), .I (g1345));
INVX1 gate3640(.O (I13466), .I (g7122));
INVX1 gate3641(.O (I9505), .I (g4300));
INVX1 gate3642(.O (g1563), .I (g639));
INVX1 gate3643(.O (g2424), .I (g1329));
INVX1 gate3644(.O (I12141), .I (g5897));
INVX1 gate3645(.O (g2795), .I (g1801));
INVX1 gate3646(.O (I8449), .I (g3630));
INVX1 gate3647(.O (I12652), .I (g6664));
INVX1 gate3648(.O (g9087), .I (I15651));
INVX1 gate3649(.O (g9105), .I (I15705));
INVX1 gate3650(.O (g5784), .I (I10397));
INVX1 gate3651(.O (g4004), .I (g2845));
INVX1 gate3652(.O (I15010), .I (g8584));
INVX1 gate3653(.O (I15918), .I (g9211));
INVX1 gate3654(.O (g9305), .I (I16033));
INVX1 gate3655(.O (g5739), .I (I10274));
INVX1 gate3656(.O (I8865), .I (g4032));
INVX1 gate3657(.O (g7496), .I (I13666));
INVX1 gate3658(.O (g4527), .I (g3466));
INVX1 gate3659(.O (g7550), .I (I13834));
INVX1 gate3660(.O (g6297), .I (I11218));
INVX1 gate3661(.O (g3999), .I (I7738));
INVX1 gate3662(.O (g4647), .I (I8856));
INVX1 gate3663(.O (g8175), .I (I14406));
INVX1 gate3664(.O (I8715), .I (g3903));
INVX1 gate3665(.O (I7595), .I (g2573));
INVX1 gate3666(.O (g8871), .I (I15199));
INVX1 gate3667(.O (g3633), .I (I7104));
INVX1 gate3668(.O (g2672), .I (I6471));
INVX1 gate3669(.O (g2231), .I (I5954));
INVX1 gate3670(.O (g7137), .I (I12993));
INVX1 gate3671(.O (I14208), .I (g7711));
INVX1 gate3672(.O (g8651), .I (I14747));
INVX1 gate3673(.O (g2477), .I (g25));
INVX1 gate3674(.O (I16017), .I (g9264));
INVX1 gate3675(.O (g2643), .I (g1589));
INVX1 gate3676(.O (g6684), .I (I11998));
INVX1 gate3677(.O (I12135), .I (g5988));
INVX1 gate3678(.O (g6639), .I (g6198));
INVX1 gate3679(.O (g5668), .I (I10151));
INVX1 gate3680(.O (g6338), .I (I11341));
INVX1 gate3681(.O (I15598), .I (g8991));
INVX1 gate3682(.O (I6509), .I (g1684));
INVX1 gate3683(.O (g5294), .I (g5087));
INVX1 gate3684(.O (g4503), .I (I8565));
INVX1 gate3685(.O (g5840), .I (I10535));
INVX1 gate3686(.O (g6963), .I (I12690));
INVX1 gate3687(.O (I7978), .I (g3574));
INVX1 gate3688(.O (g6791), .I (I12244));
INVX1 gate3689(.O (g2205), .I (g13));
INVX1 gate3690(.O (I12406), .I (g6773));
INVX1 gate3691(.O (g6309), .I (I11254));
INVX1 gate3692(.O (g5190), .I (g4938));
INVX1 gate3693(.O (g4925), .I (g4114));
INVX1 gate3694(.O (I5657), .I (g921));
INVX1 gate3695(.O (I12361), .I (g6765));
INVX1 gate3696(.O (I7417), .I (g3659));
INVX1 gate3697(.O (g3732), .I (g2533));
INVX1 gate3698(.O (I6018), .I (g462));
INVX1 gate3699(.O (g1557), .I (I5432));
INVX1 gate3700(.O (g2634), .I (g1578));
INVX1 gate3701(.O (g3753), .I (g2540));
INVX1 gate3702(.O (I10614), .I (g5302));
INVX1 gate3703(.O (g6808), .I (I12295));
INVX1 gate3704(.O (I9573), .I (g4701));
INVX1 gate3705(.O (g9045), .I (I15539));
INVX1 gate3706(.O (I10436), .I (g5213));
INVX1 gate3707(.O (g724), .I (I5401));
INVX1 gate3708(.O (I14614), .I (g7832));
INVX1 gate3709(.O (g7266), .I (I13238));
INVX1 gate3710(.O (g2551), .I (g1360));
INVX1 gate3711(.O (I14436), .I (g7904));
INVX1 gate3712(.O (g2104), .I (I5879));
INVX1 gate3713(.O (g3944), .I (I7635));
INVX1 gate3714(.O (I11693), .I (g6076));
INVX1 gate3715(.O (g5156), .I (I9594));
INVX1 gate3716(.O (g9373), .I (I16145));
INVX1 gate3717(.O (g9091), .I (I15663));
INVX1 gate3718(.O (g4120), .I (I7967));
INVX1 gate3719(.O (I16023), .I (g9267));
INVX1 gate3720(.O (I7629), .I (g3633));
INVX1 gate3721(.O (g6759), .I (I12148));
INVX1 gate3722(.O (I10274), .I (g5524));
INVX1 gate3723(.O (I14073), .I (g7627));
INVX1 gate3724(.O (I6093), .I (g468));
INVX1 gate3725(.O (I8268), .I (g2801));
INVX1 gate3726(.O (I13009), .I (g6935));
INVX1 gate3727(.O (g1948), .I (g1250));
INVX1 gate3728(.O (g8809), .I (I15065));
INVX1 gate3729(.O (g7142), .I (I13012));
INVX1 gate3730(.O (g6201), .I (I10946));
INVX1 gate3731(.O (g2926), .I (g2325));
INVX1 gate3732(.O (g7342), .I (I13444));
INVX1 gate3733(.O (I11008), .I (g5693));
INVX1 gate3734(.O (g9369), .I (I16135));
INVX1 gate3735(.O (I10565), .I (g5402));
INVX1 gate3736(.O (g6957), .I (I12672));
INVX1 gate3737(.O (g7255), .I (I13209));
INVX1 gate3738(.O (g4617), .I (I8766));
INVX1 gate3739(.O (I8452), .I (g2816));
INVX1 gate3740(.O (g649), .I (I5380));
INVX1 gate3741(.O (g8672), .I (I14810));
INVX1 gate3742(.O (g3316), .I (I6930));
INVX1 gate3743(.O (g9059), .I (I15571));
INVX1 gate3744(.O (I11476), .I (g6194));
INVX1 gate3745(.O (I11485), .I (g6137));
INVX1 gate3746(.O (I7800), .I (g2605));
INVX1 gate3747(.O (g6449), .I (I11596));
INVX1 gate3748(.O (g2273), .I (I6024));
INVX1 gate3749(.O (g1814), .I (g630));
INVX1 gate3750(.O (g6865), .I (I12466));
INVX1 gate3751(.O (I7554), .I (g2573));
INVX1 gate3752(.O (g7097), .I (I12881));
INVX1 gate3753(.O (g7726), .I (I14049));
INVX1 gate3754(.O (I13454), .I (g7147));
INVX1 gate3755(.O (g7497), .I (I13669));
INVX1 gate3756(.O (I10292), .I (g5577));
INVX1 gate3757(.O (g2044), .I (I5861));
INVX1 gate3758(.O (g7354), .I (I13478));
INVX1 gate3759(.O (g5163), .I (I9615));
INVX1 gate3760(.O (g6604), .I (I11818));
INVX1 gate3761(.O (g5810), .I (I10463));
INVX1 gate3762(.O (I13570), .I (g7198));
INVX1 gate3763(.O (I6021), .I (g495));
INVX1 gate3764(.O (g6498), .I (I11666));
INVX1 gate3765(.O (g2269), .I (I6012));
INVX1 gate3766(.O (g1773), .I (g610));
INVX1 gate3767(.O (I8486), .I (g2824));
INVX1 gate3768(.O (I10409), .I (g5204));
INVX1 gate3769(.O (g4547), .I (g3466));
INVX1 gate3770(.O (g5053), .I (g4438));
INVX1 gate3771(.O (g6833), .I (I12370));
INVX1 gate3772(.O (I8730), .I (g3987));
INVX1 gate3773(.O (g3533), .I (g2397));
INVX1 gate3774(.O (g5453), .I (g4680));
INVX1 gate3775(.O (g2862), .I (I6578));
INVX1 gate3776(.O (I15631), .I (g9003));
INVX1 gate3777(.O (I12463), .I (g6682));
INVX1 gate3778(.O (g4892), .I (I9250));
INVX1 gate3779(.O (I11239), .I (g6173));
INVX1 gate3780(.O (g2712), .I (g2039));
INVX1 gate3781(.O (I14136), .I (g7633));
INVX1 gate3782(.O (g9227), .I (I15947));
INVX1 gate3783(.O (g1769), .I (I5609));
INVX1 gate3784(.O (I9126), .I (g3870));
INVX1 gate3785(.O (I7902), .I (g2709));
INVX1 gate3786(.O (g2543), .I (g1348));
INVX1 gate3787(.O (g6896), .I (I12561));
INVX1 gate3788(.O (I13238), .I (g6900));
INVX1 gate3789(.O (I9760), .I (g4838));
INVX1 gate3790(.O (g3013), .I (I6764));
INVX1 gate3791(.O (g1918), .I (g822));
INVX1 gate3792(.O (g1967), .I (g1432));
INVX1 gate3793(.O (g7112), .I (I12924));
INVX1 gate3794(.O (g7267), .I (I13241));
INVX1 gate3795(.O (I5966), .I (g278));
INVX1 gate3796(.O (g5157), .I (I9597));
INVX1 gate3797(.O (g2961), .I (I6711));
INVX1 gate3798(.O (g4738), .I (I9050));
INVX1 gate3799(.O (g8754), .I (g8524));
INVX1 gate3800(.O (I5471), .I (g1029));
INVX1 gate3801(.O (g6019), .I (g5367));
INVX1 gate3802(.O (g6362), .I (I11413));
INVX1 gate3803(.O (I13185), .I (g7020));
INVX1 gate3804(.O (I6723), .I (g2052));
INVX1 gate3805(.O (I13092), .I (g7047));
INVX1 gate3806(.O (g7293), .I (I13311));
INVX1 gate3807(.O (g2927), .I (I6663));
INVX1 gate3808(.O (I12514), .I (g6605));
INVX1 gate3809(.O (I5948), .I (g378));
INVX1 gate3810(.O (g3936), .I (I7605));
INVX1 gate3811(.O (I13518), .I (g7141));
INVX1 gate3812(.O (g7129), .I (I12973));
INVX1 gate3813(.O (I15571), .I (g8982));
INVX1 gate3814(.O (I15308), .I (g8799));
INVX1 gate3815(.O (g1822), .I (g761));
INVX1 gate3816(.O (g7329), .I (I13407));
INVX1 gate3817(.O (g7761), .I (I14154));
INVX1 gate3818(.O (g4907), .I (g4087));
INVX1 gate3819(.O (g2885), .I (g2239));
INVX1 gate3820(.O (g4035), .I (I7814));
INVX1 gate3821(.O (g2660), .I (I6451));
INVX1 gate3822(.O (g2946), .I (g2365));
INVX1 gate3823(.O (I12421), .I (g6486));
INVX1 gate3824(.O (I14109), .I (g7590));
INVX1 gate3825(.O (g7727), .I (I14052));
INVX1 gate3826(.O (I15495), .I (g8973));
INVX1 gate3827(.O (g4482), .I (I8520));
INVX1 gate3828(.O (I7964), .I (g3488));
INVX1 gate3829(.O (g2903), .I (g2286));
INVX1 gate3830(.O (g5626), .I (g4748));
INVX1 gate3831(.O (g7592), .I (I13921));
INVX1 gate3832(.O (I8766), .I (g3960));
INVX1 gate3833(.O (I9588), .I (g4704));
INVX1 gate3834(.O (g6486), .I (I11648));
INVX1 gate3835(.O (I8105), .I (g3339));
INVX1 gate3836(.O (I10283), .I (g5643));
INVX1 gate3837(.O (g4656), .I (I8883));
INVX1 gate3838(.O (g7746), .I (I14109));
INVX1 gate3839(.O (g6730), .I (I12098));
INVX1 gate3840(.O (g9188), .I (I15842));
INVX1 gate3841(.O (g7221), .I (I13157));
INVX1 gate3842(.O (I15687), .I (g9071));
INVX1 gate3843(.O (g9388), .I (I16180));
INVX1 gate3844(.O (g3922), .I (I7561));
INVX1 gate3845(.O (I15985), .I (g9237));
INVX1 gate3846(.O (I14492), .I (g7829));
INVX1 gate3847(.O (g9216), .I (I15924));
INVX1 gate3848(.O (g6385), .I (I11482));
INVX1 gate3849(.O (g6881), .I (I12514));
INVX1 gate3850(.O (I12541), .I (g6614));
INVX1 gate3851(.O (I8748), .I (g3997));
INVX1 gate3852(.O (g4915), .I (g4094));
INVX1 gate3853(.O (I11215), .I (g6156));
INVX1 gate3854(.O (g9028), .I (I15498));
INVX1 gate3855(.O (g6070), .I (g5317));
INVX1 gate3856(.O (I11729), .I (g5772));
INVX1 gate3857(.O (g1895), .I (I5775));
INVX1 gate3858(.O (g6897), .I (I12564));
INVX1 gate3859(.O (g1837), .I (g1007));
INVX1 gate3860(.O (I13577), .I (g7186));
INVX1 gate3861(.O (g9030), .I (I15504));
INVX1 gate3862(.O (g6025), .I (g5367));
INVX1 gate3863(.O (I6673), .I (g2246));
INVX1 gate3864(.O (g6425), .I (I11556));
INVX1 gate3865(.O (I14381), .I (g7596));
INVX1 gate3866(.O (I13728), .I (g7439));
INVX1 gate3867(.O (g5683), .I (I10180));
INVX1 gate3868(.O (I12325), .I (g6755));
INVX1 gate3869(.O (I9633), .I (g4800));
INVX1 gate3870(.O (g2288), .I (I6048));
INVX1 gate3871(.O (I7118), .I (g2484));
INVX1 gate3872(.O (I7167), .I (g2505));
INVX1 gate3873(.O (I14091), .I (g7589));
INVX1 gate3874(.O (g2382), .I (I6248));
INVX1 gate3875(.O (g7068), .I (g6556));
INVX1 gate3876(.O (I12829), .I (g6441));
INVX1 gate3877(.O (I12535), .I (g6599));
INVX1 gate3878(.O (I15669), .I (g9045));
INVX1 gate3879(.O (g3784), .I (g1768));
INVX1 gate3880(.O (I10796), .I (g5397));
INVX1 gate3881(.O (g8014), .I (g7564));
INVX1 gate3882(.O (I9103), .I (g4374));
INVX1 gate3883(.O (I12358), .I (g6761));
INVX1 gate3884(.O (I13438), .I (g7143));
INVX1 gate3885(.O (g3739), .I (g2536));
INVX1 gate3886(.O (I6669), .I (g1698));
INVX1 gate3887(.O (g4663), .I (I8904));
INVX1 gate3888(.O (I6368), .I (g20));
INVX1 gate3889(.O (g2916), .I (I6646));
INVX1 gate3890(.O (I15842), .I (g9171));
INVX1 gate3891(.O (I8373), .I (g3783));
INVX1 gate3892(.O (g5735), .I (I10262));
INVX1 gate3893(.O (g1788), .I (g984));
INVX1 gate3894(.O (g3995), .I (I7728));
INVX1 gate3895(.O (g3937), .I (g2845));
INVX1 gate3896(.O (g8903), .I (I15315));
INVX1 gate3897(.O (g3079), .I (g1603));
INVX1 gate3898(.O (g5782), .I (I10393));
INVX1 gate3899(.O (g4002), .I (g3192));
INVX1 gate3900(.O (I10390), .I (g5195));
INVX1 gate3901(.O (I13906), .I (g7358));
INVX1 gate3902(.O (I11284), .I (g5795));
INVX1 gate3903(.O (I13284), .I (g7156));
INVX1 gate3904(.O (g6131), .I (g5529));
INVX1 gate3905(.O (g7576), .I (I13873));
INVX1 gate3906(.O (g6331), .I (I11320));
INVX1 gate3907(.O (g5075), .I (I9443));
INVX1 gate3908(.O (g3840), .I (I7323));
INVX1 gate3909(.O (g2947), .I (I6695));
INVX1 gate3910(.O (g7716), .I (I14025));
INVX1 gate3911(.O (g7149), .I (I13031));
INVX1 gate3912(.O (g2798), .I (g1787));
INVX1 gate3913(.O (I11622), .I (g5847));
INVX1 gate3914(.O (g1842), .I (g764));
INVX1 gate3915(.O (g7349), .I (I13463));
INVX1 gate3916(.O (g6635), .I (I11897));
INVX1 gate3917(.O (I13622), .I (g7279));
INVX1 gate3918(.O (g9108), .I (I15714));
INVX1 gate3919(.O (g3390), .I (I6949));
INVX1 gate3920(.O (g9308), .I (I16040));
INVX1 gate3921(.O (I8868), .I (g4035));
INVX1 gate3922(.O (g5627), .I (g4673));
INVX1 gate3923(.O (g6682), .I (I11994));
INVX1 gate3924(.O (g6766), .I (I12167));
INVX1 gate3925(.O (g6087), .I (I10705));
INVX1 gate3926(.O (I12173), .I (g5918));
INVX1 gate3927(.O (g8178), .I (I14413));
INVX1 gate3928(.O (g6305), .I (I11242));
INVX1 gate3929(.O (g6801), .I (I12274));
INVX1 gate3930(.O (I6856), .I (g449));
INVX1 gate3931(.O (g4590), .I (g2932));
INVX1 gate3932(.O (I10522), .I (g5243));
INVX1 gate3933(.O (I15830), .I (g9180));
INVX1 gate3934(.O (I8718), .I (g3909));
INVX1 gate3935(.O (g3501), .I (g2185));
INVX1 gate3936(.O (I9443), .I (g4564));
INVX1 gate3937(.O (g5526), .I (g5086));
INVX1 gate3938(.O (g7198), .I (I13126));
INVX1 gate3939(.O (g4657), .I (I8886));
INVX1 gate3940(.O (g7747), .I (I14112));
INVX1 gate3941(.O (g7855), .I (I14267));
INVX1 gate3942(.O (g9217), .I (I15927));
INVX1 gate3943(.O (g2873), .I (g1779));
INVX1 gate3944(.O (g1854), .I (g773));
INVX1 gate3945(.O (g2632), .I (g1576));
INVX1 gate3946(.O (I9116), .I (g4297));
INVX1 gate3947(.O (I8261), .I (g3643));
INVX1 gate3948(.O (g4556), .I (g2895));
INVX1 gate3949(.O (g9066), .I (I15592));
INVX1 gate3950(.O (I13653), .I (g7246));
INVX1 gate3951(.O (g5084), .I (g4477));
INVX1 gate3952(.O (g5603), .I (g4938));
INVX1 gate3953(.O (g1941), .I (I5812));
INVX1 gate3954(.O (I6474), .I (g1941));
INVX1 gate3955(.O (g2495), .I (g26));
INVX1 gate3956(.O (I8793), .I (g3923));
INVX1 gate3957(.O (I9034), .I (g4317));
INVX1 gate3958(.O (g2653), .I (I6443));
INVX1 gate3959(.O (g7241), .I (I13185));
INVX1 gate3960(.O (g6755), .I (I12138));
INVX1 gate3961(.O (g2208), .I (I5923));
INVX1 gate3962(.O (g3942), .I (I7629));
INVX1 gate3963(.O (I12760), .I (g6685));
INVX1 gate3964(.O (g5439), .I (g5058));
INVX1 gate3965(.O (g4928), .I (g4119));
INVX1 gate3966(.O (I10862), .I (g5364));
INVX1 gate3967(.O (g6226), .I (g5658));
INVX1 gate3968(.O (g4930), .I (g4121));
INVX1 gate3969(.O (g8916), .I (I15334));
INVX1 gate3970(.O (g2869), .I (g2224));
INVX1 gate3971(.O (I15610), .I (g8995));
INVX1 gate3972(.O (I15705), .I (g9068));
INVX1 gate3973(.O (I10949), .I (g5513));
INVX1 gate3974(.O (g9048), .I (I15546));
INVX1 gate3975(.O (g4899), .I (g4080));
INVX1 gate3976(.O (g4464), .I (I8486));
INVX1 gate3977(.O (I9347), .I (g3896));
INVX1 gate3978(.O (g1708), .I (I5552));
INVX1 gate3979(.O (I9681), .I (g4811));
INVX1 gate3980(.O (g7524), .I (I13752));
INVX1 gate3981(.O (g6173), .I (I10882));
INVX1 gate3982(.O (g2752), .I (g2389));
INVX1 gate3983(.O (g3954), .I (I7655));
INVX1 gate3984(.O (g6373), .I (I11446));
INVX1 gate3985(.O (I10702), .I (g5529));
INVX1 gate3986(.O (I15678), .I (g9060));
INVX1 gate3987(.O (g9133), .I (I15773));
INVX1 gate3988(.O (g2917), .I (g2309));
INVX1 gate3989(.O (g9333), .I (g9323));
INVX1 gate3990(.O (g7119), .I (I12945));
INVX1 gate3991(.O (g1812), .I (I5682));
INVX1 gate3992(.O (g7319), .I (g7124));
INVX1 gate3993(.O (I14904), .I (g8629));
INVX1 gate3994(.O (I8721), .I (g3918));
INVX1 gate3995(.O (g1958), .I (g786));
INVX1 gate3996(.O (g2265), .I (I6000));
INVX1 gate3997(.O (g6369), .I (I11434));
INVX1 gate3998(.O (g7352), .I (I13472));
INVX1 gate3999(.O (g7577), .I (I13876));
INVX1 gate4000(.O (g6007), .I (g5494));
INVX1 gate4001(.O (I12927), .I (g7014));
INVX1 gate4002(.O (g9196), .I (g9185));
INVX1 gate4003(.O (g7717), .I (I14028));
INVX1 gate4004(.O (g6059), .I (g5317));
INVX1 gate4005(.O (g6868), .I (I12475));
INVX1 gate4006(.O (g5616), .I (g4938));
INVX1 gate4007(.O (g3568), .I (g1935));
INVX1 gate4008(.O (g8873), .I (I15205));
INVX1 gate4009(.O (I13484), .I (g7128));
INVX1 gate4010(.O (g1829), .I (I5715));
INVX1 gate4011(.O (g8632), .I (I14712));
INVX1 gate4012(.O (I5842), .I (g68));
INVX1 gate4013(.O (I15065), .I (g8636));
INVX1 gate4014(.O (g6767), .I (I12170));
INVX1 gate4015(.O (g2364), .I (I6192));
INVX1 gate4016(.O (I12649), .I (g6457));
INVX1 gate4017(.O (g2233), .I (I5960));
INVX1 gate4018(.O (I10183), .I (g5129));
INVX1 gate4019(.O (g1911), .I (I5789));
INVX1 gate4020(.O (I10397), .I (g5200));
INVX1 gate4021(.O (g7211), .I (I13147));
INVX1 gate4022(.O (I5392), .I (g694));
INVX1 gate4023(.O (g3912), .I (g3192));
INVX1 gate4024(.O (I14397), .I (g7686));
INVX1 gate4025(.O (g4089), .I (I7888));
INVX1 gate4026(.O (I12903), .I (g6905));
INVX1 gate4027(.O (g2454), .I (I6294));
INVX1 gate4028(.O (I11200), .I (g6251));
INVX1 gate4029(.O (g8869), .I (I15193));
INVX1 gate4030(.O (g4489), .I (g2826));
INVX1 gate4031(.O (g2770), .I (g2210));
INVX1 gate4032(.O (g6793), .I (I12250));
INVX1 gate4033(.O (I10509), .I (g5237));
INVX1 gate4034(.O (g9018), .I (I15478));
INVX1 gate4035(.O (g4557), .I (g2896));
INVX1 gate4036(.O (g5764), .I (I10369));
INVX1 gate4037(.O (g7599), .I (g7450));
INVX1 gate4038(.O (g9067), .I (I15595));
INVX1 gate4039(.O (g1974), .I (g803));
INVX1 gate4040(.O (I10933), .I (g5668));
INVX1 gate4041(.O (g7274), .I (I13258));
INVX1 gate4042(.O (I15218), .I (g8801));
INVX1 gate4043(.O (g6015), .I (I10617));
INVX1 gate4044(.O (g4071), .I (I7850));
INVX1 gate4045(.O (I6000), .I (g202));
INVX1 gate4046(.O (I7341), .I (g2931));
INVX1 gate4047(.O (g2532), .I (I6358));
INVX1 gate4048(.O (g8752), .I (g8564));
INVX1 gate4049(.O (g6227), .I (I11018));
INVX1 gate4050(.O (g3929), .I (I7588));
INVX1 gate4051(.O (I13921), .I (g7362));
INVX1 gate4052(.O (I6326), .I (g1443));
INVX1 gate4053(.O (I14851), .I (g8630));
INVX1 gate4054(.O (g8917), .I (I15337));
INVX1 gate4055(.O (g1796), .I (g617));
INVX1 gate4056(.O (g4242), .I (I8161));
INVX1 gate4057(.O (g7125), .I (I12965));
INVX1 gate4058(.O (g9093), .I (I15669));
INVX1 gate4059(.O (I8428), .I (g3611));
INVX1 gate4060(.O (g6246), .I (I11055));
INVX1 gate4061(.O (I7691), .I (g3651));
INVX1 gate4062(.O (I15160), .I (g8631));
INVX1 gate4063(.O (I13813), .I (g7314));
INVX1 gate4064(.O (g8042), .I (I14325));
INVX1 gate4065(.O (g5224), .I (g5114));
INVX1 gate4066(.O (g7280), .I (I13274));
INVX1 gate4067(.O (g8442), .I (I14623));
INVX1 gate4068(.O (g6721), .I (g6257));
INVX1 gate4069(.O (g8786), .I (g8545));
INVX1 gate4070(.O (g5120), .I (I9512));
INVX1 gate4071(.O (I12262), .I (g6656));
INVX1 gate4072(.O (g2389), .I (g1230));
INVX1 gate4073(.O (g9181), .I (g9177));
INVX1 gate4074(.O (g2706), .I (g1821));
INVX1 gate4075(.O (g7544), .I (I13816));
INVX1 gate4076(.O (I8826), .I (g4023));
INVX1 gate4077(.O (g9381), .I (I16165));
INVX1 gate4078(.O (I5812), .I (g1243));
INVX1 gate4079(.O (g7483), .I (g7226));
INVX1 gate4080(.O (I15915), .I (g9194));
INVX1 gate4081(.O (I9460), .I (g3941));
INVX1 gate4082(.O (I9597), .I (g4738));
INVX1 gate4083(.O (I6183), .I (g6));
INVX1 gate4084(.O (g4350), .I (I8315));
INVX1 gate4085(.O (g2888), .I (I6608));
INVX1 gate4086(.O (I6608), .I (g1612));
INVX1 gate4087(.O (g9197), .I (g9186));
INVX1 gate4088(.O (I6220), .I (g126));
INVX1 gate4089(.O (I10574), .I (g5426));
INVX1 gate4090(.O (g2371), .I (g944));
INVX1 gate4091(.O (I8910), .I (g4200));
INVX1 gate4092(.O (g2787), .I (g1807));
INVX1 gate4093(.O (g4438), .I (I8446));
INVX1 gate4094(.O (g7106), .I (I12906));
INVX1 gate4095(.O (I11732), .I (g6076));
INVX1 gate4096(.O (g5617), .I (g4969));
INVX1 gate4097(.O (g8770), .I (g8545));
INVX1 gate4098(.O (g6502), .I (I11672));
INVX1 gate4099(.O (I14205), .I (g7710));
INVX1 gate4100(.O (g7306), .I (I13350));
INVX1 gate4101(.O (g5789), .I (I10412));
INVX1 gate4102(.O (g4009), .I (I7758));
INVX1 gate4103(.O (g2956), .I (g2375));
INVX1 gate4104(.O (I16119), .I (g9351));
INVX1 gate4105(.O (I14311), .I (g7566));
INVX1 gate4106(.O (g7790), .I (I14227));
INVX1 gate4107(.O (g5516), .I (g4924));
INVX1 gate4108(.O (I15595), .I (g8990));
INVX1 gate4109(.O (g6940), .I (I12639));
INVX1 gate4110(.O (I5911), .I (g216));
INVX1 gate4111(.O (I8308), .I (g3674));
INVX1 gate4112(.O (g7061), .I (g6650));
INVX1 gate4113(.O (g7187), .I (I13103));
INVX1 gate4114(.O (I7311), .I (g2879));
INVX1 gate4115(.O (g5987), .I (g5294));
INVX1 gate4116(.O (g1849), .I (I5732));
INVX1 gate4117(.O (g3778), .I (g2145));
INVX1 gate4118(.O (I13692), .I (g7343));
INVX1 gate4119(.O (I13761), .I (g7418));
INVX1 gate4120(.O (g642), .I (I5377));
INVX1 gate4121(.O (I8883), .I (g4198));
INVX1 gate4122(.O (g7756), .I (I14139));
INVX1 gate4123(.O (g6388), .I (I11491));
INVX1 gate4124(.O (I10592), .I (g5444));
INVX1 gate4125(.O (g5299), .I (I9804));
INVX1 gate4126(.O (I9840), .I (g4702));
INVX1 gate4127(.O (g3735), .I (g1961));
INVX1 gate4128(.O (g4918), .I (g4103));
INVX1 gate4129(.O (g6216), .I (I10987));
INVX1 gate4130(.O (g1781), .I (g622));
INVX1 gate4131(.O (I6051), .I (g440));
INVX1 gate4132(.O (I7374), .I (g3084));
INVX1 gate4133(.O (I10780), .I (g5445));
INVX1 gate4134(.O (g8012), .I (I14305));
INVX1 gate4135(.O (I6127), .I (g471));
INVX1 gate4136(.O (I6451), .I (g1895));
INVX1 gate4137(.O (g6028), .I (g5529));
INVX1 gate4138(.O (I14780), .I (g8284));
INVX1 gate4139(.O (I12247), .I (g6646));
INVX1 gate4140(.O (g6671), .I (I11971));
INVX1 gate4141(.O (g7904), .I (I14276));
INVX1 gate4142(.O (g1797), .I (g627));
INVX1 gate4143(.O (g2639), .I (g1583));
INVX1 gate4144(.O (g7046), .I (I12806));
INVX1 gate4145(.O (I11329), .I (g5825));
INVX1 gate4146(.O (g3075), .I (g2216));
INVX1 gate4147(.O (g2963), .I (g2383));
INVX1 gate4148(.O (g4229), .I (I8140));
INVX1 gate4149(.O (I10350), .I (g5707));
INVX1 gate4150(.O (I13329), .I (g7247));
INVX1 gate4151(.O (g7446), .I (I13595));
INVX1 gate4152(.O (g7514), .I (I13722));
INVX1 gate4153(.O (g3949), .I (I7644));
INVX1 gate4154(.O (g2309), .I (I6084));
INVX1 gate4155(.O (g9101), .I (I15693));
INVX1 gate4156(.O (I7545), .I (g3589));
INVX1 gate4157(.O (I12388), .I (g6403));
INVX1 gate4158(.O (g9301), .I (g9260));
INVX1 gate4159(.O (g4822), .I (I9177));
INVX1 gate4160(.O (g7145), .I (I13023));
INVX1 gate4161(.O (g8029), .I (I14318));
INVX1 gate4162(.O (I7380), .I (g3461));
INVX1 gate4163(.O (g7345), .I (I13451));
INVX1 gate4164(.O (I12098), .I (g5956));
INVX1 gate4165(.O (g8787), .I (g8564));
INVX1 gate4166(.O (I16036), .I (g9282));
INVX1 gate4167(.O (I7832), .I (g2768));
INVX1 gate4168(.O (g5738), .I (I10271));
INVX1 gate4169(.O (g6826), .I (I12349));
INVX1 gate4170(.O (g7763), .I (I14160));
INVX1 gate4171(.O (g3526), .I (g2185));
INVX1 gate4172(.O (g8956), .I (I15382));
INVX1 gate4173(.O (g3998), .I (g3097));
INVX1 gate4174(.O (g8675), .I (I14819));
INVX1 gate4175(.O (g5709), .I (g4841));
INVX1 gate4176(.O (I8333), .I (g3721));
INVX1 gate4177(.O (g6741), .I (I12117));
INVX1 gate4178(.O (I15589), .I (g8988));
INVX1 gate4179(.O (g3084), .I (I6820));
INVX1 gate4180(.O (g3603), .I (g2092));
INVX1 gate4181(.O (I5377), .I (g635));
INVX1 gate4182(.O (g785), .I (I5407));
INVX1 gate4183(.O (g5478), .I (g5025));
INVX1 gate4184(.O (I13241), .I (g7030));
INVX1 gate4185(.O (I14413), .I (g7723));
INVX1 gate4186(.O (g1694), .I (g21));
INVX1 gate4187(.O (g7107), .I (I12909));
INVX1 gate4188(.O (g4921), .I (g4202));
INVX1 gate4189(.O (g7307), .I (I13353));
INVX1 gate4190(.O (g3850), .I (I7353));
INVX1 gate4191(.O (I15836), .I (g9165));
INVX1 gate4192(.O (g2957), .I (g2376));
INVX1 gate4193(.O (I8196), .I (g3654));
INVX1 gate4194(.O (g7159), .I (I13051));
INVX1 gate4195(.O (I7931), .I (g2780));
INVX1 gate4196(.O (g1852), .I (g887));
INVX1 gate4197(.O (g1923), .I (I5801));
INVX1 gate4198(.O (I6072), .I (g1211));
INVX1 gate4199(.O (g6108), .I (g5345));
INVX1 gate4200(.O (g7359), .I (I13493));
INVX1 gate4201(.O (I9250), .I (g4134));
INVX1 gate4202(.O (g5435), .I (g5121));
INVX1 gate4203(.O (g6308), .I (I11251));
INVX1 gate4204(.O (g5517), .I (g4925));
INVX1 gate4205(.O (g5690), .I (g4748));
INVX1 gate4206(.O (I9363), .I (g4258));
INVX1 gate4207(.O (g7223), .I (I13161));
INVX1 gate4208(.O (g5482), .I (g4915));
INVX1 gate4209(.O (g1701), .I (I5545));
INVX1 gate4210(.O (g6883), .I (I12520));
INVX1 gate4211(.O (I9053), .I (g4327));
INVX1 gate4212(.O (g8684), .I (I14848));
INVX1 gate4213(.O (g3583), .I (g2128));
INVX1 gate4214(.O (g4895), .I (g4078));
INVX1 gate4215(.O (g8639), .I (I14725));
INVX1 gate4216(.O (I6443), .I (g1774));
INVX1 gate4217(.O (g7757), .I (I14142));
INVX1 gate4218(.O (I7905), .I (g2863));
INVX1 gate4219(.O (I11683), .I (g5988));
INVX1 gate4220(.O (g4620), .I (I8775));
INVX1 gate4221(.O (g8791), .I (g8585));
INVX1 gate4222(.O (g4462), .I (I8480));
INVX1 gate4223(.O (g2498), .I (I6333));
INVX1 gate4224(.O (g6217), .I (g5649));
INVX1 gate4225(.O (g3919), .I (I7554));
INVX1 gate4226(.O (g6758), .I (I12145));
INVX1 gate4227(.O (g6589), .I (g6083));
INVX1 gate4228(.O (g1886), .I (I5766));
INVX1 gate4229(.O (I7204), .I (g2520));
INVX1 gate4230(.O (I16009), .I (g9261));
INVX1 gate4231(.O (I15616), .I (g8997));
INVX1 gate4232(.O (I5781), .I (g979));
INVX1 gate4233(.O (g2833), .I (I6561));
INVX1 gate4234(.O (g7522), .I (I13746));
INVX1 gate4235(.O (g7115), .I (I12933));
INVX1 gate4236(.O (g7251), .I (I13203));
INVX1 gate4237(.O (g8808), .I (I15062));
INVX1 gate4238(.O (I6434), .I (g1830));
INVX1 gate4239(.O (g3952), .I (I7651));
INVX1 gate4240(.O (g7315), .I (I13373));
INVX1 gate4241(.O (g7811), .I (I14238));
INVX1 gate4242(.O (g7047), .I (g6498));
INVX1 gate4243(.O (g9368), .I (I16132));
INVX1 gate4244(.O (I8994), .I (g4565));
INVX1 gate4245(.O (I10046), .I (g4840));
INVX1 gate4246(.O (g6861), .I (I12454));
INVX1 gate4247(.O (g6365), .I (I11422));
INVX1 gate4248(.O (g2584), .I (g1646));
INVX1 gate4249(.O (I14046), .I (g7492));
INVX1 gate4250(.O (g4788), .I (I9103));
INVX1 gate4251(.O (g6048), .I (g5246));
INVX1 gate4252(.O (I11515), .I (g5897));
INVX1 gate4253(.O (I11991), .I (g5939));
INVX1 gate4254(.O (g2539), .I (I6363));
INVX1 gate4255(.O (g2896), .I (g2269));
INVX1 gate4256(.O (g3561), .I (I7041));
INVX1 gate4257(.O (g9058), .I (I15568));
INVX1 gate4258(.O (I13515), .I (g7152));
INVX1 gate4259(.O (g8759), .I (g8524));
INVX1 gate4260(.O (I13882), .I (g7350));
INVX1 gate4261(.O (g6711), .I (I12059));
INVX1 gate4262(.O (g1870), .I (I5751));
INVX1 gate4263(.O (I11407), .I (g5841));
INVX1 gate4264(.O (I13407), .I (g7271));
INVX1 gate4265(.O (g1825), .I (I5709));
INVX1 gate4266(.O (g6827), .I (I12352));
INVX1 gate4267(.O (g3527), .I (g1616));
INVX1 gate4268(.O (g8957), .I (I15385));
INVX1 gate4269(.O (g6133), .I (I10766));
INVX1 gate4270(.O (g6333), .I (I11326));
INVX1 gate4271(.O (I14282), .I (g7709));
INVX1 gate4272(.O (g3647), .I (g2424));
INVX1 gate4273(.O (I9929), .I (g5052));
INVX1 gate4274(.O (g2162), .I (I5901));
INVX1 gate4275(.O (I7973), .I (g3071));
INVX1 gate4276(.O (g2268), .I (I6009));
INVX1 gate4277(.O (g6774), .I (I12193));
INVX1 gate4278(.O (g2362), .I (I6186));
INVX1 gate4279(.O (I12629), .I (g6523));
INVX1 gate4280(.O (g3764), .I (g2039));
INVX1 gate4281(.O (g4085), .I (I7878));
INVX1 gate4282(.O (I12451), .I (g6524));
INVX1 gate4283(.O (g6846), .I (I12409));
INVX1 gate4284(.O (I12472), .I (g6591));
INVX1 gate4285(.O (I12220), .I (g6645));
INVX1 gate4286(.O (g8865), .I (I15181));
INVX1 gate4287(.O (g3546), .I (I7029));
INVX1 gate4288(.O (g5002), .I (g4335));
INVX1 gate4289(.O (I14743), .I (g8174));
INVX1 gate4290(.O (I8847), .I (g4025));
INVX1 gate4291(.O (g2052), .I (I5865));
INVX1 gate4292(.O (g5402), .I (g5000));
INVX1 gate4293(.O (g5824), .I (I10497));
INVX1 gate4294(.O (g7595), .I (I13930));
INVX1 gate4295(.O (g6803), .I (I12280));
INVX1 gate4296(.O (g2452), .I (g23));
INVX1 gate4297(.O (g8604), .I (I14677));
INVX1 gate4298(.O (g3503), .I (g2407));
INVX1 gate4299(.O (g3970), .I (g2845));
INVX1 gate4300(.O (g1768), .I (g605));
INVX1 gate4301(.O (g9074), .I (I15616));
INVX1 gate4302(.O (g6538), .I (I11714));
INVX1 gate4303(.O (I13441), .I (g7146));
INVX1 gate4304(.O (I5852), .I (g1202));
INVX1 gate4305(.O (I5923), .I (g252));
INVX1 gate4306(.O (I11206), .I (g6133));
INVX1 gate4307(.O (I7323), .I (g2905));
INVX1 gate4308(.O (g6780), .I (I12211));
INVX1 gate4309(.O (g6509), .I (I11689));
INVX1 gate4310(.O (g1806), .I (I5670));
INVX1 gate4311(.O (g1943), .I (g1025));
INVX1 gate4312(.O (I6820), .I (g1707));
INVX1 gate4313(.O (g7243), .I (I13189));
INVX1 gate4314(.O (I6936), .I (g1878));
INVX1 gate4315(.O (I11725), .I (g6036));
INVX1 gate4316(.O (I12776), .I (g6739));
INVX1 gate4317(.O (I13725), .I (g7437));
INVX1 gate4318(.O (g2728), .I (g2256));
INVX1 gate4319(.O (g2486), .I (g959));
INVX1 gate4320(.O (g6662), .I (I11964));
INVX1 gate4321(.O (g6018), .I (g5494));
INVX1 gate4322(.O (I6317), .I (g1339));
INVX1 gate4323(.O (g1887), .I (g83));
INVX1 gate4324(.O (I16176), .I (g9385));
INVX1 gate4325(.O (I13758), .I (g7414));
INVX1 gate4326(.O (I15693), .I (g9048));
INVX1 gate4327(.O (I12355), .I (g6756));
INVX1 gate4328(.O (I13435), .I (g7170));
INVX1 gate4329(.O (g1934), .I (g154));
INVX1 gate4330(.O (g2185), .I (I5914));
INVX1 gate4331(.O (g6290), .I (I11197));
INVX1 gate4332(.O (g4640), .I (I8835));
INVX1 gate4333(.O (g2881), .I (g2235));
INVX1 gate4334(.O (I7648), .I (g2712));
INVX1 gate4335(.O (I16154), .I (g9370));
INVX1 gate4336(.O (I7875), .I (g3819));
INVX1 gate4337(.O (I12370), .I (g6758));
INVX1 gate4338(.O (g4031), .I (I7804));
INVX1 gate4339(.O (g7130), .I (I12976));
INVX1 gate4340(.O (I7655), .I (g2734));
INVX1 gate4341(.O (g3617), .I (g1655));
INVX1 gate4342(.O (g6093), .I (g5345));
INVX1 gate4343(.O (I11744), .I (g6120));
INVX1 gate4344(.O (g7542), .I (I13810));
INVX1 gate4345(.O (g2470), .I (g42));
INVX1 gate4346(.O (g7330), .I (I13410));
INVX1 gate4347(.O (g2897), .I (g2270));
INVX1 gate4348(.O (g6493), .I (I11659));
INVX1 gate4349(.O (g6256), .I (I11069));
INVX1 gate4350(.O (I12151), .I (g5847));
INVX1 gate4351(.O (g6816), .I (I12319));
INVX1 gate4352(.O (g5785), .I (I10400));
INVX1 gate4353(.O (I12996), .I (g6934));
INVX1 gate4354(.O (g4005), .I (I7746));
INVX1 gate4355(.O (I13940), .I (g7355));
INVX1 gate4356(.O (I8101), .I (g3259));
INVX1 gate4357(.O (I8817), .I (g3935));
INVX1 gate4358(.O (I14662), .I (g7783));
INVX1 gate4359(.O (g3987), .I (I7716));
INVX1 gate4360(.O (g3771), .I (g1853));
INVX1 gate4361(.O (I11848), .I (g6159));
INVX1 gate4362(.O (I9782), .I (g4720));
INVX1 gate4363(.O (I11398), .I (g5823));
INVX1 gate4364(.O (I12367), .I (g6754));
INVX1 gate4365(.O (I12394), .I (g6759));
INVX1 gate4366(.O (I6060), .I (g580));
INVX1 gate4367(.O (g6381), .I (I11470));
INVX1 gate4368(.O (g4286), .I (g3790));
INVX1 gate4369(.O (I11652), .I (g5939));
INVX1 gate4370(.O (g6847), .I (I12412));
INVX1 gate4371(.O (I6460), .I (g2104));
INVX1 gate4372(.O (I6597), .I (g1970));
INVX1 gate4373(.O (I10482), .I (g5228));
INVX1 gate4374(.O (g3547), .I (g2345));
INVX1 gate4375(.O (g6700), .I (g6244));
INVX1 gate4376(.O (g6397), .I (I11512));
INVX1 gate4377(.O (I10552), .I (g5396));
INVX1 gate4378(.O (I8751), .I (g4009));
INVX1 gate4379(.O (g3892), .I (g3131));
INVX1 gate4380(.O (I11263), .I (g5784));
INVX1 gate4381(.O (I10204), .I (g5060));
INVX1 gate4382(.O (I9627), .I (g4777));
INVX1 gate4383(.O (g2131), .I (g1300));
INVX1 gate4384(.O (I6784), .I (g2052));
INVX1 gate4385(.O (g2006), .I (g806));
INVX1 gate4386(.O (g2331), .I (g933));
INVX1 gate4387(.O (I12319), .I (g6741));
INVX1 gate4388(.O (g4733), .I (g4202));
INVX1 gate4389(.O (I11332), .I (g5832));
INVX1 gate4390(.O (g5844), .I (I10545));
INVX1 gate4391(.O (I13332), .I (g7241));
INVX1 gate4392(.O (g6263), .I (g5688));
INVX1 gate4393(.O (g4270), .I (g2573));
INVX1 gate4394(.O (I5972), .I (g356));
INVX1 gate4395(.O (g2635), .I (g1579));
INVX1 gate4396(.O (g1807), .I (g619));
INVX1 gate4397(.O (g6950), .I (I12659));
INVX1 gate4398(.O (g8881), .I (g8683));
INVX1 gate4399(.O (g9126), .I (I15756));
INVX1 gate4400(.O (g4610), .I (I8745));
INVX1 gate4401(.O (g2105), .I (g1444));
INVX1 gate4402(.O (I7667), .I (g3052));
INVX1 gate4403(.O (g3945), .I (g3097));
INVX1 gate4404(.O (I12059), .I (g5874));
INVX1 gate4405(.O (I10786), .I (g5452));
INVX1 gate4406(.O (I12025), .I (g5918));
INVX1 gate4407(.O (g2487), .I (I6323));
INVX1 gate4408(.O (I9084), .I (g4358));
INVX1 gate4409(.O (g5731), .I (I10250));
INVX1 gate4410(.O (I9603), .I (g4719));
INVX1 gate4411(.O (I13962), .I (g7413));
INVX1 gate4412(.O (I14786), .I (g8606));
INVX1 gate4413(.O (g7512), .I (I13716));
INVX1 gate4414(.O (I9484), .I (g3957));
INVX1 gate4415(.O (g3991), .I (g3160));
INVX1 gate4416(.O (g7090), .I (g6525));
INVX1 gate4417(.O (I6294), .I (g1330));
INVX1 gate4418(.O (I9850), .I (g4798));
INVX1 gate4419(.O (g594), .I (I5368));
INVX1 gate4420(.O (I10356), .I (g5711));
INVX1 gate4421(.O (I15382), .I (g8883));
INVX1 gate4422(.O (I11500), .I (g6219));
INVX1 gate4423(.O (g6562), .I (I11736));
INVX1 gate4424(.O (g7366), .I (I13512));
INVX1 gate4425(.O (g4069), .I (I7844));
INVX1 gate4426(.O (I15519), .I (g9019));
INVX1 gate4427(.O (g5071), .I (g4438));
INVX1 gate4428(.O (g3078), .I (g1603));
INVX1 gate4429(.O (g3340), .I (g2474));
INVX1 gate4430(.O (I10826), .I (g5434));
INVX1 gate4431(.O (I15675), .I (g9058));
INVX1 gate4432(.O (I10380), .I (g5448));
INVX1 gate4433(.O (g5705), .I (g4841));
INVX1 gate4434(.O (g5471), .I (I9889));
INVX1 gate4435(.O (g7056), .I (g6520));
INVX1 gate4436(.O (g6631), .I (I11887));
INVX1 gate4437(.O (g4540), .I (g2882));
INVX1 gate4438(.O (g2226), .I (g1320));
INVX1 gate4439(.O (I7548), .I (g3590));
INVX1 gate4440(.O (I10998), .I (g5672));
INVX1 gate4441(.O (I12044), .I (g5847));
INVX1 gate4442(.O (g6723), .I (I12085));
INVX1 gate4443(.O (g7456), .I (g7174));
INVX1 gate4444(.O (I13048), .I (g6956));
INVX1 gate4445(.O (g7529), .I (I13767));
INVX1 gate4446(.O (g6257), .I (g5685));
INVX1 gate4447(.O (g3959), .I (g3097));
INVX1 gate4448(.O (g1815), .I (g760));
INVX1 gate4449(.O (g6101), .I (g5317));
INVX1 gate4450(.O (g7148), .I (I13028));
INVX1 gate4451(.O (g6817), .I (I12322));
INVX1 gate4452(.O (g9183), .I (g9161));
INVX1 gate4453(.O (g6301), .I (I11230));
INVX1 gate4454(.O (g7348), .I (I13460));
INVX1 gate4455(.O (g3517), .I (g2283));
INVX1 gate4456(.O (I11004), .I (g5613));
INVX1 gate4457(.O (g3082), .I (g1680));
INVX1 gate4458(.O (g9383), .I (g9380));
INVX1 gate4459(.O (I8772), .I (g4011));
INVX1 gate4460(.O (I7804), .I (g3029));
INVX1 gate4461(.O (g9220), .I (g9205));
INVX1 gate4462(.O (I11221), .I (g6167));
INVX1 gate4463(.O (g7155), .I (I13039));
INVX1 gate4464(.O (g7355), .I (I13481));
INVX1 gate4465(.O (g6605), .I (I11821));
INVX1 gate4466(.O (I7792), .I (g3038));
INVX1 gate4467(.O (I12301), .I (g6703));
INVX1 gate4468(.O (g8678), .I (I14828));
INVX1 gate4469(.O (g1726), .I (g158));
INVX1 gate4470(.O (g3876), .I (g3466));
INVX1 gate4471(.O (g8131), .I (I14378));
INVX1 gate4472(.O (I12120), .I (g5939));
INVX1 gate4473(.O (g2373), .I (I6217));
INVX1 gate4474(.O (g2091), .I (g819));
INVX1 gate4475(.O (g8406), .I (I14614));
INVX1 gate4476(.O (I13613), .I (g7273));
INVX1 gate4477(.O (g1960), .I (g1268));
INVX1 gate4478(.O (g5814), .I (I10475));
INVX1 gate4479(.O (g7260), .I (g7064));
INVX1 gate4480(.O (g6751), .I (I12128));
INVX1 gate4481(.O (g5150), .I (I9576));
INVX1 gate4482(.O (I8011), .I (g3225));
INVX1 gate4483(.O (I9561), .I (g4695));
INVX1 gate4484(.O (g8682), .I (I14844));
INVX1 gate4485(.O (g8766), .I (g8545));
INVX1 gate4486(.O (g5038), .I (g4457));
INVX1 gate4487(.O (I5395), .I (g698));
INVX1 gate4488(.O (I8856), .I (g3955));
INVX1 gate4489(.O (g2283), .I (I6033));
INVX1 gate4490(.O (g7063), .I (I12826));
INVX1 gate4491(.O (I12699), .I (g6504));
INVX1 gate4492(.O (g9161), .I (I15803));
INVX1 gate4493(.O (I16138), .I (g9358));
INVX1 gate4494(.O (I13106), .I (g7056));
INVX1 gate4495(.O (g9361), .I (I16119));
INVX1 gate4496(.O (g2007), .I (g1223));
INVX1 gate4497(.O (I13605), .I (g7197));
INVX1 gate4498(.O (I10448), .I (g5335));
INVX1 gate4499(.O (g7463), .I (g7239));
INVX1 gate4500(.O (g5009), .I (g4344));
INVX1 gate4501(.O (g2407), .I (I6286));
INVX1 gate4502(.O (I6163), .I (g402));
INVX1 gate4503(.O (I14448), .I (g7792));
INVX1 gate4504(.O (g2920), .I (I6652));
INVX1 gate4505(.O (g2868), .I (g2223));
INVX1 gate4506(.O (I6363), .I (g16));
INVX1 gate4507(.O (I15501), .I (g8975));
INVX1 gate4508(.O (g9051), .I (I15553));
INVX1 gate4509(.O (I15729), .I (g9073));
INVX1 gate4510(.O (g2459), .I (I6299));
INVX1 gate4511(.O (I15577), .I (g8984));
INVX1 gate4512(.O (g4898), .I (g4079));
INVX1 gate4513(.O (g6441), .I (I11586));
INVX1 gate4514(.O (I13463), .I (g7264));
INVX1 gate4515(.O (g9127), .I (I15759));
INVX1 gate4516(.O (g2767), .I (I6509));
INVX1 gate4517(.O (g4900), .I (I9258));
INVX1 gate4518(.O (g1783), .I (I5633));
INVX1 gate4519(.O (I7908), .I (g3516));
INVX1 gate4520(.O (g5769), .I (I10380));
INVX1 gate4521(.O (I11951), .I (g5847));
INVX1 gate4522(.O (I11371), .I (g5840));
INVX1 gate4523(.O (g8755), .I (g8545));
INVX1 gate4524(.O (g636), .I (I5371));
INVX1 gate4525(.O (g7279), .I (I13271));
INVX1 gate4526(.O (g8226), .I (I14457));
INVX1 gate4527(.O (g5836), .I (g5529));
INVX1 gate4528(.O (g4510), .I (g2840));
INVX1 gate4529(.O (I13234), .I (g6898));
INVX1 gate4530(.O (g4245), .I (I8172));
INVX1 gate4531(.O (I12427), .I (g6553));
INVX1 gate4532(.O (g7720), .I (I14035));
INVX1 gate4533(.O (g7118), .I (I12942));
INVX1 gate4534(.O (g5918), .I (I10574));
INVX1 gate4535(.O (g2793), .I (I6532));
INVX1 gate4536(.O (g7367), .I (I13515));
INVX1 gate4537(.O (I12632), .I (g6514));
INVX1 gate4538(.O (g9103), .I (I15699));
INVX1 gate4539(.O (g9303), .I (g9301));
INVX1 gate4540(.O (g1676), .I (g727));
INVX1 gate4541(.O (g2015), .I (g33));
INVX1 gate4542(.O (I8480), .I (g3640));
INVX1 gate4543(.O (g6368), .I (I11431));
INVX1 gate4544(.O (g7057), .I (g6644));
INVX1 gate4545(.O (g8173), .I (I14400));
INVX1 gate4546(.O (g4344), .I (g3124));
INVX1 gate4547(.O (g6772), .I (I12187));
INVX1 gate4548(.O (I6157), .I (g246));
INVX1 gate4549(.O (I12403), .I (g6769));
INVX1 gate4550(.O (I12547), .I (g6708));
INVX1 gate4551(.O (g1828), .I (g769));
INVX1 gate4552(.O (g2664), .I (I6463));
INVX1 gate4553(.O (g2246), .I (I5989));
INVX1 gate4554(.O (g4259), .I (I8196));
INVX1 gate4555(.O (g5822), .I (I10491));
INVX1 gate4556(.O (g6890), .I (I12541));
INVX1 gate4557(.O (g7549), .I (I13831));
INVX1 gate4558(.O (g1830), .I (I5718));
INVX1 gate4559(.O (g4694), .I (I8977));
INVX1 gate4560(.O (I15622), .I (g8999));
INVX1 gate4561(.O (g1727), .I (g596));
INVX1 gate4562(.O (g3590), .I (I7064));
INVX1 gate4563(.O (g3877), .I (g2960));
INVX1 gate4564(.O (I10433), .I (g5212));
INVX1 gate4565(.O (I5692), .I (g906));
INVX1 gate4566(.O (g8602), .I (g8094));
INVX1 gate4567(.O (I10387), .I (g5194));
INVX1 gate4568(.O (I12226), .I (g6636));
INVX1 gate4569(.O (I14433), .I (g8061));
INVX1 gate4570(.O (g7686), .I (I13979));
INVX1 gate4571(.O (g8407), .I (g8013));
INVX1 gate4572(.O (g4088), .I (I7885));
INVX1 gate4573(.O (I12481), .I (g6616));
INVX1 gate4574(.O (g9072), .I (I15610));
INVX1 gate4575(.O (g3657), .I (I7145));
INVX1 gate4576(.O (g4923), .I (g4112));
INVX1 gate4577(.O (g2721), .I (g1803));
INVX1 gate4578(.O (g6505), .I (I11677));
INVX1 gate4579(.O (g8868), .I (I15190));
INVX1 gate4580(.O (I14148), .I (g7543));
INVX1 gate4581(.O (g6011), .I (g5494));
INVX1 gate4582(.O (I5960), .I (g187));
INVX1 gate4583(.O (g1746), .I (g290));
INVX1 gate4584(.O (I14097), .I (g7595));
INVX1 gate4585(.O (g6856), .I (I12439));
INVX1 gate4586(.O (g4701), .I (I8994));
INVX1 gate4587(.O (I10646), .I (g5364));
INVX1 gate4588(.O (g8767), .I (g8564));
INVX1 gate4589(.O (g9043), .I (I15533));
INVX1 gate4590(.O (g3556), .I (I7036));
INVX1 gate4591(.O (I13012), .I (g7071));
INVX1 gate4592(.O (I10343), .I (g5704));
INVX1 gate4593(.O (I14646), .I (g7790));
INVX1 gate4594(.O (g3928), .I (g3097));
INVX1 gate4595(.O (I16052), .I (g9291));
INVX1 gate4596(.O (g8582), .I (g8094));
INVX1 gate4597(.O (g9116), .I (I15738));
INVX1 gate4598(.O (g6074), .I (g5317));
INVX1 gate4599(.O (g3930), .I (g3097));
INVX1 gate4600(.O (g2502), .I (I6337));
INVX1 gate4601(.O (g9316), .I (g9302));
INVX1 gate4602(.O (I11473), .I (g6069));
INVX1 gate4603(.O (I13541), .I (g7209));
INVX1 gate4604(.O (g4886), .I (g4071));
INVX1 gate4605(.O (I10369), .I (g5716));
INVX1 gate4606(.O (g9034), .I (I15516));
INVX1 gate4607(.O (I12490), .I (g6625));
INVX1 gate4608(.O (g8015), .I (g7689));
INVX1 gate4609(.O (g2940), .I (I6686));
INVX1 gate4610(.O (g8227), .I (I14460));
INVX1 gate4611(.O (g4114), .I (I7953));
INVX1 gate4612(.O (g7253), .I (g7049));
INVX1 gate4613(.O (I11359), .I (g5810));
INVX1 gate4614(.O (I12376), .I (g6766));
INVX1 gate4615(.O (I12385), .I (g6397));
INVX1 gate4616(.O (I13359), .I (g7255));
INVX1 gate4617(.O (I9892), .I (g4879));
INVX1 gate4618(.O (g5462), .I (g4886));
INVX1 gate4619(.O (g2689), .I (g1670));
INVX1 gate4620(.O (g6573), .I (g5868));
INVX1 gate4621(.O (g6863), .I (I12460));
INVX1 gate4622(.O (I11920), .I (g5874));
INVX1 gate4623(.O (I12980), .I (g6929));
INVX1 gate4624(.O (I7878), .I (g2829));
INVX1 gate4625(.O (g8664), .I (I14786));
INVX1 gate4626(.O (I8760), .I (g3931));
INVX1 gate4627(.O (I11434), .I (g5789));
INVX1 gate4628(.O (g3563), .I (g2007));
INVX1 gate4629(.O (I10412), .I (g5205));
INVX1 gate4630(.O (g2216), .I (I5933));
INVX1 gate4631(.O (g6713), .I (I12065));
INVX1 gate4632(.O (g1677), .I (g1532));
INVX1 gate4633(.O (g7519), .I (I13737));
INVX1 gate4634(.O (g7740), .I (I14091));
INVX1 gate4635(.O (g4650), .I (I8865));
INVX1 gate4636(.O (I7658), .I (g2562));
INVX1 gate4637(.O (I5401), .I (g723));
INVX1 gate4638(.O (I12888), .I (g6948));
INVX1 gate4639(.O (I13828), .I (g7321));
INVX1 gate4640(.O (I5676), .I (g911));
INVX1 gate4641(.O (I14133), .I (g7574));
INVX1 gate4642(.O (g2671), .I (I6468));
INVX1 gate4643(.O (g9210), .I (g9200));
INVX1 gate4644(.O (g1576), .I (g691));
INVX1 gate4645(.O (g6569), .I (I11747));
INVX1 gate4646(.O (g1866), .I (g71));
INVX1 gate4647(.O (I7882), .I (g2700));
INVX1 gate4648(.O (g5788), .I (I10409));
INVX1 gate4649(.O (g4008), .I (I7755));
INVX1 gate4650(.O (I10896), .I (g5475));
INVX1 gate4651(.O (I6894), .I (g1863));
INVX1 gate4652(.O (I11344), .I (g5820));
INVX1 gate4653(.O (g3844), .I (I7335));
INVX1 gate4654(.O (I13344), .I (g7210));
INVX1 gate4655(.O (I15484), .I (g8918));
INVX1 gate4656(.O (g1848), .I (g772));
INVX1 gate4657(.O (I10716), .I (g5537));
INVX1 gate4658(.O (I13682), .I (g7251));
INVX1 gate4659(.O (g4594), .I (g2941));
INVX1 gate4660(.O (g5842), .I (I10541));
INVX1 gate4661(.O (g2826), .I (g2183));
INVX1 gate4662(.O (g1747), .I (g599));
INVX1 gate4663(.O (g1855), .I (g866));
INVX1 gate4664(.O (I6075), .I (g2));
INVX1 gate4665(.O (g6857), .I (I12442));
INVX1 gate4666(.O (g7586), .I (I13903));
INVX1 gate4667(.O (I9907), .I (g4837));
INVX1 gate4668(.O (I13173), .I (g7089));
INVX1 gate4669(.O (g5192), .I (g4841));
INVX1 gate4670(.O (I10582), .I (g5437));
INVX1 gate4671(.O (g3557), .I (g1773));
INVX1 gate4672(.O (g5085), .I (I9457));
INVX1 gate4673(.O (g4806), .I (I9139));
INVX1 gate4674(.O (I7981), .I (g3555));
INVX1 gate4675(.O (I6949), .I (g2148));
INVX1 gate4676(.O (I12190), .I (g5918));
INVX1 gate4677(.O (g3966), .I (g3160));
INVX1 gate4678(.O (I8977), .I (g3877));
INVX1 gate4679(.O (g2910), .I (I6636));
INVX1 gate4680(.O (g3071), .I (g1948));
INVX1 gate4681(.O (g3705), .I (I7204));
INVX1 gate4682(.O (g9117), .I (I15741));
INVX1 gate4683(.O (I12520), .I (g6622));
INVX1 gate4684(.O (g2638), .I (g1582));
INVX1 gate4685(.O (g4065), .I (I7838));
INVX1 gate4686(.O (g9317), .I (g9306));
INVX1 gate4687(.O (I8161), .I (g3517));
INVX1 gate4688(.O (g8689), .I (I14857));
INVX1 gate4689(.O (g4122), .I (I7973));
INVX1 gate4690(.O (I15921), .I (g9206));
INVX1 gate4691(.O (g4465), .I (g3677));
INVX1 gate4692(.O (g7141), .I (I13009));
INVX1 gate4693(.O (I14925), .I (g8381));
INVX1 gate4694(.O (g3948), .I (g3131));
INVX1 gate4695(.O (g4934), .I (g4125));
INVX1 gate4696(.O (g7341), .I (I13441));
INVX1 gate4697(.O (g8216), .I (I14427));
INVX1 gate4698(.O (I6646), .I (g2246));
INVX1 gate4699(.O (g2308), .I (I6081));
INVX1 gate4700(.O (I7132), .I (g2554));
INVX1 gate4701(.O (I13134), .I (g7017));
INVX1 gate4702(.O (I7332), .I (g2947));
INVX1 gate4703(.O (I8665), .I (g3051));
INVX1 gate4704(.O (I12211), .I (g6502));
INVX1 gate4705(.O (I14112), .I (g7560));
INVX1 gate4706(.O (g6326), .I (I11305));
INVX1 gate4707(.O (g7525), .I (I13755));
INVX1 gate4708(.O (g7710), .I (I14009));
INVX1 gate4709(.O (g3955), .I (I7658));
INVX1 gate4710(.O (I7680), .I (g2712));
INVX1 gate4711(.O (I11506), .I (g6189));
INVX1 gate4712(.O (I14378), .I (g7691));
INVX1 gate4713(.O (g2883), .I (g2237));
INVX1 gate4714(.O (I6084), .I (g240));
INVX1 gate4715(.O (I7353), .I (g2833));
INVX1 gate4716(.O (g8671), .I (I14807));
INVX1 gate4717(.O (I11028), .I (g5642));
INVX1 gate4718(.O (I13506), .I (g7148));
INVX1 gate4719(.O (I12088), .I (g5874));
INVX1 gate4720(.O (I6039), .I (g207));
INVX1 gate4721(.O (g4033), .I (g3192));
INVX1 gate4722(.O (I13028), .I (g7087));
INVX1 gate4723(.O (g6760), .I (I12151));
INVX1 gate4724(.O (I14603), .I (g7827));
INVX1 gate4725(.O (g5520), .I (g4928));
INVX1 gate4726(.O (I15184), .I (g8684));
INVX1 gate4727(.O (g4096), .I (I7911));
INVX1 gate4728(.O (g8564), .I (g7951));
INVX1 gate4729(.O (g3038), .I (g2092));
INVX1 gate4730(.O (g1818), .I (I5692));
INVX1 gate4731(.O (g1577), .I (g695));
INVX1 gate4732(.O (g1867), .I (g878));
INVX1 gate4733(.O (g9060), .I (I15574));
INVX1 gate4734(.O (I9310), .I (g4268));
INVX1 gate4735(.O (I7558), .I (g2734));
INVX1 gate4736(.O (I10681), .I (g5686));
INVX1 gate4737(.O (g5812), .I (I10469));
INVX1 gate4738(.O (g6183), .I (I10914));
INVX1 gate4739(.O (g7158), .I (I13048));
INVX1 gate4740(.O (g2365), .I (I6195));
INVX1 gate4741(.O (I12659), .I (g6459));
INVX1 gate4742(.O (g6383), .I (I11476));
INVX1 gate4743(.O (g7358), .I (I13490));
INVX1 gate4744(.O (g5176), .I (I9654));
INVX1 gate4745(.O (g4195), .I (I8094));
INVX1 gate4746(.O (I9663), .I (g4809));
INVX1 gate4747(.O (g6220), .I (I11001));
INVX1 gate4748(.O (g7506), .I (I13698));
INVX1 gate4749(.O (I15732), .I (g9076));
INVX1 gate4750(.O (g4891), .I (g4076));
INVX1 gate4751(.O (I13927), .I (g7366));
INVX1 gate4752(.O (g4913), .I (g4092));
INVX1 gate4753(.O (I12250), .I (g6651));
INVX1 gate4754(.O (g658), .I (I5386));
INVX1 gate4755(.O (g8910), .I (I15324));
INVX1 gate4756(.O (I16100), .I (g9338));
INVX1 gate4757(.O (g6779), .I (I12208));
INVX1 gate4758(.O (I14857), .I (g8657));
INVX1 gate4759(.O (g3769), .I (g2548));
INVX1 gate4760(.O (I6952), .I (g1896));
INVX1 gate4761(.O (g8638), .I (I14722));
INVX1 gate4762(.O (g3836), .I (I7311));
INVX1 gate4763(.O (g5829), .I (I10512));
INVX1 gate4764(.O (g7587), .I (I13906));
INVX1 gate4765(.O (I13649), .I (g7281));
INVX1 gate4766(.O (g5286), .I (g4714));
INVX1 gate4767(.O (g1975), .I (g1253));
INVX1 gate4768(.O (I5747), .I (g1260));
INVX1 gate4769(.O (g4807), .I (I9142));
INVX1 gate4770(.O (g6977), .I (g6664));
INVX1 gate4771(.O (g7111), .I (I12921));
INVX1 gate4772(.O (I5855), .I (g71));
INVX1 gate4773(.O (I5398), .I (g702));
INVX1 gate4774(.O (g3918), .I (I7551));
INVX1 gate4775(.O (g2774), .I (g1813));
INVX1 gate4776(.O (g7275), .I (I13261));
INVX1 gate4777(.O (g7311), .I (I13365));
INVX1 gate4778(.O (g3967), .I (I7680));
INVX1 gate4779(.O (I6561), .I (g1715));
INVX1 gate4780(.O (I11648), .I (g6028));
INVX1 gate4781(.O (I10690), .I (g5538));
INVX1 gate4782(.O (g6588), .I (g5836));
INVX1 gate4783(.O (I11491), .I (g6010));
INVX1 gate4784(.O (I11903), .I (g5939));
INVX1 gate4785(.O (g9079), .I (I15631));
INVX1 gate4786(.O (I13903), .I (g7357));
INVX1 gate4787(.O (g8883), .I (I15225));
INVX1 gate4788(.O (g6161), .I (I10842));
INVX1 gate4789(.O (I7492), .I (g3561));
INVX1 gate4790(.O (g6361), .I (I11410));
INVX1 gate4791(.O (g4266), .I (I8202));
INVX1 gate4792(.O (g2396), .I (g1033));
INVX1 gate4793(.O (I7864), .I (g3812));
INVX1 gate4794(.O (I10548), .I (g5260));
INVX1 gate4795(.O (I13755), .I (g7317));
INVX1 gate4796(.O (g5733), .I (I10256));
INVX1 gate4797(.O (g7174), .I (g7097));
INVX1 gate4798(.O (g6051), .I (g5246));
INVX1 gate4799(.O (g3993), .I (g3192));
INVX1 gate4800(.O (g8217), .I (I14430));
INVX1 gate4801(.O (I13770), .I (g7491));
INVX1 gate4802(.O (I11981), .I (g6246));
INVX1 gate4803(.O (I9657), .I (g4784));
INVX1 gate4804(.O (I12968), .I (g6925));
INVX1 gate4805(.O (g1821), .I (g631));
INVX1 gate4806(.O (I15329), .I (g8793));
INVX1 gate4807(.O (g6327), .I (I11308));
INVX1 gate4808(.O (g2780), .I (I6517));
INVX1 gate4809(.O (I6764), .I (g1955));
INVX1 gate4810(.O (g3822), .I (g1815));
INVX1 gate4811(.O (g5610), .I (g4938));
INVX1 gate4812(.O (g2509), .I (g37));
INVX1 gate4813(.O (I15539), .I (g9005));
INVX1 gate4814(.O (g5073), .I (g4477));
INVX1 gate4815(.O (g5796), .I (I10427));
INVX1 gate4816(.O (I8565), .I (g3071));
INVX1 gate4817(.O (g5473), .I (g4903));
INVX1 gate4818(.O (g7284), .I (I13284));
INVX1 gate4819(.O (g6146), .I (I10801));
INVX1 gate4820(.O (g4081), .I (I7870));
INVX1 gate4821(.O (g7239), .I (g6945));
INVX1 gate4822(.O (g6346), .I (I11365));
INVX1 gate4823(.O (g7545), .I (I13819));
INVX1 gate4824(.O (I6970), .I (g1872));
INVX1 gate4825(.O (g2662), .I (I6457));
INVX1 gate4826(.O (g5124), .I (I9520));
INVX1 gate4827(.O (g7180), .I (I13092));
INVX1 gate4828(.O (g6103), .I (g5317));
INVX1 gate4829(.O (g4692), .I (I8971));
INVX1 gate4830(.O (g7591), .I (I13918));
INVX1 gate4831(.O (g6303), .I (I11236));
INVX1 gate4832(.O (g2467), .I (I6305));
INVX1 gate4833(.O (I9064), .I (g4302));
INVX1 gate4834(.O (I13767), .I (g7486));
INVX1 gate4835(.O (I13794), .I (g7346));
INVX1 gate4836(.O (I11395), .I (g5812));
INVX1 gate4837(.O (g5469), .I (g4898));
INVX1 gate4838(.O (g2290), .I (I6054));
INVX1 gate4839(.O (I7262), .I (g2514));
INVX1 gate4840(.O (I10128), .I (g4688));
INVX1 gate4841(.O (g6696), .I (I12022));
INVX1 gate4842(.O (g3921), .I (I7558));
INVX1 gate4843(.O (I9785), .I (g4747));
INVX1 gate4844(.O (I5577), .I (g172));
INVX1 gate4845(.O (g4960), .I (g4259));
INVX1 gate4846(.O (g7420), .I (I13537));
INVX1 gate4847(.O (I11633), .I (g5897));
INVX1 gate4848(.O (g5177), .I (I9657));
INVX1 gate4849(.O (I12894), .I (g7009));
INVX1 gate4850(.O (g7507), .I (I13701));
INVX1 gate4851(.O (g8774), .I (I14964));
INVX1 gate4852(.O (g5206), .I (g4938));
INVX1 gate4853(.O (I7623), .I (g3631));
INVX1 gate4854(.O (g2256), .I (g1324));
INVX1 gate4855(.O (I11191), .I (g6155));
INVX1 gate4856(.O (g2816), .I (g1685));
INVX1 gate4857(.O (I13719), .I (g7334));
INVX1 gate4858(.O (g6508), .I (I11686));
INVX1 gate4859(.O (g6944), .I (I12643));
INVX1 gate4860(.O (g3837), .I (I7314));
INVX1 gate4861(.O (g6072), .I (g5345));
INVX1 gate4862(.O (I11718), .I (g6115));
INVX1 gate4863(.O (g3062), .I (g2100));
INVX1 gate4864(.O (I14298), .I (g7678));
INVX1 gate4865(.O (g9032), .I (I15510));
INVX1 gate4866(.O (I5386), .I (g648));
INVX1 gate4867(.O (g3462), .I (g1743));
INVX1 gate4868(.O (g1756), .I (g533));
INVX1 gate4869(.O (g2381), .I (I6245));
INVX1 gate4870(.O (I5975), .I (g381));
INVX1 gate4871(.O (I11832), .I (g6274));
INVX1 gate4872(.O (g8780), .I (g8524));
INVX1 gate4873(.O (g9053), .I (I15557));
INVX1 gate4874(.O (I12202), .I (g6481));
INVX1 gate4875(.O (g4112), .I (I7947));
INVX1 gate4876(.O (g7905), .I (I14279));
INVX1 gate4877(.O (g4267), .I (I8205));
INVX1 gate4878(.O (g2700), .I (g1744));
INVX1 gate4879(.O (I7651), .I (g2573));
INVX1 gate4880(.O (I16107), .I (g9337));
INVX1 gate4881(.O (I8820), .I (g3952));
INVX1 gate4882(.O (I11440), .I (g6009));
INVX1 gate4883(.O (g2397), .I (g1272));
INVX1 gate4884(.O (I12496), .I (g6592));
INVX1 gate4885(.O (g5199), .I (g4841));
INVX1 gate4886(.O (g1904), .I (g1021));
INVX1 gate4887(.O (I12111), .I (g5956));
INVX1 gate4888(.O (g6316), .I (I11275));
INVX1 gate4889(.O (g7515), .I (I13725));
INVX1 gate4890(.O (I11861), .I (g5747));
INVX1 gate4891(.O (g8662), .I (I14780));
INVX1 gate4892(.O (g5781), .I (I10390));
INVX1 gate4893(.O (g4001), .I (g3160));
INVX1 gate4894(.O (g6034), .I (I10639));
INVX1 gate4895(.O (g8018), .I (I14315));
INVX1 gate4896(.O (I13861), .I (g7330));
INVX1 gate4897(.O (I9089), .I (g4566));
INVX1 gate4898(.O (g8067), .I (I14342));
INVX1 gate4899(.O (g2263), .I (g1394));
INVX1 gate4900(.O (g7100), .I (I12888));
INVX1 gate4901(.O (I13247), .I (g6906));
INVX1 gate4902(.O (I6299), .I (g47));
INVX1 gate4903(.O (g7300), .I (I13332));
INVX1 gate4904(.O (I11389), .I (g5766));
INVX1 gate4905(.O (I11926), .I (g6190));
INVX1 gate4906(.O (I12986), .I (g6931));
INVX1 gate4907(.O (g5797), .I (I10430));
INVX1 gate4908(.O (I15414), .I (g8900));
INVX1 gate4909(.O (I13045), .I (g6955));
INVX1 gate4910(.O (g6147), .I (I10804));
INVX1 gate4911(.O (I5984), .I (g540));
INVX1 gate4912(.O (g9157), .I (g9141));
INVX1 gate4913(.O (g6347), .I (I11368));
INVX1 gate4914(.O (I5939), .I (g275));
INVX1 gate4915(.O (I13099), .I (g7054));
INVX1 gate4916(.O (g3842), .I (I7329));
INVX1 gate4917(.O (I13388), .I (g7149));
INVX1 gate4918(.O (g8093), .I (I14370));
INVX1 gate4919(.O (g6681), .I (I11991));
INVX1 gate4920(.O (I11701), .I (g5772));
INVX1 gate4921(.O (g8493), .I (g8041));
INVX1 gate4922(.O (I13701), .I (g7349));
INVX1 gate4923(.O (I10512), .I (g5238));
INVX1 gate4924(.O (g3085), .I (g1945));
INVX1 gate4925(.O (I8775), .I (g4019));
INVX1 gate4926(.O (I7838), .I (g2781));
INVX1 gate4927(.O (I8922), .I (g4229));
INVX1 gate4928(.O (I11251), .I (g6152));
INVX1 gate4929(.O (I11272), .I (g5758));
INVX1 gate4930(.O (g7750), .I (I14121));
INVX1 gate4931(.O (g3485), .I (g1737));
INVX1 gate4932(.O (g2562), .I (g1652));
INVX1 gate4933(.O (g1695), .I (g778));
INVX1 gate4934(.O (g6697), .I (I12025));
INVX1 gate4935(.O (g1637), .I (g1087));
INVX1 gate4936(.O (g5144), .I (I9558));
INVX1 gate4937(.O (g4592), .I (g2938));
INVX1 gate4938(.O (g5344), .I (I9819));
INVX1 gate4939(.O (g6210), .I (I10969));
INVX1 gate4940(.O (I5636), .I (g891));
INVX1 gate4941(.O (g2631), .I (g1586));
INVX1 gate4942(.O (g4746), .I (I9076));
INVX1 gate4943(.O (I12877), .I (g6700));
INVX1 gate4944(.O (g8181), .I (I14420));
INVX1 gate4945(.O (g6596), .I (I11800));
INVX1 gate4946(.O (g5207), .I (g4673));
INVX1 gate4947(.O (g8381), .I (I14603));
INVX1 gate4948(.O (g3854), .I (I7365));
INVX1 gate4949(.O (g2817), .I (g1849));
INVX1 gate4950(.O (g3941), .I (I7626));
INVX1 gate4951(.O (I7672), .I (g3062));
INVX1 gate4952(.O (I16135), .I (g9357));
INVX1 gate4953(.O (g4703), .I (I8998));
INVX1 gate4954(.O (g5819), .I (I10482));
INVX1 gate4955(.O (g8685), .I (I14851));
INVX1 gate4956(.O (g7440), .I (I13577));
INVX1 gate4957(.O (I10445), .I (g5418));
INVX1 gate4958(.O (I7523), .I (g2562));
INVX1 gate4959(.O (I14445), .I (g8067));
INVX1 gate4960(.O (I12196), .I (g6471));
INVX1 gate4961(.O (I6078), .I (g95));
INVX1 gate4962(.O (g2605), .I (g1639));
INVX1 gate4963(.O (I13140), .I (g6954));
INVX1 gate4964(.O (I9350), .I (g4503));
INVX1 gate4965(.O (g7123), .I (I12961));
INVX1 gate4966(.O (g8421), .I (g8017));
INVX1 gate4967(.O (g5088), .I (I9466));
INVX1 gate4968(.O (I8784), .I (g3949));
INVX1 gate4969(.O (I13997), .I (g7432));
INVX1 gate4970(.O (I8739), .I (g3910));
INVX1 gate4971(.O (g1757), .I (g604));
INVX1 gate4972(.O (g5488), .I (I9910));
INVX1 gate4973(.O (g4932), .I (g4202));
INVX1 gate4974(.O (I12526), .I (g6626));
INVX1 gate4975(.O (I15759), .I (g9082));
INVX1 gate4976(.O (g5701), .I (g5120));
INVX1 gate4977(.O (g6820), .I (I12331));
INVX1 gate4978(.O (g4624), .I (I8787));
INVX1 gate4979(.O (I9009), .I (g4591));
INVX1 gate4980(.O (I6959), .I (g1558));
INVX1 gate4981(.O (g3520), .I (g1616));
INVX1 gate4982(.O (g6936), .I (I12629));
INVX1 gate4983(.O (g3219), .I (I6872));
INVX1 gate4984(.O (I6517), .I (g1687));
INVX1 gate4985(.O (g3640), .I (I7112));
INVX1 gate4986(.O (I16049), .I (g9288));
INVX1 gate4987(.O (g6117), .I (I10739));
INVX1 gate4988(.O (g1811), .I (I5679));
INVX1 gate4989(.O (g6317), .I (I11278));
INVX1 gate4990(.O (I7551), .I (g2712));
INVX1 gate4991(.O (I7104), .I (g2479));
INVX1 gate4992(.O (g3812), .I (g1750));
INVX1 gate4993(.O (I12457), .I (g6671));
INVX1 gate4994(.O (g7528), .I (I13764));
INVX1 gate4995(.O (I14722), .I (g8076));
INVX1 gate4996(.O (g7151), .I (I13035));
INVX1 gate4997(.O (g3958), .I (g3097));
INVX1 gate4998(.O (g7351), .I (I13469));
INVX1 gate4999(.O (g4677), .I (I8932));
INVX1 gate5000(.O (g6601), .I (g6083));
INVX1 gate5001(.O (g7530), .I (I13770));
INVX1 gate5002(.O (I12866), .I (g6483));
INVX1 gate5003(.O (I8190), .I (g3545));
INVX1 gate5004(.O (g8562), .I (g8094));
INVX1 gate5005(.O (I9918), .I (g4968));
INVX1 gate5006(.O (I10271), .I (g5487));
INVX1 gate5007(.O (g5114), .I (I9502));
INVX1 gate5008(.O (g4576), .I (g2913));
INVX1 gate5009(.O (I15940), .I (g9213));
INVX1 gate5010(.O (I13447), .I (g7261));
INVX1 gate5011(.O (g8631), .I (I14709));
INVX1 gate5012(.O (g2673), .I (I6474));
INVX1 gate5013(.O (g6775), .I (I12196));
INVX1 gate5014(.O (g3829), .I (I7290));
INVX1 gate5015(.O (g6922), .I (g6525));
INVX1 gate5016(.O (I5763), .I (g1207));
INVX1 gate5017(.O (g3911), .I (I7526));
INVX1 gate5018(.O (I6214), .I (g7));
INVX1 gate5019(.O (g6581), .I (I11773));
INVX1 gate5020(.O (g5825), .I (I10500));
INVX1 gate5021(.O (I14342), .I (g7582));
INVX1 gate5022(.O (g8605), .I (I14680));
INVX1 gate5023(.O (I14145), .I (g7542));
INVX1 gate5024(.O (I12256), .I (g6647));
INVX1 gate5025(.O (I14031), .I (g7448));
INVX1 gate5026(.O (g4198), .I (I8101));
INVX1 gate5027(.O (I7044), .I (g2402));
INVX1 gate5028(.O (g6597), .I (I11803));
INVX1 gate5029(.O (g9075), .I (I15619));
INVX1 gate5030(.O (I13451), .I (g7262));
INVX1 gate5031(.O (I13472), .I (g7266));
INVX1 gate5032(.O (I14199), .I (g7704));
INVX1 gate5033(.O (I12280), .I (g6684));
INVX1 gate5034(.O (g3974), .I (g3131));
INVX1 gate5035(.O (I6663), .I (g2246));
INVX1 gate5036(.O (I13628), .I (g7248));
INVX1 gate5037(.O (g8751), .I (g8545));
INVX1 gate5038(.O (g2458), .I (g30));
INVX1 gate5039(.O (I5359), .I (g3839));
INVX1 gate5040(.O (g6784), .I (I12223));
INVX1 gate5041(.O (g2743), .I (g1808));
INVX1 gate5042(.O (g3610), .I (g2424));
INVX1 gate5043(.O (g2890), .I (g2264));
INVX1 gate5044(.O (g5768), .I (I10377));
INVX1 gate5045(.O (I10528), .I (g5245));
INVX1 gate5046(.O (I16033), .I (g9282));
INVX1 gate5047(.O (g8585), .I (g7993));
INVX1 gate5048(.O (g1612), .I (I5475));
INVX1 gate5049(.O (I10393), .I (g5196));
INVX1 gate5050(.O (g7172), .I (g7092));
INVX1 gate5051(.O (g1017), .I (I5419));
INVX1 gate5052(.O (I7712), .I (g3657));
INVX1 gate5053(.O (I14330), .I (g7538));
INVX1 gate5054(.O (g2505), .I (g28));
INVX1 gate5055(.O (g8041), .I (g7701));
INVX1 gate5056(.O (I15962), .I (g9218));
INVX1 gate5057(.O (g2011), .I (I5847));
INVX1 gate5058(.O (g3124), .I (g1857));
INVX1 gate5059(.O (g5806), .I (I10451));
INVX1 gate5060(.O (I5416), .I (g8868));
INVX1 gate5061(.O (g1935), .I (g1280));
INVX1 gate5062(.O (g3980), .I (g3192));
INVX1 gate5063(.O (g6937), .I (I12632));
INVX1 gate5064(.O (g7143), .I (g6996));
INVX1 gate5065(.O (I11591), .I (g5814));
INVX1 gate5066(.O (g2734), .I (g2170));
INVX1 gate5067(.O (g7343), .I (I13447));
INVX1 gate5068(.O (I13776), .I (g7497));
INVX1 gate5069(.O (g9039), .I (I15527));
INVX1 gate5070(.O (g4524), .I (g2869));
INVX1 gate5071(.O (g6294), .I (I11209));
INVX1 gate5072(.O (g6840), .I (I12391));
INVX1 gate5073(.O (g4644), .I (I8847));
INVX1 gate5074(.O (I6590), .I (g2467));
INVX1 gate5075(.O (I13147), .I (g7024));
INVX1 gate5076(.O (g8673), .I (I14813));
INVX1 gate5077(.O (g3540), .I (g2424));
INVX1 gate5078(.O (I15833), .I (g9162));
INVX1 gate5079(.O (g4119), .I (I7964));
INVX1 gate5080(.O (I9837), .I (g4781));
INVX1 gate5081(.O (g6190), .I (I10933));
INVX1 gate5082(.O (g2074), .I (I5872));
INVX1 gate5083(.O (I6657), .I (g1701));
INVX1 gate5084(.O (g6390), .I (I11497));
INVX1 gate5085(.O (g7134), .I (I12986));
INVX1 gate5086(.O (I12885), .I (g6946));
INVX1 gate5087(.O (g7334), .I (I13422));
INVX1 gate5088(.O (I13825), .I (g7318));
INVX1 gate5089(.O (g2992), .I (g1833));
INVX1 gate5090(.O (g4258), .I (I8193));
INVX1 gate5091(.O (I11858), .I (g6165));
INVX1 gate5092(.O (g4577), .I (g2914));
INVX1 gate5093(.O (g6501), .I (I11669));
INVX1 gate5094(.O (g7548), .I (I13828));
INVX1 gate5095(.O (g8669), .I (I14801));
INVX1 gate5096(.O (g4867), .I (I9209));
INVX1 gate5097(.O (I13858), .I (g7329));
INVX1 gate5098(.O (I14709), .I (g8198));
INVX1 gate5099(.O (I10259), .I (g5362));
INVX1 gate5100(.O (g6156), .I (I10829));
INVX1 gate5101(.O (I12511), .I (g6598));
INVX1 gate5102(.O (g6356), .I (I11395));
INVX1 gate5103(.O (g5433), .I (g5024));
INVX1 gate5104(.O (I10708), .I (g5545));
INVX1 gate5105(.O (g7555), .I (I13843));
INVX1 gate5106(.O (g1800), .I (g1477));
INVX1 gate5107(.O (I12763), .I (g6686));
INVX1 gate5108(.O (g3287), .I (I6911));
INVX1 gate5109(.O (g8772), .I (g8585));
INVX1 gate5110(.O (I7885), .I (g2837));
INVX1 gate5111(.O (I5654), .I (g921));
INVX1 gate5112(.O (I8357), .I (g1182));
INVX1 gate5113(.O (I6930), .I (g1876));
INVX1 gate5114(.O (g2573), .I (g1649));
INVX1 gate5115(.O (g2863), .I (g1778));
INVX1 gate5116(.O (g7792), .I (I14231));
INVX1 gate5117(.O (g2480), .I (g44));
INVX1 gate5118(.O (I15613), .I (g8996));
INVX1 gate5119(.O (I9788), .I (g4711));
INVX1 gate5120(.O (g8743), .I (g8524));
INVX1 gate5121(.O (g3849), .I (I7350));
INVX1 gate5122(.O (g6704), .I (I12044));
INVX1 gate5123(.O (I15947), .I (g9221));
INVX1 gate5124(.O (g5845), .I (I10548));
INVX1 gate5125(.O (g4599), .I (I8712));
INVX1 gate5126(.O (g5137), .I (I9539));
INVX1 gate5127(.O (g5395), .I (I9840));
INVX1 gate5128(.O (g8856), .I (I15160));
INVX1 gate5129(.O (g7113), .I (I12927));
INVX1 gate5130(.O (g3898), .I (g3160));
INVX1 gate5131(.O (g8734), .I (I14904));
INVX1 gate5132(.O (g4026), .I (g3192));
INVX1 gate5133(.O (g7313), .I (I13369));
INVX1 gate5134(.O (g4274), .I (I8218));
INVX1 gate5135(.O (g4426), .I (I8428));
INVX1 gate5136(.O (I7036), .I (g2454));
INVX1 gate5137(.O (g6250), .I (g5679));
INVX1 gate5138(.O (g6810), .I (I12301));
INVX1 gate5139(.O (g4614), .I (I8757));
INVX1 gate5140(.O (g6363), .I (I11416));
INVX1 gate5141(.O (g4370), .I (I8351));
INVX1 gate5142(.O (I5978), .I (g414));
INVX1 gate5143(.O (g3510), .I (g2185));
INVX1 gate5144(.O (I10810), .I (g5403));
INVX1 gate5145(.O (g6032), .I (g5494));
INVX1 gate5146(.O (I11446), .I (g6062));
INVX1 gate5147(.O (g4125), .I (I7978));
INVX1 gate5148(.O (I14810), .I (g8481));
INVX1 gate5149(.O (I11227), .I (g6130));
INVX1 gate5150(.O (g6432), .I (I11569));
INVX1 gate5151(.O (g5807), .I (I10454));
INVX1 gate5152(.O (I14657), .I (g7782));
INVX1 gate5153(.O (g7094), .I (g6525));
INVX1 gate5154(.O (I12307), .I (g6712));
INVX1 gate5155(.O (I11025), .I (g5638));
INVX1 gate5156(.O (I12085), .I (g5971));
INVX1 gate5157(.O (g2976), .I (I6728));
INVX1 gate5158(.O (I7335), .I (g2910));
INVX1 gate5159(.O (g1823), .I (g768));
INVX1 gate5160(.O (g7494), .I (g7260));
INVX1 gate5161(.O (g7518), .I (I13734));
INVX1 gate5162(.O (g5266), .I (I9782));
INVX1 gate5163(.O (g6568), .I (I11744));
INVX1 gate5164(.O (g4544), .I (g2886));
INVX1 gate5165(.O (I11203), .I (g6129));
INVX1 gate5166(.O (I5542), .I (g1272));
INVX1 gate5167(.O (I13203), .I (g7088));
INVX1 gate5168(.O (g7776), .I (I14199));
INVX1 gate5169(.O (g1649), .I (g1217));
INVX1 gate5170(.O (I7749), .I (g3692));
INVX1 gate5171(.O (g7593), .I (I13924));
INVX1 gate5172(.O (g3819), .I (g1748));
INVX1 gate5173(.O (g4636), .I (I8823));
INVX1 gate5174(.O (g3694), .I (g2174));
INVX1 gate5175(.O (g2326), .I (I6121));
INVX1 gate5176(.O (I14792), .I (g8583));
INVX1 gate5177(.O (I9520), .I (g3995));
INVX1 gate5178(.O (g6357), .I (I11398));
INVX1 gate5179(.O (g4106), .I (I7931));
INVX1 gate5180(.O (I15507), .I (g8968));
INVX1 gate5181(.O (I12942), .I (g7023));
INVX1 gate5182(.O (g3852), .I (I7359));
INVX1 gate5183(.O (I6471), .I (g1923));
INVX1 gate5184(.O (g3923), .I (I7564));
INVX1 gate5185(.O (g4306), .I (I8273));
INVX1 gate5186(.O (I8778), .I (g3922));
INVX1 gate5187(.O (I11281), .I (g5785));
INVX1 gate5188(.O (I12268), .I (g6661));
INVX1 gate5189(.O (g9320), .I (g9307));
INVX1 gate5190(.O (g5481), .I (g4914));
INVX1 gate5191(.O (g3488), .I (g1727));
INVX1 gate5192(.O (I7947), .I (g3485));
INVX1 gate5193(.O (I13281), .I (g7155));
INVX1 gate5194(.O (g1698), .I (I5542));
INVX1 gate5195(.O (I6242), .I (g1554));
INVX1 gate5196(.O (I16173), .I (g9382));
INVX1 gate5197(.O (I12655), .I (g6458));
INVX1 gate5198(.O (I11377), .I (g5811));
INVX1 gate5199(.O (g7264), .I (I13234));
INVX1 gate5200(.O (g5726), .I (I10243));
INVX1 gate5201(.O (g5154), .I (I9588));
INVX1 gate5202(.O (I10919), .I (g5479));
INVX1 gate5203(.O (I9005), .I (g4585));
INVX1 gate5204(.O (g7160), .I (I13054));
INVX1 gate5205(.O (g7360), .I (I13496));
INVX1 gate5206(.O (I11562), .I (g5939));
INVX1 gate5207(.O (I11645), .I (g5874));
INVX1 gate5208(.O (I13562), .I (g7179));
INVX1 gate5209(.O (g7521), .I (I13743));
INVX1 gate5210(.O (g4622), .I (I8781));
INVX1 gate5211(.O (g4027), .I (g2845));
INVX1 gate5212(.O (g2183), .I (I5908));
INVX1 gate5213(.O (g3951), .I (I7648));
INVX1 gate5214(.O (g7050), .I (g6618));
INVX1 gate5215(.O (I6254), .I (g536));
INVX1 gate5216(.O (g2383), .I (I6251));
INVX1 gate5217(.O (g2924), .I (g2314));
INVX1 gate5218(.O (I12839), .I (g6630));
INVX1 gate5219(.O (I12930), .I (g7019));
INVX1 gate5220(.O (I8949), .I (g4116));
INVX1 gate5221(.O (I7632), .I (g3634));
INVX1 gate5222(.O (I7095), .I (g2539));
INVX1 gate5223(.O (I12993), .I (g6933));
INVX1 gate5224(.O (I10545), .I (g5259));
INVX1 gate5225(.O (g6626), .I (I11870));
INVX1 gate5226(.O (I11290), .I (g5818));
INVX1 gate5227(.O (I13290), .I (g7158));
INVX1 gate5228(.O (I7495), .I (g3562));
INVX1 gate5229(.O (I14079), .I (g7579));
INVX1 gate5230(.O (g4904), .I (g4085));
INVX1 gate5231(.O (g4200), .I (I8105));
INVX1 gate5232(.O (I13698), .I (g7348));
INVX1 gate5233(.O (I7302), .I (g2825));
INVX1 gate5234(.O (I12965), .I (g6924));
INVX1 gate5235(.O (I12131), .I (g5918));
INVX1 gate5236(.O (g9299), .I (I16023));
INVX1 gate5237(.O (I6009), .I (g359));
INVX1 gate5238(.O (g3870), .I (g3466));
INVX1 gate5239(.O (I8998), .I (g4576));
INVX1 gate5240(.O (I5512), .I (g557));
INVX1 gate5241(.O (g4003), .I (g3192));
INVX1 gate5242(.O (I9974), .I (g4676));
INVX1 gate5243(.O (g5112), .I (I9496));
INVX1 gate5244(.O (g3825), .I (g1826));
INVX1 gate5245(.O (g3650), .I (I7126));
INVX1 gate5246(.O (g5267), .I (I9785));
INVX1 gate5247(.O (I12487), .I (g6623));
INVX1 gate5248(.O (g4841), .I (g4250));
INVX1 gate5249(.O (g2161), .I (g1454));
INVX1 gate5250(.O (I8084), .I (g3706));
INVX1 gate5251(.O (g1652), .I (g1220));
INVX1 gate5252(.O (g2361), .I (I6183));
INVX1 gate5253(.O (I7752), .I (g3591));
INVX1 gate5254(.O (I12502), .I (g6604));
INVX1 gate5255(.O (g4191), .I (I8084));
INVX1 gate5256(.O (g1843), .I (g771));
INVX1 gate5257(.O (g8760), .I (g8545));
INVX1 gate5258(.O (g3008), .I (g1816));
INVX1 gate5259(.O (I8850), .I (g4031));
INVX1 gate5260(.O (g2665), .I (g1661));
INVX1 gate5261(.O (g7289), .I (I13299));
INVX1 gate5262(.O (g7777), .I (I14202));
INVX1 gate5263(.O (g6683), .I (g6237));
INVX1 gate5264(.O (g5401), .I (I9845));
INVX1 gate5265(.O (I10125), .I (g5127));
INVX1 gate5266(.O (g4695), .I (I8980));
INVX1 gate5267(.O (I10532), .I (g5253));
INVX1 gate5268(.O (g4637), .I (I8826));
INVX1 gate5269(.O (I5649), .I (g1389));
INVX1 gate5270(.O (g7835), .I (I14257));
INVX1 gate5271(.O (g2327), .I (I6124));
INVX1 gate5272(.O (g5129), .I (I9531));
INVX1 gate5273(.O (g6778), .I (I12205));
INVX1 gate5274(.O (g5761), .I (I10356));
INVX1 gate5275(.O (g3768), .I (g2253));
INVX1 gate5276(.O (I10783), .I (g5542));
INVX1 gate5277(.O (g6894), .I (g6525));
INVX1 gate5278(.O (I13403), .I (g7269));
INVX1 gate5279(.O (I13547), .I (g1170));
INVX1 gate5280(.O (g4307), .I (g3700));
INVX1 gate5281(.O (g4536), .I (g2877));
INVX1 gate5282(.O (g2999), .I (g1823));
INVX1 gate5283(.O (I14783), .I (g8324));
INVX1 gate5284(.O (g3972), .I (I7691));
INVX1 gate5285(.O (g1686), .I (I5531));
INVX1 gate5286(.O (g5828), .I (I10509));
INVX1 gate5287(.O (g2346), .I (I6154));
INVX1 gate5288(.O (g2633), .I (g1577));
INVX1 gate5289(.O (I12469), .I (g6586));
INVX1 gate5290(.O (g9244), .I (I15974));
INVX1 gate5291(.O (I10561), .I (g5265));
INVX1 gate5292(.O (I6229), .I (g486));
INVX1 gate5293(.O (g8608), .I (I14687));
INVX1 gate5294(.O (g8220), .I (I14439));
INVX1 gate5295(.O (I10353), .I (g5710));
INVX1 gate5296(.O (I12286), .I (g6696));
INVX1 gate5297(.O (g6782), .I (I12217));
INVX1 gate5298(.O (I7164), .I (g2157));
INVX1 gate5299(.O (I10295), .I (g5523));
INVX1 gate5300(.O (I8919), .I (g4196));
INVX1 gate5301(.O (g3943), .I (I7632));
INVX1 gate5302(.O (g9140), .I (I15784));
INVX1 gate5303(.O (I9177), .I (g4299));
INVX1 gate5304(.O (g9078), .I (I15628));
INVX1 gate5305(.O (g9340), .I (I16090));
INVX1 gate5306(.O (I13481), .I (g7254));
INVX1 gate5307(.O (g5592), .I (g4969));
INVX1 gate5308(.O (I14680), .I (g7810));
INVX1 gate5309(.O (g6661), .I (I11961));
INVX1 gate5310(.O (g6075), .I (g5345));
INVX1 gate5311(.O (g4016), .I (g3192));
INVX1 gate5312(.O (I8952), .I (g4197));
INVX1 gate5313(.O (g699), .I (I5395));
INVX1 gate5314(.O (I12038), .I (g5847));
INVX1 gate5315(.O (g5746), .I (I10295));
INVX1 gate5316(.O (g6475), .I (I11633));
INVX1 gate5317(.O (g9035), .I (I15519));
INVX1 gate5318(.O (g1670), .I (g1489));
INVX1 gate5319(.O (g3465), .I (I6963));
INVX1 gate5320(.O (g8977), .I (I15433));
INVX1 gate5321(.O (I7296), .I (g2915));
INVX1 gate5322(.O (g3934), .I (I7599));
INVX1 gate5323(.O (g9082), .I (I15638));
INVX1 gate5324(.O (g3230), .I (I6887));
INVX1 gate5325(.O (g4522), .I (g2867));
INVX1 gate5326(.O (g4115), .I (I7956));
INVX1 gate5327(.O (g4251), .I (I8180));
INVX1 gate5328(.O (g6292), .I (I11203));
INVX1 gate5329(.O (I12187), .I (g5897));
INVX1 gate5330(.O (g4811), .I (I9158));
INVX1 gate5331(.O (g4642), .I (I8841));
INVX1 gate5332(.O (g7541), .I (I13807));
INVX1 gate5333(.O (g2944), .I (g2363));
INVX1 gate5334(.O (g2240), .I (I5981));
INVX1 gate5335(.O (g1938), .I (g1288));
INVX1 gate5336(.O (g1813), .I (g620));
INVX1 gate5337(.O (g6646), .I (I11920));
INVX1 gate5338(.O (g7132), .I (I12980));
INVX1 gate5339(.O (I8986), .I (g4552));
INVX1 gate5340(.O (g8665), .I (I14789));
INVX1 gate5341(.O (g7332), .I (I13416));
INVX1 gate5342(.O (I13490), .I (g7130));
INVX1 gate5343(.O (g1909), .I (g998));
INVX1 gate5344(.O (g7353), .I (I13475));
INVX1 gate5345(.O (g6603), .I (I11815));
INVX1 gate5346(.O (g3096), .I (I6834));
INVX1 gate5347(.O (I5872), .I (g77));
INVX1 gate5348(.O (I13956), .I (g7499));
INVX1 gate5349(.O (g5468), .I (I9884));
INVX1 gate5350(.O (g6850), .I (I12421));
INVX1 gate5351(.O (g3496), .I (I6974));
INVX1 gate5352(.O (g7744), .I (I14103));
INVX1 gate5353(.O (g4654), .I (I8877));
INVX1 gate5354(.O (I13103), .I (g7055));
INVX1 gate5355(.O (g3845), .I (I7338));
INVX1 gate5356(.O (g2316), .I (I6109));
INVX1 gate5357(.O (g9214), .I (I15918));
INVX1 gate5358(.O (I5989), .I (g1460));
INVX1 gate5359(.O (I7389), .I (g3496));
INVX1 gate5360(.O (I11824), .I (g6283));
INVX1 gate5361(.O (g5677), .I (I10166));
INVX1 gate5362(.O (I7706), .I (g2584));
INVX1 gate5363(.O (I13888), .I (g7335));
INVX1 gate5364(.O (g3891), .I (g3097));
INVX1 gate5365(.O (I8925), .I (g4482));
INVX1 gate5366(.O (g3913), .I (g2834));
INVX1 gate5367(.O (I10289), .I (g5569));
INVX1 gate5368(.O (g9110), .I (I15720));
INVX1 gate5369(.O (g9310), .I (I16046));
INVX1 gate5370(.O (g6702), .I (I12038));
INVX1 gate5371(.O (g7558), .I (I13850));
INVX1 gate5372(.O (I7888), .I (g3505));
INVX1 gate5373(.O (g4595), .I (g2942));
INVX1 gate5374(.O (g4537), .I (g2878));
INVX1 gate5375(.O (I15927), .I (g9208));
INVX1 gate5376(.O (I7029), .I (g2392));
INVX1 gate5377(.O (g1687), .I (g10));
INVX1 gate5378(.O (I7371), .I (g3050));
INVX1 gate5379(.O (g2347), .I (I6157));
INVX1 gate5380(.O (I12666), .I (g6476));
INVX1 gate5381(.O (g5149), .I (I9573));
INVX1 gate5382(.O (I14288), .I (g7705));
INVX1 gate5383(.O (I14224), .I (g7722));
INVX1 gate5384(.O (I9344), .I (g4341));
INVX1 gate5385(.O (I12217), .I (g6631));
INVX1 gate5386(.O (I7956), .I (g2810));
INVX1 gate5387(.O (g1586), .I (g730));
INVX1 gate5388(.O (I6788), .I (g1681));
INVX1 gate5389(.O (I12478), .I (g6603));
INVX1 gate5390(.O (g2533), .I (g1336));
INVX1 gate5391(.O (g8753), .I (I14925));
INVX1 gate5392(.O (g3859), .I (I7380));
INVX1 gate5393(.O (g4612), .I (I8751));
INVX1 gate5394(.O (g7511), .I (I13713));
INVX1 gate5395(.O (g4017), .I (g2845));
INVX1 gate5396(.O (I15648), .I (g9044));
INVX1 gate5397(.O (g2914), .I (g2308));
INVX1 gate5398(.O (I8277), .I (g3504));
INVX1 gate5399(.O (g5198), .I (g4969));
INVX1 gate5400(.O (I9819), .I (g4691));
INVX1 gate5401(.O (g8072), .I (I14349));
INVX1 gate5402(.O (g9236), .I (I15962));
INVX1 gate5403(.O (g2210), .I (g1326));
INVX1 gate5404(.O (g6616), .I (I11848));
INVX1 gate5405(.O (g4935), .I (g4202));
INVX1 gate5406(.O (g7092), .I (I12866));
INVX1 gate5407(.O (I5670), .I (g941));
INVX1 gate5408(.O (I15604), .I (g8993));
INVX1 gate5409(.O (g7492), .I (I13656));
INVX1 gate5410(.O (I14816), .I (g8642));
INVX1 gate5411(.O (g1570), .I (g665));
INVX1 gate5412(.O (g1860), .I (g162));
INVX1 gate5413(.O (g8443), .I (g8015));
INVX1 gate5414(.O (I6192), .I (g327));
INVX1 gate5415(.O (g7574), .I (I13869));
INVX1 gate5416(.O (g6004), .I (g5494));
INVX1 gate5417(.O (I15770), .I (g9121));
INVX1 gate5418(.O (I10687), .I (g5674));
INVX1 gate5419(.O (g4629), .I (I8802));
INVX1 gate5420(.O (I10976), .I (g5726));
INVX1 gate5421(.O (g6404), .I (I11525));
INVX1 gate5422(.O (I12223), .I (g6655));
INVX1 gate5423(.O (g4328), .I (g3086));
INVX1 gate5424(.O (I14687), .I (g7826));
INVX1 gate5425(.O (g7714), .I (I14019));
INVX1 gate5426(.O (g6647), .I (I11923));
INVX1 gate5427(.O (g4130), .I (I7987));
INVX1 gate5428(.O (g4542), .I (g2884));
INVX1 gate5429(.O (I10752), .I (g5618));
INVX1 gate5430(.O (g3815), .I (g1822));
INVX1 gate5431(.O (I7338), .I (g2923));
INVX1 gate5432(.O (g6764), .I (I12161));
INVX1 gate5433(.O (I14374), .I (g7693));
INVX1 gate5434(.O (I10643), .I (g5267));
INVX1 gate5435(.O (g3692), .I (I7198));
INVX1 gate5436(.O (I13088), .I (g7045));
INVX1 gate5437(.O (g9222), .I (I15940));
INVX1 gate5438(.O (I14643), .I (g7837));
INVX1 gate5439(.O (g2936), .I (I6680));
INVX1 gate5440(.O (g3497), .I (g2185));
INVX1 gate5441(.O (g5524), .I (I9938));
INVX1 gate5442(.O (g7580), .I (I13885));
INVX1 gate5443(.O (g4800), .I (I9123));
INVX1 gate5444(.O (g5644), .I (g4748));
INVX1 gate5445(.O (I15845), .I (g9174));
INVX1 gate5446(.O (g3960), .I (I7667));
INVX1 gate5447(.O (I8892), .I (g4115));
INVX1 gate5448(.O (g1879), .I (I5763));
INVX1 gate5449(.O (g4554), .I (g2892));
INVX1 gate5450(.O (I11497), .I (g6014));
INVX1 gate5451(.O (g9064), .I (I15586));
INVX1 gate5452(.O (I15990), .I (g9239));
INVX1 gate5453(.O (I5552), .I (g1284));
INVX1 gate5454(.O (g7262), .I (I13228));
INVX1 gate5455(.O (g5152), .I (I9582));
INVX1 gate5456(.O (g5258), .I (I9774));
INVX1 gate5457(.O (I14260), .I (g7717));
INVX1 gate5458(.O (g7736), .I (I14079));
INVX1 gate5459(.O (g5818), .I (I10479));
INVX1 gate5460(.O (I10842), .I (g5701));
INVX1 gate5461(.O (g6224), .I (I11011));
INVX1 gate5462(.O (g5577), .I (I10046));
INVX1 gate5463(.O (I14668), .I (g7787));
INVX1 gate5464(.O (I11659), .I (g5897));
INVX1 gate5465(.O (g5717), .I (g4969));
INVX1 gate5466(.O (I13126), .I (g6949));
INVX1 gate5467(.O (I13659), .I (g7232));
INVX1 gate5468(.O (I8945), .I (g4106));
INVX1 gate5469(.O (I11987), .I (g6278));
INVX1 gate5470(.O (g6320), .I (I11287));
INVX1 gate5471(.O (I12373), .I (g6763));
INVX1 gate5472(.O (I6431), .I (g1825));
INVX1 gate5473(.O (I13250), .I (g7036));
INVX1 gate5474(.O (I14489), .I (g7829));
INVX1 gate5475(.O (g2922), .I (g2313));
INVX1 gate5476(.O (g1587), .I (g734));
INVX1 gate5477(.O (g3783), .I (I7255));
INVX1 gate5478(.O (g8013), .I (g7561));
INVX1 gate5479(.O (I10525), .I (g5244));
INVX1 gate5480(.O (I10488), .I (g5230));
INVX1 gate5481(.O (I16061), .I (g9294));
INVX1 gate5482(.O (I10424), .I (g5209));
INVX1 gate5483(.O (g7476), .I (g7229));
INVX1 gate5484(.O (I8709), .I (g4191));
INVX1 gate5485(.O (g3979), .I (I7702));
INVX1 gate5486(.O (I14424), .I (g7652));
INVX1 gate5487(.O (I6376), .I (g38));
INVX1 gate5488(.O (g5186), .I (I9684));
INVX1 gate5489(.O (I10558), .I (g5264));
INVX1 gate5490(.O (I8140), .I (g3429));
INVX1 gate5491(.O (I12936), .I (g7015));
INVX1 gate5492(.O (g9237), .I (I15965));
INVX1 gate5493(.O (I9136), .I (g4280));
INVX1 gate5494(.O (I11296), .I (g5831));
INVX1 gate5495(.O (I9336), .I (g4493));
INVX1 gate5496(.O (g6617), .I (I11851));
INVX1 gate5497(.O (g6789), .I (I12238));
INVX1 gate5498(.O (I13296), .I (g7161));
INVX1 gate5499(.O (g4512), .I (g2842));
INVX1 gate5500(.O (g2460), .I (I6302));
INVX1 gate5501(.O (I7098), .I (g2477));
INVX1 gate5502(.O (I8907), .I (g4095));
INVX1 gate5503(.O (I11338), .I (g5798));
INVX1 gate5504(.O (g7722), .I (I14039));
INVX1 gate5505(.O (I12334), .I (g6713));
INVX1 gate5506(.O (I13338), .I (g7190));
INVX1 gate5507(.O (I9594), .I (g4718));
INVX1 gate5508(.O (I7498), .I (g2752));
INVX1 gate5509(.O (g5026), .I (I9366));
INVX1 gate5510(.O (I6286), .I (g1307));
INVX1 gate5511(.O (g3676), .I (g2380));
INVX1 gate5512(.O (g9194), .I (g9182));
INVX1 gate5513(.O (g5426), .I (g5013));
INVX1 gate5514(.O (I6911), .I (g1869));
INVX1 gate5515(.O (I8517), .I (g3014));
INVX1 gate5516(.O (g7285), .I (I13287));
INVX1 gate5517(.O (g2784), .I (g2340));
INVX1 gate5518(.O (g5170), .I (I9636));
INVX1 gate5519(.O (g3761), .I (g1772));
INVX1 gate5520(.O (g4056), .I (g3082));
INVX1 gate5521(.O (g7500), .I (I13676));
INVX1 gate5522(.O (I11060), .I (g5453));
INVX1 gate5523(.O (g9089), .I (I15657));
INVX1 gate5524(.O (I13060), .I (g6959));
INVX1 gate5525(.O (g6299), .I (I11224));
INVX1 gate5526(.O (g5821), .I (I10488));
INVX1 gate5527(.O (I11197), .I (g6122));
INVX1 gate5528(.O (g3828), .I (I7287));
INVX1 gate5529(.O (g4649), .I (I8862));
INVX1 gate5530(.O (I7584), .I (g3062));
INVX1 gate5531(.O (I11855), .I (g5751));
INVX1 gate5532(.O (I6733), .I (g1718));
INVX1 gate5533(.O (g3830), .I (I7293));
INVX1 gate5534(.O (I6974), .I (g2528));
INVX1 gate5535(.O (I15388), .I (g8898));
INVX1 gate5536(.O (I15324), .I (g8779));
INVX1 gate5537(.O (I6270), .I (g492));
INVX1 gate5538(.O (g2937), .I (g2346));
INVX1 gate5539(.O (I11870), .I (g5752));
INVX1 gate5540(.O (g7139), .I (I12999));
INVX1 gate5541(.O (g9071), .I (I15607));
INVX1 gate5542(.O (g5939), .I (I10579));
INVX1 gate5543(.O (I10705), .I (g5463));
INVX1 gate5544(.O (g6892), .I (I12547));
INVX1 gate5545(.O (g1832), .I (g763));
INVX1 gate5546(.O (g2479), .I (g32));
INVX1 gate5547(.O (g7339), .I (I13435));
INVX1 gate5548(.O (I13527), .I (g7217));
INVX1 gate5549(.O (g2668), .I (g1662));
INVX1 gate5550(.O (I14042), .I (g7470));
INVX1 gate5551(.O (g1853), .I (g766));
INVX1 gate5552(.O (g2840), .I (g2207));
INVX1 gate5553(.O (g4698), .I (I8989));
INVX1 gate5554(.O (g8775), .I (g8564));
INVX1 gate5555(.O (g3746), .I (g2100));
INVX1 gate5556(.O (g5083), .I (g4457));
INVX1 gate5557(.O (g7838), .I (I14264));
INVX1 gate5558(.O (I5879), .I (g1267));
INVX1 gate5559(.O (g7024), .I (I12782));
INVX1 gate5560(.O (g7424), .I (I13547));
INVX1 gate5561(.O (I7362), .I (g2933));
INVX1 gate5562(.O (I12909), .I (g7046));
INVX1 gate5563(.O (I14270), .I (g7703));
INVX1 gate5564(.O (g7737), .I (I14082));
INVX1 gate5565(.O (I10678), .I (g5566));
INVX1 gate5566(.O (I6124), .I (g399));
INVX1 gate5567(.O (g8581), .I (g8094));
INVX1 gate5568(.O (I14124), .I (g7591));
INVX1 gate5569(.O (g6945), .I (I12646));
INVX1 gate5570(.O (I12117), .I (g5918));
INVX1 gate5571(.O (g1794), .I (I5646));
INVX1 gate5572(.O (I11503), .I (g6220));
INVX1 gate5573(.O (g2501), .I (g27));
INVX1 gate5574(.O (I11867), .I (g6286));
INVX1 gate5575(.O (I11894), .I (g5956));
INVX1 gate5576(.O (I10460), .I (g5219));
INVX1 gate5577(.O (I13894), .I (g7353));
INVX1 gate5578(.O (g4463), .I (I8483));
INVX1 gate5579(.O (I14460), .I (g7789));
INVX1 gate5580(.O (g6244), .I (g5670));
INVX1 gate5581(.O (g7077), .I (g6676));
INVX1 gate5582(.O (I9496), .I (g3971));
INVX1 gate5583(.O (g7231), .I (I13173));
INVX1 gate5584(.O (g3932), .I (I7595));
INVX1 gate5585(.O (g5790), .I (I10415));
INVX1 gate5586(.O (g7523), .I (I13749));
INVX1 gate5587(.O (I9845), .I (g4728));
INVX1 gate5588(.O (g6140), .I (I10783));
INVX1 gate5589(.O (g3953), .I (g3160));
INVX1 gate5590(.O (g6340), .I (I11347));
INVX1 gate5591(.O (I11714), .I (g5772));
INVX1 gate5592(.O (g9350), .I (I16100));
INVX1 gate5593(.O (g5187), .I (I9687));
INVX1 gate5594(.O (g5061), .I (I9425));
INVX1 gate5595(.O (I14267), .I (g7695));
INVX1 gate5596(.O (I14294), .I (g7553));
INVX1 gate5597(.O (g6478), .I (I11638));
INVX1 gate5598(.O (g8784), .I (g8545));
INVX1 gate5599(.O (g2942), .I (g2350));
INVX1 gate5600(.O (g5461), .I (g4885));
INVX1 gate5601(.O (g4279), .I (g3340));
INVX1 gate5602(.O (I11707), .I (g5988));
INVX1 gate5603(.O (g7205), .I (I13131));
INVX1 gate5604(.O (I13707), .I (g7420));
INVX1 gate5605(.O (I13819), .I (g7426));
INVX1 gate5606(.O (g5756), .I (I10343));
INVX1 gate5607(.O (g6035), .I (g5494));
INVX1 gate5608(.O (g6959), .I (I12678));
INVX1 gate5609(.O (I7728), .I (g3675));
INVX1 gate5610(.O (I11257), .I (g5805));
INVX1 gate5611(.O (g5622), .I (g4938));
INVX1 gate5612(.O (g4619), .I (I8772));
INVX1 gate5613(.O (g5027), .I (I9369));
INVX1 gate5614(.O (g6517), .I (I11701));
INVX1 gate5615(.O (I11818), .I (g6276));
INVX1 gate5616(.O (g3677), .I (g2485));
INVX1 gate5617(.O (g5427), .I (g5115));
INVX1 gate5618(.O (I15871), .I (g9184));
INVX1 gate5619(.O (I11055), .I (g5696));
INVX1 gate5620(.O (I13979), .I (g7415));
INVX1 gate5621(.O (I5374), .I (g634));
INVX1 gate5622(.O (I13496), .I (g7133));
INVX1 gate5623(.O (g7742), .I (I14097));
INVX1 gate5624(.O (g4652), .I (I8871));
INVX1 gate5625(.O (g7551), .I (I13837));
INVX1 gate5626(.O (g7104), .I (I12900));
INVX1 gate5627(.O (g6876), .I (I12499));
INVX1 gate5628(.O (g7099), .I (I12885));
INVX1 gate5629(.O (g4057), .I (I7832));
INVX1 gate5630(.O (g7304), .I (I13344));
INVX1 gate5631(.O (g8668), .I (I14798));
INVX1 gate5632(.O (I11978), .I (g6186));
INVX1 gate5633(.O (I6849), .I (g368));
INVX1 gate5634(.O (g3866), .I (g2945));
INVX1 gate5635(.O (g2954), .I (g2374));
INVX1 gate5636(.O (g4457), .I (I8477));
INVX1 gate5637(.O (g7499), .I (g7258));
INVX1 gate5638(.O (I8877), .I (g4274));
INVX1 gate5639(.O (g2810), .I (g1922));
INVX1 gate5640(.O (g2363), .I (I6189));
INVX1 gate5641(.O (g6656), .I (I11948));
INVX1 gate5642(.O (g9212), .I (I15912));
INVX1 gate5643(.O (I12639), .I (g6506));
INVX1 gate5644(.O (I16151), .I (g9369));
INVX1 gate5645(.O (g3716), .I (g2522));
INVX1 gate5646(.O (g5514), .I (g4922));
INVX1 gate5647(.O (I5545), .I (g1276));
INVX1 gate5648(.O (g5403), .I (g5088));
INVX1 gate5649(.O (g5145), .I (I9561));
INVX1 gate5650(.O (g2453), .I (I6291));
INVX1 gate5651(.O (I5380), .I (g645));
INVX1 gate5652(.O (g5841), .I (I10538));
INVX1 gate5653(.O (g3848), .I (I7347));
INVX1 gate5654(.O (g1750), .I (g602));
INVX1 gate5655(.O (I6900), .I (g1866));
INVX1 gate5656(.O (I12265), .I (g6660));
INVX1 gate5657(.O (g7754), .I (I14133));
INVX1 gate5658(.O (I10160), .I (g5139));
INVX1 gate5659(.O (g5763), .I (I10366));
INVX1 gate5660(.O (I9142), .I (g4236));
INVX1 gate5661(.O (g5191), .I (g4969));
INVX1 gate5662(.O (g8156), .I (I14394));
INVX1 gate5663(.O (g3855), .I (I7368));
INVX1 gate5664(.O (I14160), .I (g7549));
INVX1 gate5665(.O (g3398), .I (I6952));
INVX1 gate5666(.O (I8928), .I (g4153));
INVX1 gate5667(.O (g7273), .I (I13255));
INVX1 gate5668(.O (I6245), .I (g142));
INVX1 gate5669(.O (I9081), .I (g4357));
INVX1 gate5670(.O (I12391), .I (g6744));
INVX1 gate5671(.O (g4598), .I (I8709));
INVX1 gate5672(.O (g6110), .I (g5335));
INVX1 gate5673(.O (g6310), .I (I11257));
INVX1 gate5674(.O (I6291), .I (g46));
INVX1 gate5675(.O (g7044), .I (g6543));
INVX1 gate5676(.O (I10617), .I (g5677));
INVX1 gate5677(.O (I15628), .I (g9001));
INVX1 gate5678(.O (g4121), .I (I7970));
INVX1 gate5679(.O (I5559), .I (g1292));
INVX1 gate5680(.O (g2157), .I (I5897));
INVX1 gate5681(.O (g7269), .I (I13247));
INVX1 gate5682(.O (g6663), .I (I11967));
INVX1 gate5683(.O (g4670), .I (I8925));
INVX1 gate5684(.O (g5159), .I (I9603));
INVX1 gate5685(.O (g4625), .I (I8790));
INVX1 gate5686(.O (g7983), .I (I14294));
INVX1 gate5687(.O (I10277), .I (g5472));
INVX1 gate5688(.O (I11018), .I (g5626));
INVX1 gate5689(.O (I13196), .I (g7008));
INVX1 gate5690(.O (I7635), .I (g3052));
INVX1 gate5691(.O (I13695), .I (g7345));
INVX1 gate5692(.O (g6824), .I (I12343));
INVX1 gate5693(.O (g7712), .I (I14015));
INVX1 gate5694(.O (g1666), .I (g1472));
INVX1 gate5695(.O (g3524), .I (g2306));
INVX1 gate5696(.O (g4253), .I (g2734));
INVX1 gate5697(.O (g2929), .I (g2327));
INVX1 gate5698(.O (g4938), .I (I9310));
INVX1 gate5699(.O (g6236), .I (I11037));
INVX1 gate5700(.O (g4813), .I (I9162));
INVX1 gate5701(.O (I12586), .I (g6643));
INVX1 gate5702(.O (g7543), .I (I13813));
INVX1 gate5703(.O (g5016), .I (I9350));
INVX1 gate5704(.O (g5757), .I (g5261));
INVX1 gate5705(.O (g8810), .I (I15068));
INVX1 gate5706(.O (g3644), .I (g2131));
INVX1 gate5707(.O (I7305), .I (g3048));
INVX1 gate5708(.O (g8363), .I (g7992));
INVX1 gate5709(.O (I15776), .I (g9127));
INVX1 gate5710(.O (I16058), .I (g9294));
INVX1 gate5711(.O (I10494), .I (g5232));
INVX1 gate5712(.O (g4909), .I (I9271));
INVX1 gate5713(.O (I12442), .I (g6542));
INVX1 gate5714(.O (I5515), .I (g567));
INVX1 gate5715(.O (I14623), .I (g7833));
INVX1 gate5716(.O (I8844), .I (g3992));
INVX1 gate5717(.O (g5522), .I (g4930));
INVX1 gate5718(.O (g5115), .I (I9505));
INVX1 gate5719(.O (g6877), .I (I12502));
INVX1 gate5720(.O (g5811), .I (I10466));
INVX1 gate5721(.O (g5642), .I (I10125));
INVX1 gate5722(.O (g2626), .I (g1571));
INVX1 gate5723(.O (g3577), .I (g2372));
INVX1 gate5724(.O (g7534), .I (I13782));
INVX1 gate5725(.O (g7729), .I (I14058));
INVX1 gate5726(.O (g3867), .I (g2946));
INVX1 gate5727(.O (I15950), .I (g9222));
INVX1 gate5728(.O (I13457), .I (g7120));
INVX1 gate5729(.O (g1655), .I (g1231));
INVX1 gate5730(.O (g6657), .I (I11951));
INVX1 gate5731(.O (I7755), .I (g3019));
INVX1 gate5732(.O (g4552), .I (g2890));
INVX1 gate5733(.O (g9062), .I (I15580));
INVX1 gate5734(.O (I11917), .I (g5897));
INVX1 gate5735(.O (g4606), .I (I8733));
INVX1 gate5736(.O (g6556), .I (I11732));
INVX1 gate5737(.O (I10418), .I (g5453));
INVX1 gate5738(.O (g6222), .I (g5654));
INVX1 gate5739(.O (I12041), .I (g5897));
INVX1 gate5740(.O (g5874), .I (I10565));
INVX1 gate5741(.O (I9001), .I (g4577));
INVX1 gate5742(.O (I14822), .I (g8649));
INVX1 gate5743(.O (g7014), .I (I12760));
INVX1 gate5744(.O (g4687), .I (I8962));
INVX1 gate5745(.O (I8966), .I (g4444));
INVX1 gate5746(.O (I12430), .I (g6432));
INVX1 gate5747(.O (I11001), .I (g5698));
INVX1 gate5748(.O (g5654), .I (g4748));
INVX1 gate5749(.O (I12493), .I (g6587));
INVX1 gate5750(.O (g7414), .I (I13527));
INVX1 gate5751(.O (I9129), .I (g4475));
INVX1 gate5752(.O (I15394), .I (g8916));
INVX1 gate5753(.O (g3975), .I (g3131));
INVX1 gate5754(.O (g6064), .I (I10681));
INVX1 gate5755(.O (g4586), .I (g2926));
INVX1 gate5756(.O (g6899), .I (g6525));
INVX1 gate5757(.O (g2683), .I (g1666));
INVX1 gate5758(.O (g6785), .I (I12226));
INVX1 gate5759(.O (I11689), .I (g5956));
INVX1 gate5760(.O (I11923), .I (g5939));
INVX1 gate5761(.O (I12340), .I (g6725));
INVX1 gate5762(.O (I12983), .I (g6930));
INVX1 gate5763(.O (g7513), .I (I13719));
INVX1 gate5764(.O (I5969), .I (g303));
INVX1 gate5765(.O (I12806), .I (g6602));
INVX1 gate5766(.O (I12684), .I (g6472));
INVX1 gate5767(.O (I7602), .I (g2562));
INVX1 gate5768(.O (g2894), .I (g2267));
INVX1 gate5769(.O (I15420), .I (g8881));
INVX1 gate5770(.O (g4570), .I (g2907));
INVX1 gate5771(.O (g4341), .I (I8308));
INVX1 gate5772(.O (g9298), .I (I16020));
INVX1 gate5773(.O (g9085), .I (I15645));
INVX1 gate5774(.O (I8814), .I (g4028));
INVX1 gate5775(.O (g1667), .I (g1481));
INVX1 gate5776(.O (g4525), .I (g2870));
INVX1 gate5777(.O (g4710), .I (I9009));
INVX1 gate5778(.O (g7178), .I (I13088));
INVX1 gate5779(.O (g2782), .I (g1616));
INVX1 gate5780(.O (g6295), .I (I11212));
INVX1 gate5781(.O (g1235), .I (I5422));
INVX1 gate5782(.O (g5612), .I (g4814));
INVX1 gate5783(.O (I12517), .I (g6613));
INVX1 gate5784(.O (g6237), .I (I11040));
INVX1 gate5785(.O (g4645), .I (I8850));
INVX1 gate5786(.O (I13157), .I (g6997));
INVX1 gate5787(.O (g2661), .I (I6454));
INVX1 gate5788(.O (g5417), .I (g5006));
INVX1 gate5789(.O (g1566), .I (g652));
INVX1 gate5790(.O (g7135), .I (I12989));
INVX1 gate5791(.O (g6844), .I (I12403));
INVX1 gate5792(.O (g7335), .I (I13425));
INVX1 gate5793(.O (I11066), .I (g5460));
INVX1 gate5794(.O (I13066), .I (g6957));
INVX1 gate5795(.O (I13231), .I (g6897));
INVX1 gate5796(.O (g7288), .I (I13296));
INVX1 gate5797(.O (g6194), .I (I10937));
INVX1 gate5798(.O (I5528), .I (g43));
INVX1 gate5799(.O (g2627), .I (g1572));
INVX1 gate5800(.O (I14118), .I (g7565));
INVX1 gate5801(.O (g5128), .I (I9528));
INVX1 gate5802(.O (I9624), .I (g4746));
INVX1 gate5803(.O (g2292), .I (I6060));
INVX1 gate5804(.O (I14022), .I (g7443));
INVX1 gate5805(.O (g6089), .I (g5317));
INVX1 gate5806(.O (I12193), .I (g6468));
INVX1 gate5807(.O (g6731), .I (I12101));
INVX1 gate5808(.O (g4607), .I (I8736));
INVX1 gate5809(.O (I8769), .I (g3999));
INVX1 gate5810(.O (I13876), .I (g7347));
INVX1 gate5811(.O (I13885), .I (g7351));
INVX1 gate5812(.O (g5542), .I (g5061));
INVX1 gate5813(.O (g7022), .I (I12776));
INVX1 gate5814(.O (g2646), .I (I6422));
INVX1 gate5815(.O (g7422), .I (I13541));
INVX1 gate5816(.O (g4659), .I (I8892));
INVX1 gate5817(.O (g7749), .I (I14118));
INVX1 gate5818(.O (g1555), .I (I5428));
INVX1 gate5819(.O (I12523), .I (g6624));
INVX1 gate5820(.O (g4358), .I (g3680));
INVX1 gate5821(.O (g1804), .I (I5664));
INVX1 gate5822(.O (I6887), .I (g2528));
INVX1 gate5823(.O (g8683), .I (g8235));
INVX1 gate5824(.O (I13854), .I (g7327));
INVX1 gate5825(.O (g6071), .I (I10694));
INVX1 gate5826(.O (g9219), .I (I15933));
INVX1 gate5827(.O (g1792), .I (g616));
INVX1 gate5828(.O (g2039), .I (g1228));
INVX1 gate5829(.O (g3061), .I (I6795));
INVX1 gate5830(.O (g3187), .I (I6860));
INVX1 gate5831(.O (g6471), .I (I11627));
INVX1 gate5832(.O (g8778), .I (I14974));
INVX1 gate5833(.O (I14276), .I (g7720));
INVX1 gate5834(.O (I14285), .I (g7625));
INVX1 gate5835(.O (g2484), .I (g45));
INVX1 gate5836(.O (g9031), .I (I15507));
INVX1 gate5837(.O (g5800), .I (I10439));
INVX1 gate5838(.O (I5410), .I (g8866));
INVX1 gate5839(.O (g3461), .I (I6959));
INVX1 gate5840(.O (g6242), .I (I11047));
INVX1 gate5841(.O (I14305), .I (g7537));
INVX1 gate5842(.O (g9252), .I (I15982));
INVX1 gate5843(.O (g4587), .I (g2928));
INVX1 gate5844(.O (I12475), .I (g6596));
INVX1 gate5845(.O (I6033), .I (g3));
INVX1 gate5846(.O (I9576), .I (g4706));
INVX1 gate5847(.O (I10466), .I (g5221));
INVX1 gate5848(.O (g6948), .I (I12655));
INVX1 gate5849(.O (g4111), .I (I7944));
INVX1 gate5850(.O (I5839), .I (g1198));
INVX1 gate5851(.O (g7560), .I (I13854));
INVX1 gate5852(.O (g4275), .I (g3790));
INVX1 gate5853(.O (g4311), .I (I8282));
INVX1 gate5854(.O (g9376), .I (I16154));
INVX1 gate5855(.O (I15738), .I (g9079));
INVX1 gate5856(.O (I15562), .I (g8979));
INVX1 gate5857(.O (I15645), .I (g9043));
INVX1 gate5858(.O (g6955), .I (I12666));
INVX1 gate5859(.O (g4615), .I (I8760));
INVX1 gate5860(.O (g3904), .I (g3160));
INVX1 gate5861(.O (g8661), .I (I14777));
INVX1 gate5862(.O (I10177), .I (g4721));
INVX1 gate5863(.O (I15699), .I (g9061));
INVX1 gate5864(.O (I6096), .I (g521));
INVX1 gate5865(.O (g6254), .I (g5683));
INVX1 gate5866(.O (g6814), .I (I12313));
INVX1 gate5867(.O (g7095), .I (I12877));
INVX1 gate5868(.O (g3514), .I (g2424));
INVX1 gate5869(.O (g2919), .I (g2311));
INVX1 gate5870(.O (g7037), .I (g6525));
INVX1 gate5871(.O (g6150), .I (g5287));
INVX1 gate5872(.O (g7495), .I (I13663));
INVX1 gate5873(.O (g1908), .I (g812));
INVX1 gate5874(.O (g7437), .I (I13570));
INVX1 gate5875(.O (g6350), .I (I11377));
INVX1 gate5876(.O (g7102), .I (I12894));
INVX1 gate5877(.O (g7208), .I (I13140));
INVX1 gate5878(.O (I6195), .I (g405));
INVX1 gate5879(.O (g7302), .I (I13338));
INVX1 gate5880(.O (I13550), .I (g1173));
INVX1 gate5881(.O (g6038), .I (I10649));
INVX1 gate5882(.O (I5667), .I (g916));
INVX1 gate5883(.O (I11314), .I (g5781));
INVX1 gate5884(.O (I6337), .I (g1348));
INVX1 gate5885(.O (g3841), .I (I7326));
INVX1 gate5886(.O (I13314), .I (g7160));
INVX1 gate5887(.O (I11287), .I (g5806));
INVX1 gate5888(.O (g2276), .I (I6029));
INVX1 gate5889(.O (I12253), .I (g6427));
INVX1 gate5890(.O (g6773), .I (I12190));
INVX1 gate5891(.O (I13287), .I (g7157));
INVX1 gate5892(.O (g1567), .I (g655));
INVX1 gate5893(.O (I16103), .I (g9339));
INVX1 gate5894(.O (g7579), .I (I13882));
INVX1 gate5895(.O (I14064), .I (g7556));
INVX1 gate5896(.O (g6009), .I (I10605));
INVX1 gate5897(.O (g3191), .I (I6868));
INVX1 gate5898(.O (g4545), .I (g2887));
INVX1 gate5899(.O (g2616), .I (g1564));
INVX1 gate5900(.O (g7719), .I (g7475));
INVX1 gate5901(.O (g2561), .I (g1555));
INVX1 gate5902(.O (g5490), .I (g4917));
INVX1 gate5903(.O (g691), .I (I5389));
INVX1 gate5904(.O (g5823), .I (I10494));
INVX1 gate5905(.O (g534), .I (I5365));
INVX1 gate5906(.O (g5166), .I (I9624));
INVX1 gate5907(.O (I11596), .I (g6228));
INVX1 gate5908(.O (g4591), .I (g2937));
INVX1 gate5909(.O (g8603), .I (I14674));
INVX1 gate5910(.O (I13054), .I (g6960));
INVX1 gate5911(.O (g8039), .I (g7696));
INVX1 gate5912(.O (g1776), .I (g608));
INVX1 gate5913(.O (g6769), .I (I12176));
INVX1 gate5914(.O (g7752), .I (I14127));
INVX1 gate5915(.O (I11431), .I (g5782));
INVX1 gate5916(.O (g9073), .I (I15613));
INVX1 gate5917(.O (g6836), .I (I12379));
INVX1 gate5918(.O (g4020), .I (I7781));
INVX1 gate5919(.O (g6212), .I (I10973));
INVX1 gate5920(.O (g2404), .I (g1276));
INVX1 gate5921(.O (I5548), .I (g1280));
INVX1 gate5922(.O (I8895), .I (g4130));
INVX1 gate5923(.O (g2647), .I (I6425));
INVX1 gate5924(.O (g5529), .I (g4689));
INVX1 gate5925(.O (g3159), .I (I6856));
INVX1 gate5926(.O (I10166), .I (g5016));
INVX1 gate5927(.O (g5148), .I (I9570));
INVX1 gate5928(.O (g3359), .I (I6946));
INVX1 gate5929(.O (g5649), .I (g4748));
INVX1 gate5930(.O (g6918), .I (I12609));
INVX1 gate5931(.O (g6967), .I (I12696));
INVX1 gate5932(.O (I5555), .I (g1288));
INVX1 gate5933(.O (I11269), .I (g5756));
INVX1 gate5934(.O (I14166), .I (g7702));
INVX1 gate5935(.O (I14009), .I (g7436));
INVX1 gate5936(.O (g2764), .I (g1802));
INVX1 gate5937(.O (g7265), .I (g7077));
INVX1 gate5938(.O (g9324), .I (I16072));
INVX1 gate5939(.O (g7042), .I (g6543));
INVX1 gate5940(.O (g2546), .I (I6368));
INVX1 gate5941(.O (I11773), .I (g6262));
INVX1 gate5942(.O (g5155), .I (I9591));
INVX1 gate5943(.O (g4559), .I (g2898));
INVX1 gate5944(.O (g9069), .I (I15601));
INVX1 gate5945(.O (I11942), .I (g6015));
INVX1 gate5946(.O (I11341), .I (g5809));
INVX1 gate5947(.O (I13773), .I (g7496));
INVX1 gate5948(.O (g3858), .I (I7377));
INVX1 gate5949(.O (g7442), .I (I13583));
INVX1 gate5950(.O (g8583), .I (I14668));
INVX1 gate5951(.O (I13341), .I (g7207));
INVX1 gate5952(.O (g4931), .I (I9301));
INVX1 gate5953(.O (I6248), .I (g411));
INVX1 gate5954(.O (I7564), .I (g2752));
INVX1 gate5955(.O (I9258), .I (g4249));
INVX1 gate5956(.O (g3757), .I (g1977));
INVX1 gate5957(.O (g2970), .I (g2394));
INVX1 gate5958(.O (g6229), .I (g5665));
INVX1 gate5959(.O (I15481), .I (g8913));
INVX1 gate5960(.O (I10485), .I (g5229));
INVX1 gate5961(.O (g6993), .I (I12731));
INVX1 gate5962(.O (g1933), .I (g1247));
INVX1 gate5963(.O (g7164), .I (I13066));
INVX1 gate5964(.O (g7364), .I (I13506));
INVX1 gate5965(.O (I6081), .I (g118));
INVX1 gate5966(.O (g2925), .I (g2324));
INVX1 gate5967(.O (g9177), .I (I15811));
INVX1 gate5968(.O (g7233), .I (g6940));
INVX1 gate5969(.O (g9206), .I (g9196));
INVX1 gate5970(.O (I10555), .I (g5529));
INVX1 gate5971(.O (I10454), .I (g5217));
INVX1 gate5972(.O (g6822), .I (I12337));
INVX1 gate5973(.O (g3522), .I (g2407));
INVX1 gate5974(.O (I14454), .I (g8177));
INVX1 gate5975(.O (g7054), .I (g6511));
INVX1 gate5976(.O (g2224), .I (I5945));
INVX1 gate5977(.O (g3642), .I (I7118));
INVX1 gate5978(.O (I13734), .I (g7422));
INVX1 gate5979(.O (g3047), .I (g1736));
INVX1 gate5980(.O (I10914), .I (g5448));
INVX1 gate5981(.O (I11335), .I (g5839));
INVX1 gate5982(.O (g7454), .I (I13610));
INVX1 gate5983(.O (g4628), .I (I8799));
INVX1 gate5984(.O (I14712), .I (g8059));
INVX1 gate5985(.O (I13335), .I (g7206));
INVX1 gate5986(.O (g7770), .I (I14181));
INVX1 gate5987(.O (g5463), .I (g5085));
INVX1 gate5988(.O (I6154), .I (g122));
INVX1 gate5989(.O (g7296), .I (I13320));
INVX1 gate5990(.O (I6354), .I (g1357));
INVX1 gate5991(.O (g4630), .I (I8805));
INVX1 gate5992(.O (I13930), .I (g7405));
INVX1 gate5993(.O (g7725), .I (I14046));
INVX1 gate5994(.O (I11838), .I (g6281));
INVX1 gate5995(.O (I5908), .I (g196));
INVX1 gate5996(.O (g4300), .I (I8261));
INVX1 gate5997(.O (g7532), .I (I13776));
INVX1 gate5998(.O (g1724), .I (I5568));
INVX1 gate5999(.O (I7308), .I (g3074));
INVX1 gate6000(.O (g3874), .I (g2957));
INVX1 gate6001(.O (I12208), .I (g6496));
INVX1 gate6002(.O (I13131), .I (g6951));
INVX1 gate6003(.O (g3654), .I (g2521));
INVX1 gate6004(.O (g9199), .I (g9188));
INVX1 gate6005(.O (I15784), .I (g9125));
INVX1 gate6006(.O (g8647), .I (I14739));
INVX1 gate6007(.O (I15956), .I (g9216));
INVX1 gate6008(.O (g2617), .I (g1565));
INVX1 gate6009(.O (g2906), .I (g2288));
INVX1 gate6010(.O (I15385), .I (g8880));
INVX1 gate6011(.O (g1878), .I (g80));
INVX1 gate6012(.O (g5167), .I (I9627));
INVX1 gate6013(.O (I14238), .I (g7608));
INVX1 gate6014(.O (g5367), .I (I9834));
INVX1 gate6015(.O (g5872), .I (I10561));
INVX1 gate6016(.O (I13487), .I (g7129));
AN2X1 gate6017(.O (g7412), .I1 (g7121), .I2 (g4841));
AN2X1 gate6018(.O (g6462), .I1 (g6215), .I2 (g2424));
AN2X1 gate6019(.O (g8925), .I1 (g4592), .I2 (g8754));
AN2X1 gate6020(.O (g4969), .I1 (g4362), .I2 (g2216));
AN2X1 gate6021(.O (g7429), .I1 (g1057), .I2 (g7212));
AN2X1 gate6022(.O (g9144), .I1 (g9123), .I2 (g6096));
AN2X1 gate6023(.O (g9344), .I1 (g9329), .I2 (g6211));
AN2X1 gate6024(.O (g4123), .I1 (g2627), .I2 (g2617));
AN2X1 gate6025(.O (g8320), .I1 (g4557), .I2 (g7951));
AN4X1 gate6026(.O (I8431), .I1 (g3430), .I2 (g3398), .I3 (g3359), .I4 (g3341));
AN2X1 gate6027(.O (g9259), .I1 (g9230), .I2 (g5639));
AN2X1 gate6028(.O (g8277), .I1 (g162), .I2 (g8042));
AN4X1 gate6029(.O (I8005), .I1 (g3430), .I2 (g3398), .I3 (g3359), .I4 (g2106));
AN2X1 gate6030(.O (g4351), .I1 (g309), .I2 (g3131));
AN2X1 gate6031(.O (g8299), .I1 (g591), .I2 (g8181));
AN2X1 gate6032(.O (g6941), .I1 (g1126), .I2 (g6582));
AN2X1 gate6033(.O (g4410), .I1 (g408), .I2 (g3160));
AN2X1 gate6034(.O (g8892), .I1 (g8681), .I2 (g4969));
AN4X1 gate6035(.O (I7994), .I1 (g3430), .I2 (g3398), .I3 (g3359), .I4 (g3341));
AN2X1 gate6036(.O (g5552), .I1 (g1114), .I2 (g4832));
AN2X1 gate6037(.O (g8945), .I1 (g4541), .I2 (g8784));
AN2X1 gate6038(.O (g8738), .I1 (g8619), .I2 (g3338));
AN2X1 gate6039(.O (g6431), .I1 (g5847), .I2 (g5494));
AN2X1 gate6040(.O (g4172), .I1 (I8057), .I2 (I8058));
AN2X1 gate6041(.O (g7449), .I1 (g7272), .I2 (g6901));
AN2X1 gate6042(.O (g8709), .I1 (g2818), .I2 (g8386));
AN2X1 gate6043(.O (g6176), .I1 (g1149), .I2 (g5198));
AN2X1 gate6044(.O (g6005), .I1 (g5557), .I2 (g2407));
AN2X1 gate6045(.O (g4343), .I1 (g306), .I2 (g3131));
AN2X1 gate6046(.O (g8078), .I1 (g7463), .I2 (g7634));
AN2X1 gate6047(.O (g8340), .I1 (g423), .I2 (g7920));
AN2X1 gate6048(.O (g6405), .I1 (g5956), .I2 (g5494));
AN2X1 gate6049(.O (g4282), .I1 (g3549), .I2 (g3568));
AN2X1 gate6050(.O (g7604), .I1 (g7456), .I2 (g3466));
AN2X1 gate6051(.O (g1714), .I1 (g1454), .I2 (g1450));
AN2X1 gate6052(.O (g5570), .I1 (g1759), .I2 (g4841));
AN2X1 gate6053(.O (g8690), .I1 (g3485), .I2 (g8363));
AN2X1 gate6054(.O (g7833), .I1 (g6461), .I2 (g7601));
AN2X1 gate6055(.O (g4334), .I1 (g225), .I2 (g3097));
AN2X1 gate6056(.O (g8876), .I1 (g8769), .I2 (g6102));
AN2X1 gate6057(.O (g6733), .I1 (g685), .I2 (g5873));
AN2X1 gate6058(.O (g6974), .I1 (g3613), .I2 (g6505));
AN2X1 gate6059(.O (g4804), .I1 (g952), .I2 (g3876));
AN2X1 gate6060(.O (g8915), .I1 (g8794), .I2 (g8239));
AN2X1 gate6061(.O (g7419), .I1 (g7230), .I2 (g3530));
AN2X1 gate6062(.O (g8310), .I1 (g573), .I2 (g8181));
AN2X1 gate6063(.O (g4494), .I1 (I8546), .I2 (I8547));
AN2X1 gate6064(.O (g8824), .I1 (g264), .I2 (g8524));
AN2X1 gate6065(.O (g8877), .I1 (g8773), .I2 (g6104));
AN2X1 gate6066(.O (g6399), .I1 (g5971), .I2 (g5494));
AN3X1 gate6067(.O (I9330), .I1 (g2784), .I2 (g2770), .I3 (g2746));
AN2X1 gate6068(.O (g9142), .I1 (g9124), .I2 (g6059));
AN2X1 gate6069(.O (g8928), .I1 (g4595), .I2 (g8757));
AN2X1 gate6070(.O (g5020), .I1 (g579), .I2 (g3937));
AN4X1 gate6071(.O (g4933), .I1 (g2746), .I2 (g2728), .I3 (g4320), .I4 (g2770));
AN2X1 gate6072(.O (g8930), .I1 (g3866), .I2 (g8760));
AN4X1 gate6073(.O (I8114), .I1 (g2162), .I2 (g2149), .I3 (g2137), .I4 (g2106));
AN2X1 gate6074(.O (g8064), .I1 (g7483), .I2 (g7634));
AN2X1 gate6075(.O (g7678), .I1 (g7367), .I2 (g4158));
AN2X1 gate6076(.O (g4724), .I1 (g828), .I2 (g4038));
AN2X1 gate6077(.O (g7087), .I1 (g6440), .I2 (g5311));
AN2X1 gate6078(.O (g4379), .I1 (g399), .I2 (g3160));
AN2X1 gate6079(.O (g8295), .I1 (g4512), .I2 (g7905));
AN2X1 gate6080(.O (g8237), .I1 (g89), .I2 (g8131));
AN2X1 gate6081(.O (g6923), .I1 (g6570), .I2 (g5612));
AN3X1 gate6082(.O (g4878), .I1 (g2573), .I2 (g2562), .I3 (I9222));
AN2X1 gate6083(.O (g8844), .I1 (g4056), .I2 (g8602));
AN4X1 gate6084(.O (I8594), .I1 (g3316), .I2 (g2057), .I3 (g2020), .I4 (g1987));
AN3X1 gate6085(.O (I9166), .I1 (g4041), .I2 (g2595), .I3 (g2584));
AN2X1 gate6086(.O (g8089), .I1 (g840), .I2 (g7658));
AN2X1 gate6087(.O (g8731), .I1 (g2743), .I2 (g8421));
AN2X1 gate6088(.O (g4271), .I1 (g3666), .I2 (g3684));
AN2X1 gate6089(.O (g6951), .I1 (g5511), .I2 (g6595));
AN2X1 gate6090(.O (g8071), .I1 (g7540), .I2 (g4969));
AN2X1 gate6091(.O (g8705), .I1 (g2798), .I2 (g8421));
AN2X1 gate6092(.O (g4799), .I1 (g951), .I2 (g4596));
AN4X1 gate6093(.O (I8033), .I1 (g3430), .I2 (g3398), .I3 (g3359), .I4 (g2106));
AN2X1 gate6094(.O (g8948), .I1 (g4570), .I2 (g8789));
AN2X1 gate6095(.O (g5969), .I1 (g5564), .I2 (g2424));
AN2X1 gate6096(.O (g7602), .I1 (g7476), .I2 (g3466));
AN2X1 gate6097(.O (g7007), .I1 (g6627), .I2 (g5072));
AN2X1 gate6098(.O (g5123), .I1 (g516), .I2 (g4033));
AN2X1 gate6099(.O (g4132), .I1 (g2637), .I2 (g2633));
AN4X1 gate6100(.O (I8496), .I1 (g3316), .I2 (g3287), .I3 (g2020), .I4 (g1987));
AN3X1 gate6101(.O (g4238), .I1 (g2695), .I2 (g2698), .I3 (I8157));
AN2X1 gate6102(.O (g8814), .I1 (g3880), .I2 (g8463));
AN2X1 gate6103(.O (g6408), .I1 (g669), .I2 (g6019));
AN2X1 gate6104(.O (g8150), .I1 (g846), .I2 (g7658));
AN2X1 gate6105(.O (g4744), .I1 (g3525), .I2 (g4296));
AN2X1 gate6106(.O (g8438), .I1 (g649), .I2 (g7793));
AN2X1 gate6107(.O (g6972), .I1 (g5661), .I2 (g6498));
AN2X1 gate6108(.O (g7415), .I1 (g7222), .I2 (g5603));
AN2X1 gate6109(.O (g8836), .I1 (g348), .I2 (g8545));
AN3X1 gate6110(.O (g4901), .I1 (g3723), .I2 (g4288), .I3 (I9261));
AN2X1 gate6111(.O (g6433), .I1 (g778), .I2 (g6134));
AN2X1 gate6112(.O (g8229), .I1 (g8180), .I2 (g5680));
AN2X1 gate6113(.O (g9349), .I1 (g9340), .I2 (g5690));
AN2X1 gate6114(.O (g8822), .I1 (g417), .I2 (g8564));
AN2X1 gate6115(.O (g6395), .I1 (g2157), .I2 (g6007));
AN2X1 gate6116(.O (g8921), .I1 (g4579), .I2 (g8747));
AN2X1 gate6117(.O (g7689), .I1 (g7367), .I2 (g4417));
AN2X1 gate6118(.O (g5334), .I1 (g4887), .I2 (g2424));
AN2X1 gate6119(.O (g5548), .I1 (g1549), .I2 (g4826));
AN2X1 gate6120(.O (g4968), .I1 (g4403), .I2 (g1760));
AN2X1 gate6121(.O (g6266), .I1 (g1481), .I2 (g5285));
AN2X1 gate6122(.O (g8837), .I1 (g426), .I2 (g8564));
AN2X1 gate6123(.O (g7030), .I1 (g6705), .I2 (g5723));
AN2X1 gate6124(.O (g8062), .I1 (g7476), .I2 (g7634));
AN2X1 gate6125(.O (g8620), .I1 (g751), .I2 (g8199));
AN2X1 gate6126(.O (g8462), .I1 (g49), .I2 (g8199));
AN2X1 gate6127(.O (g9119), .I1 (g9049), .I2 (g5345));
AN4X1 gate6128(.O (I8001), .I1 (g2074), .I2 (g3287), .I3 (g2020), .I4 (g1987));
AN2X1 gate6129(.O (g7564), .I1 (g7367), .I2 (g4172));
AN2X1 gate6130(.O (g9258), .I1 (g9227), .I2 (g5628));
AN4X1 gate6131(.O (I8401), .I1 (g3316), .I2 (g3287), .I3 (g3264), .I4 (g3238));
AN2X1 gate6132(.O (g4175), .I1 (g1110), .I2 (g3502));
AN2X1 gate6133(.O (g4375), .I1 (g219), .I2 (g3097));
AN2X1 gate6134(.O (g5313), .I1 (g4820), .I2 (g2407));
AN2X1 gate6135(.O (g6726), .I1 (g5897), .I2 (g5367));
AN2X1 gate6136(.O (g6154), .I1 (g1499), .I2 (g5713));
AN2X1 gate6137(.O (g8842), .I1 (g429), .I2 (g8564));
AN2X1 gate6138(.O (g7609), .I1 (g7467), .I2 (g3466));
AN2X1 gate6139(.O (g8298), .I1 (g553), .I2 (g8181));
AN2X1 gate6140(.O (g5094), .I1 (g535), .I2 (g4004));
AN2X1 gate6141(.O (g9274), .I1 (g4748), .I2 (g9255));
AN2X1 gate6142(.O (g4139), .I1 (I8000), .I2 (I8001));
AN2X1 gate6143(.O (g4384), .I1 (g246), .I2 (g3097));
AN2X1 gate6144(.O (g4838), .I1 (g4517), .I2 (g1760));
AN2X1 gate6145(.O (g8854), .I1 (g443), .I2 (g8564));
AN2X1 gate6146(.O (g7217), .I1 (g1142), .I2 (g6941));
AN2X1 gate6147(.O (g8941), .I1 (g3882), .I2 (g8776));
AN2X1 gate6148(.O (g4424), .I1 (g489), .I2 (g3192));
AN2X1 gate6149(.O (g6979), .I1 (g5095), .I2 (g6511));
AN2X1 gate6150(.O (g5593), .I1 (g4110), .I2 (g4969));
AN3X1 gate6151(.O (g6112), .I1 (g5673), .I2 (g4841), .I3 (g5541));
AN2X1 gate6152(.O (g4077), .I1 (g1284), .I2 (g3582));
AN2X1 gate6153(.O (g6001), .I1 (g5540), .I2 (g2407));
AN2X1 gate6154(.O (g6401), .I1 (g5971), .I2 (g5367));
AN2X1 gate6155(.O (g8708), .I1 (g3557), .I2 (g8407));
AN2X1 gate6156(.O (g7827), .I1 (g7575), .I2 (g7173));
AN2X1 gate6157(.O (g5050), .I1 (g587), .I2 (g3970));
AN2X1 gate6158(.O (g1725), .I1 (g1409), .I2 (g1416));
AN2X1 gate6159(.O (g6727), .I1 (g681), .I2 (g5846));
AN2X1 gate6160(.O (g8405), .I1 (g741), .I2 (g8018));
AN2X1 gate6161(.O (g4099), .I1 (g117), .I2 (g3647));
AN2X1 gate6162(.O (g4304), .I1 (g2784), .I2 (g3779));
AN2X1 gate6163(.O (g8829), .I1 (g267), .I2 (g8524));
AN2X1 gate6164(.O (g8286), .I1 (g180), .I2 (g8156));
AN2X1 gate6165(.O (g8911), .I1 (g8798), .I2 (g7688));
AN2X1 gate6166(.O (g8733), .I1 (g2996), .I2 (g8493));
AN2X1 gate6167(.O (g8270), .I1 (g110), .I2 (g8131));
AN2X1 gate6168(.O (g8610), .I1 (g665), .I2 (g7887));
AN2X1 gate6169(.O (g9345), .I1 (g9330), .I2 (g6217));
AN3X1 gate6170(.O (g4269), .I1 (g2354), .I2 (g3563), .I3 (I8209));
AN4X1 gate6171(.O (I8524), .I1 (g3316), .I2 (g2057), .I3 (g3264), .I4 (g1987));
AN2X1 gate6172(.O (g2781), .I1 (g1600), .I2 (g976));
AN2X1 gate6173(.O (g8069), .I1 (g7456), .I2 (g7634));
AN2X1 gate6174(.O (g4712), .I1 (g1179), .I2 (g4276));
AN2X1 gate6175(.O (g7181), .I1 (g6124), .I2 (g7039));
AN2X1 gate6176(.O (g9159), .I1 (g9138), .I2 (g6074));
AN2X1 gate6177(.O (g9359), .I1 (g4748), .I2 (g9340));
AN2X1 gate6178(.O (g8377), .I1 (g507), .I2 (g7966));
AN2X1 gate6179(.O (g7197), .I1 (g7093), .I2 (g5055));
AN2X1 gate6180(.O (g7700), .I1 (g7367), .I2 (g4494));
AN2X1 gate6181(.O (g7021), .I1 (g3390), .I2 (g6673));
AN2X1 gate6182(.O (g4729), .I1 (g1504), .I2 (g4059));
AN2X1 gate6183(.O (g4961), .I1 (g377), .I2 (g3904));
AN2X1 gate6184(.O (g9016), .I1 (g8904), .I2 (g8239));
AN2X1 gate6185(.O (g8287), .I1 (g4500), .I2 (g7855));
AN4X1 gate6186(.O (I8186), .I1 (g3778), .I2 (g3549), .I3 (g3568), .I4 (g3583));
AN2X1 gate6187(.O (g5132), .I1 (I9534), .I2 (I9535));
AN2X1 gate6188(.O (g8849), .I1 (g513), .I2 (g8585));
AN4X1 gate6189(.O (I7995), .I1 (g2074), .I2 (g3287), .I3 (g2020), .I4 (g3238));
AN2X1 gate6190(.O (g9251), .I1 (g4748), .I2 (g9230));
AN2X1 gate6191(.O (g4414), .I1 (I8412), .I2 (I8413));
AN3X1 gate6192(.O (g3313), .I1 (g2334), .I2 (g2316), .I3 (g2298));
AN2X1 gate6193(.O (g7631), .I1 (g7367), .I2 (g4187));
AN2X1 gate6194(.O (g8291), .I1 (g122), .I2 (g8111));
AN2X1 gate6195(.O (g3094), .I1 (g945), .I2 (g1898));
AN2X1 gate6196(.O (g4436), .I1 (g492), .I2 (g3192));
AN2X1 gate6197(.O (g6577), .I1 (g6142), .I2 (g4160));
AN2X1 gate6198(.O (g7605), .I1 (g7435), .I2 (g5607));
AN2X1 gate6199(.O (g4378), .I1 (g321), .I2 (g3131));
AN2X1 gate6200(.O (g4135), .I1 (I7994), .I2 (I7995));
AN2X1 gate6201(.O (g5092), .I1 (g456), .I2 (g4002));
AN2X1 gate6202(.O (g4182), .I1 (I8071), .I2 (I8072));
AN4X1 gate6203(.O (g4288), .I1 (g3563), .I2 (g3579), .I3 (g3603), .I4 (I8240));
AN2X1 gate6204(.O (g9272), .I1 (g4748), .I2 (g9248));
AN2X1 gate6205(.O (g8259), .I1 (g4538), .I2 (g7855));
AN2X1 gate6206(.O (g5714), .I1 (g1532), .I2 (g4733));
AN2X1 gate6207(.O (g8088), .I1 (g837), .I2 (g7658));
AN2X1 gate6208(.O (g8852), .I1 (g362), .I2 (g8545));
AN2X1 gate6209(.O (g8923), .I1 (g4587), .I2 (g8751));
AN4X1 gate6210(.O (I8461), .I1 (g3316), .I2 (g3287), .I3 (g2020), .I4 (g3238));
AN2X1 gate6211(.O (g7041), .I1 (g6734), .I2 (g5206));
AN2X1 gate6212(.O (g4422), .I1 (g411), .I2 (g3160));
AN2X1 gate6213(.O (g8701), .I1 (g2700), .I2 (g8363));
AN2X1 gate6214(.O (g2768), .I1 (g1597), .I2 (g973));
AN2X1 gate6215(.O (g9328), .I1 (g9324), .I2 (g6465));
AN2X1 gate6216(.O (g4798), .I1 (g4216), .I2 (g1760));
AN2X1 gate6217(.O (g9130), .I1 (g9054), .I2 (g5345));
AN2X1 gate6218(.O (g6125), .I1 (g5548), .I2 (g4202));
AN2X1 gate6219(.O (g2972), .I1 (g2397), .I2 (g2407));
AN4X1 gate6220(.O (I8046), .I1 (g2074), .I2 (g2057), .I3 (g3264), .I4 (g1987));
AN2X1 gate6221(.O (g8951), .I1 (g8785), .I2 (g6072));
AN2X1 gate6222(.O (g8314), .I1 (g443), .I2 (g7920));
AN2X1 gate6223(.O (g4437), .I1 (g540), .I2 (g2845));
AN2X1 gate6224(.O (g8825), .I1 (g342), .I2 (g8545));
AN2X1 gate6225(.O (g8650), .I1 (g591), .I2 (g8094));
AN3X1 gate6226(.O (g4302), .I1 (g3086), .I2 (g3659), .I3 (g3124));
AN2X1 gate6227(.O (g1728), .I1 (g1432), .I2 (g1439));
AN2X1 gate6228(.O (g8336), .I1 (g420), .I2 (g7920));
AN2X1 gate6229(.O (g6061), .I1 (g5257), .I2 (g1616));
AN2X1 gate6230(.O (g8943), .I1 (g4560), .I2 (g8781));
AN2X1 gate6231(.O (g6046), .I1 (g1073), .I2 (g5592));
AN4X1 gate6232(.O (I8115), .I1 (g2074), .I2 (g3287), .I3 (g3264), .I4 (g1987));
AN4X1 gate6233(.O (I8642), .I1 (g3430), .I2 (g3398), .I3 (g3359), .I4 (g2106));
AN2X1 gate6234(.O (g8322), .I1 (g4559), .I2 (g7993));
AN3X1 gate6235(.O (g6003), .I1 (g3716), .I2 (g5633), .I3 (I10597));
AN2X1 gate6236(.O (g8934), .I1 (g3873), .I2 (g8766));
AN2X1 gate6237(.O (g9348), .I1 (g9333), .I2 (g6229));
AN2X1 gate6238(.O (g7713), .I1 (g4403), .I2 (g7367));
AN2X1 gate6239(.O (g6145), .I1 (g1489), .I2 (g5705));
AN2X1 gate6240(.O (g4054), .I1 (g3767), .I2 (g2424));
AN2X1 gate6241(.O (g4454), .I1 (g544), .I2 (g2845));
AN2X1 gate6242(.O (g5077), .I1 (g236), .I2 (g3988));
AN2X1 gate6243(.O (g4532), .I1 (I8617), .I2 (I8618));
AN2X1 gate6244(.O (g6107), .I1 (g5478), .I2 (g1849));
AN2X1 gate6245(.O (g8845), .I1 (g432), .I2 (g8564));
AN3X1 gate6246(.O (I9202), .I1 (g2605), .I2 (g4044), .I3 (g2584));
AN2X1 gate6247(.O (g8337), .I1 (g498), .I2 (g7966));
AN2X1 gate6248(.O (g4412), .I1 (g486), .I2 (g3192));
AN2X1 gate6249(.O (g5104), .I1 (g274), .I2 (g4010));
AN2X1 gate6250(.O (g6757), .I1 (g5874), .I2 (g5412));
AN2X1 gate6251(.O (g9279), .I1 (g9255), .I2 (g5665));
AN2X1 gate6252(.O (g4389), .I1 (g480), .I2 (g3192));
AN4X1 gate6253(.O (I8612), .I1 (g3430), .I2 (g3398), .I3 (g3359), .I4 (g3341));
AN2X1 gate6254(.O (g6416), .I1 (g710), .I2 (g6026));
AN4X1 gate6255(.O (I8417), .I1 (g3430), .I2 (g3398), .I3 (g3359), .I4 (g2106));
AN2X1 gate6256(.O (g9118), .I1 (g9046), .I2 (g5345));
AN2X1 gate6257(.O (g4787), .I1 (g953), .I2 (g4547));
AN2X1 gate6258(.O (g6047), .I1 (g1477), .I2 (g5596));
AN2X1 gate6259(.O (g8266), .I1 (g2157), .I2 (g8042));
AN2X1 gate6260(.O (g6447), .I1 (g734), .I2 (g6073));
AN2X1 gate6261(.O (g4956), .I1 (g295), .I2 (g3892));
AN2X1 gate6262(.O (g2979), .I1 (g1494), .I2 (g1733));
AN2X1 gate6263(.O (g5044), .I1 (g234), .I2 (g3959));
AN2X1 gate6264(.O (g8081), .I1 (g834), .I2 (g7658));
AN2X1 gate6265(.O (g8815), .I1 (g258), .I2 (g8524));
AN2X1 gate6266(.O (g7183), .I1 (g6132), .I2 (g7042));
AN2X1 gate6267(.O (g7608), .I1 (g7367), .I2 (g4169));
AN2X1 gate6268(.O (g8692), .I1 (g3462), .I2 (g8363));
AN2X1 gate6269(.O (g8726), .I1 (g2795), .I2 (g8386));
AN2X1 gate6270(.O (g4138), .I1 (g2638), .I2 (g2634));
AN2X1 gate6271(.O (g4109), .I1 (g990), .I2 (g3790));
AN2X1 gate6272(.O (g4791), .I1 (g949), .I2 (g4562));
AN2X1 gate6273(.O (g4707), .I1 (g812), .I2 (g4062));
AN2X1 gate6274(.O (g6417), .I1 (g718), .I2 (g6027));
AN4X1 gate6275(.O (I8090), .I1 (g3316), .I2 (g2057), .I3 (g2020), .I4 (g3238));
AN4X1 gate6276(.O (I8490), .I1 (g3430), .I2 (g3398), .I3 (g3359), .I4 (g3341));
AN2X1 gate6277(.O (g4201), .I1 (I8108), .I2 (I8109));
AN2X1 gate6278(.O (g8267), .I1 (g154), .I2 (g8042));
AN2X1 gate6279(.O (g8312), .I1 (g365), .I2 (g7870));
AN2X1 gate6280(.O (g6629), .I1 (g6023), .I2 (g4841));
AN3X1 gate6281(.O (g4957), .I1 (g2746), .I2 (g2728), .I3 (g4320));
AN2X1 gate6282(.O (g4049), .I1 (g141), .I2 (g3514));
AN4X1 gate6283(.O (I8456), .I1 (g3316), .I2 (g3287), .I3 (g2020), .I4 (g1987));
AN4X1 gate6284(.O (I8529), .I1 (g3316), .I2 (g2057), .I3 (g3264), .I4 (g3238));
AN2X1 gate6285(.O (g8293), .I1 (g4510), .I2 (g7855));
AN2X1 gate6286(.O (g8329), .I1 (g527), .I2 (g7966));
AN2X1 gate6287(.O (g7696), .I1 (g7367), .I2 (g4469));
AN2X1 gate6288(.O (g5513), .I1 (g4889), .I2 (g5071));
AN2X1 gate6289(.O (g4098), .I1 (g985), .I2 (g3790));
AN2X1 gate6290(.O (g6554), .I1 (g5762), .I2 (g1616));
AN2X1 gate6291(.O (g8828), .I1 (g4573), .I2 (g8541));
AN2X1 gate6292(.O (g8830), .I1 (g345), .I2 (g8545));
AN2X1 gate6293(.O (g8727), .I1 (g2724), .I2 (g8421));
AN2X1 gate6294(.O (g5436), .I1 (g1541), .I2 (g4926));
AN2X1 gate6295(.O (g7240), .I1 (g6719), .I2 (g6894));
AN4X1 gate6296(.O (I8063), .I1 (g2162), .I2 (g2149), .I3 (g2137), .I4 (g2106));
AN2X1 gate6297(.O (g8703), .I1 (g3574), .I2 (g8407));
AN2X1 gate6298(.O (g4268), .I1 (g2216), .I2 (g2655));
AN2X1 gate6299(.O (g8932), .I1 (g3868), .I2 (g8762));
AN2X1 gate6300(.O (g6166), .I1 (g1509), .I2 (g5725));
AN2X1 gate6301(.O (g8624), .I1 (g754), .I2 (g8199));
AN2X1 gate6302(.O (g8953), .I1 (g8758), .I2 (g6093));
AN2X1 gate6303(.O (g4052), .I1 (g1276), .I2 (g3522));
AN2X1 gate6304(.O (g8068), .I1 (g7687), .I2 (g5610));
AN2X1 gate6305(.O (g4452), .I1 (g437), .I2 (g3160));
AN3X1 gate6306(.O (g6056), .I1 (g3760), .I2 (g5286), .I3 (g1695));
AN2X1 gate6307(.O (g6456), .I1 (g6116), .I2 (g2407));
AN4X1 gate6308(.O (I8057), .I1 (g3430), .I2 (g3398), .I3 (g3359), .I4 (g3341));
AN2X1 gate6309(.O (g7681), .I1 (g7444), .I2 (g5099));
AN2X1 gate6310(.O (g9158), .I1 (g9137), .I2 (g6070));
AN2X1 gate6311(.O (g5560), .I1 (g3390), .I2 (g5036));
AN2X1 gate6312(.O (g4086), .I1 (g103), .I2 (g3629));
AN2X1 gate6313(.O (g4728), .I1 (g190), .I2 (g4179));
AN2X1 gate6314(.O (g4486), .I1 (I8528), .I2 (I8529));
AN2X1 gate6315(.O (g8716), .I1 (g3506), .I2 (g8443));
AN2X1 gate6316(.O (g7596), .I1 (g7428), .I2 (g7028));
AN2X1 gate6317(.O (g4504), .I1 (I8568), .I2 (I8569));
AN2X1 gate6318(.O (g4185), .I1 (g2636), .I2 (g2632));
AN2X1 gate6319(.O (g9275), .I1 (g9241), .I2 (g5645));
AN2X1 gate6320(.O (g4385), .I1 (g300), .I2 (g3131));
AN2X1 gate6321(.O (g8848), .I1 (g281), .I2 (g8524));
AN2X1 gate6322(.O (g5579), .I1 (g4090), .I2 (g4841));
AN2X1 gate6323(.O (g4425), .I1 (g536), .I2 (g2845));
AN2X1 gate6324(.O (g2386), .I1 (g1130), .I2 (g1092));
AN2X1 gate6325(.O (g5442), .I1 (g4679), .I2 (g4202));
AN2X1 gate6326(.O (g6057), .I1 (g1061), .I2 (g5617));
AN2X1 gate6327(.O (g4131), .I1 (g2630), .I2 (g2622));
AN2X1 gate6328(.O (g8319), .I1 (g255), .I2 (g7838));
AN4X1 gate6329(.O (I8552), .I1 (g3316), .I2 (g2057), .I3 (g3264), .I4 (g1987));
AN2X1 gate6330(.O (g8258), .I1 (g142), .I2 (g8111));
AN2X1 gate6331(.O (g6971), .I1 (g6424), .I2 (g4969));
AN2X1 gate6332(.O (g8717), .I1 (g2764), .I2 (g8421));
AN2X1 gate6333(.O (g7597), .I1 (g7316), .I2 (g4841));
AN2X1 gate6334(.O (g7079), .I1 (g4259), .I2 (g6677));
AN2X1 gate6335(.O (g8274), .I1 (g4580), .I2 (g7951));
AN2X1 gate6336(.O (g4445), .I1 (I8455), .I2 (I8456));
AN2X1 gate6337(.O (g4091), .I1 (g129), .I2 (g3639));
AN2X1 gate6338(.O (g4491), .I1 (g557), .I2 (g2845));
AN2X1 gate6339(.O (g8325), .I1 (g184), .I2 (g8156));
AN2X1 gate6340(.O (g8821), .I1 (g339), .I2 (g8545));
AN2X1 gate6341(.O (g4169), .I1 (I8052), .I2 (I8053));
AN2X1 gate6342(.O (g5029), .I1 (g212), .I2 (g3945));
AN2X1 gate6343(.O (g4369), .I1 (g580), .I2 (g2845));
AN2X1 gate6344(.O (g8280), .I1 (g114), .I2 (g8111));
AN2X1 gate6345(.O (g8939), .I1 (g3879), .I2 (g8772));
AN2X1 gate6346(.O (g4407), .I1 (g252), .I2 (g3097));
AN2X1 gate6347(.O (g4059), .I1 (g1499), .I2 (g2979));
AN2X1 gate6348(.O (g4868), .I1 (g4227), .I2 (g4160));
AN2X1 gate6349(.O (g8306), .I1 (g4525), .I2 (g7951));
AN2X1 gate6350(.O (g4793), .I1 (g3887), .I2 (g4202));
AN2X1 gate6351(.O (g8461), .I1 (g658), .I2 (g7793));
AN2X1 gate6352(.O (g8622), .I1 (g738), .I2 (g7811));
AN2X1 gate6353(.O (g4246), .I1 (g1106), .I2 (g3226));
AN2X1 gate6354(.O (g8403), .I1 (g639), .I2 (g7793));
AN2X1 gate6355(.O (g8841), .I1 (g351), .I2 (g8545));
AN2X1 gate6356(.O (g5049), .I1 (g474), .I2 (g3969));
AN4X1 gate6357(.O (I8020), .I1 (g2074), .I2 (g3287), .I3 (g2020), .I4 (g1987));
AN2X1 gate6358(.O (g8695), .I1 (g2709), .I2 (g8363));
AN2X1 gate6359(.O (g8307), .I1 (g432), .I2 (g7920));
AN2X1 gate6360(.O (g9278), .I1 (g9252), .I2 (g5658));
AN2X1 gate6361(.O (g4388), .I1 (g402), .I2 (g3160));
AN2X1 gate6362(.O (g8359), .I1 (g642), .I2 (g7793));
AN2X1 gate6363(.O (g4216), .I1 (I8114), .I2 (I8115));
AN2X1 gate6364(.O (g9143), .I1 (g9122), .I2 (g6089));
AN2X1 gate6365(.O (g9343), .I1 (g9328), .I2 (g1738));
AN2X1 gate6366(.O (g7626), .I1 (g7463), .I2 (g3466));
AN2X1 gate6367(.O (g8858), .I1 (g524), .I2 (g8585));
AN2X1 gate6368(.O (g4430), .I1 (I8436), .I2 (I8437));
AN4X1 gate6369(.O (I9534), .I1 (g3019), .I2 (g3029), .I3 (g3038), .I4 (g3052));
AN2X1 gate6370(.O (g9334), .I1 (g9318), .I2 (g6205));
AN2X1 gate6371(.O (g8315), .I1 (g4544), .I2 (g7993));
AN2X1 gate6372(.O (g4826), .I1 (g1545), .I2 (g4239));
AN2X1 gate6373(.O (g6239), .I1 (g1514), .I2 (g5314));
AN2X1 gate6374(.O (g5019), .I1 (g312), .I2 (g3933));
AN2X1 gate6375(.O (g2935), .I1 (g1612), .I2 (g1077));
AN2X1 gate6376(.O (g7683), .I1 (g1061), .I2 (g7429));
AN2X1 gate6377(.O (g5452), .I1 (g4876), .I2 (g3499));
AN2X1 gate6378(.O (g8654), .I1 (g570), .I2 (g8094));
AN2X1 gate6379(.O (g6420), .I1 (g5918), .I2 (g5367));
AN2X1 gate6380(.O (g4108), .I1 (g782), .I2 (g3655));
AN3X1 gate6381(.O (g4883), .I1 (g3746), .I2 (g3723), .I3 (g4288));
AN4X1 gate6382(.O (I8040), .I1 (g3430), .I2 (g3398), .I3 (g3359), .I4 (g3341));
AN2X1 gate6383(.O (g4066), .I1 (g1280), .I2 (g3532));
AN2X1 gate6384(.O (g8272), .I1 (g158), .I2 (g8042));
AN2X1 gate6385(.O (g4466), .I1 (I8490), .I2 (I8491));
AN2X1 gate6386(.O (g8978), .I1 (g8909), .I2 (g5587));
AN2X1 gate6387(.O (g8612), .I1 (g673), .I2 (g7887));
AN3X1 gate6388(.O (g3429), .I1 (g1454), .I2 (g1838), .I3 (g1444));
AN2X1 gate6389(.O (g6204), .I1 (g5542), .I2 (g5294));
AN2X1 gate6390(.O (g4365), .I1 (g237), .I2 (g3097));
AN2X1 gate6391(.O (g4048), .I1 (g1288), .I2 (g3513));
AN2X1 gate6392(.O (g8935), .I1 (g3874), .I2 (g8767));
AN2X1 gate6393(.O (g5425), .I1 (g1528), .I2 (g4916));
AN2X1 gate6394(.O (g4448), .I1 (I8460), .I2 (I8461));
AN2X1 gate6395(.O (g4711), .I1 (g190), .I2 (g4072));
AN4X1 gate6396(.O (I8528), .I1 (g3430), .I2 (g3398), .I3 (g3359), .I4 (g2106));
AN2X1 gate6397(.O (g8328), .I1 (g4571), .I2 (g7993));
AN2X1 gate6398(.O (g4133), .I1 (g2631), .I2 (g2623));
AN2X1 gate6399(.O (g4333), .I1 (g1087), .I2 (g2782));
AN2X1 gate6400(.O (g8542), .I1 (g661), .I2 (g7887));
AN2X1 gate6401(.O (g8330), .I1 (g261), .I2 (g7838));
AN2X1 gate6402(.O (g4396), .I1 (g459), .I2 (g3192));
AN2X1 gate6403(.O (g9160), .I1 (g9139), .I2 (g6092));
AN2X1 gate6404(.O (g6040), .I1 (g1462), .I2 (g5578));
AN2X1 gate6405(.O (g5105), .I1 (g354), .I2 (g4013));
AN2X1 gate6406(.O (g7616), .I1 (g7367), .I2 (g4517));
AN2X1 gate6407(.O (g7561), .I1 (g7367), .I2 (g4163));
AN2X1 gate6408(.O (g4067), .I1 (g133), .I2 (g3539));
AN4X1 gate6409(.O (I8618), .I1 (g2074), .I2 (g3287), .I3 (g3264), .I4 (g3238));
AN3X1 gate6410(.O (I8143), .I1 (g2674), .I2 (g2677), .I3 (g2680));
AN2X1 gate6411(.O (g3049), .I1 (g2274), .I2 (g1844));
AN2X1 gate6412(.O (g8090), .I1 (g843), .I2 (g7658));
AN2X1 gate6413(.O (g6151), .I1 (g1494), .I2 (g5709));
AN2X1 gate6414(.O (g8823), .I1 (g4561), .I2 (g8512));
AN2X1 gate6415(.O (g5045), .I1 (g293), .I2 (g3961));
AN2X1 gate6416(.O (g5091), .I1 (g397), .I2 (g4001));
AN2X1 gate6417(.O (g4181), .I1 (g1142), .I2 (g3512));
AN2X1 gate6418(.O (g8456), .I1 (g703), .I2 (g7811));
AN2X1 gate6419(.O (g9271), .I1 (g4748), .I2 (g9244));
AN2X1 gate6420(.O (g4397), .I1 (g483), .I2 (g3192));
AN2X1 gate6421(.O (g8851), .I1 (g284), .I2 (g8524));
AN2X1 gate6422(.O (g4421), .I1 (g333), .I2 (g3131));
AN2X1 gate6423(.O (g8698), .I1 (g3774), .I2 (g8342));
AN2X1 gate6424(.O (g8260), .I1 (g138), .I2 (g8111));
AN2X1 gate6425(.O (g5767), .I1 (g5344), .I2 (g3079));
AN2X1 gate6426(.O (g6172), .I1 (g1514), .I2 (g5192));
AN2X1 gate6427(.O (g9238), .I1 (g4748), .I2 (g9223));
AN2X1 gate6428(.O (g8720), .I1 (g3825), .I2 (g8421));
AN2X1 gate6429(.O (g4101), .I1 (g108), .I2 (g3649));
AN2X1 gate6430(.O (g8318), .I1 (g183), .I2 (g8156));
AN2X1 gate6431(.O (g8652), .I1 (g563), .I2 (g8094));
AN2X1 gate6432(.O (g8843), .I1 (g507), .I2 (g8585));
AN4X1 gate6433(.O (I8593), .I1 (g3430), .I2 (g3398), .I3 (g3359), .I4 (g2106));
AN2X1 gate6434(.O (g8457), .I1 (g724), .I2 (g7811));
AN3X1 gate6435(.O (I10597), .I1 (g3769), .I2 (g3754), .I3 (g3735));
AN2X1 gate6436(.O (g1753), .I1 (g819), .I2 (g815));
AN2X1 gate6437(.O (g8686), .I1 (g3819), .I2 (g8342));
AN2X1 gate6438(.O (g7709), .I1 (g7367), .I2 (g4529));
AN2X1 gate6439(.O (g8321), .I1 (g446), .I2 (g7920));
AN2X1 gate6440(.O (g6908), .I1 (g6478), .I2 (g5246));
AN2X1 gate6441(.O (g4168), .I1 (g1106), .I2 (g3500));
AN2X1 gate6442(.O (g6567), .I1 (g6265), .I2 (g2424));
AN2X1 gate6443(.O (g4368), .I1 (g318), .I2 (g3131));
AN2X1 gate6444(.O (g8938), .I1 (g3878), .I2 (g8771));
AN2X1 gate6445(.O (g5428), .I1 (g775), .I2 (g4707));
AN2X1 gate6446(.O (g8813), .I1 (g255), .I2 (g8524));
AN2X1 gate6447(.O (g5030), .I1 (g233), .I2 (g3946));
AN2X1 gate6448(.O (g4058), .I1 (g3656), .I2 (g2407));
AN2X1 gate6449(.O (g4743), .I1 (g3518), .I2 (g4286));
AN2X1 gate6450(.O (g8740), .I1 (g2966), .I2 (g8493));
AN2X1 gate6451(.O (g6965), .I1 (g55), .I2 (g6489));
AN2X1 gate6452(.O (g4411), .I1 (g462), .I2 (g3192));
AN2X1 gate6453(.O (g8687), .I1 (g3488), .I2 (g8363));
AN2X1 gate6454(.O (g6160), .I1 (g1504), .I2 (g5718));
AN2X1 gate6455(.O (g3226), .I1 (g1102), .I2 (g1919));
AN2X1 gate6456(.O (g4074), .I1 (g137), .I2 (g3573));
AN2X1 gate6457(.O (g5108), .I1 (g539), .I2 (g4017));
AN2X1 gate6458(.O (g6641), .I1 (g5939), .I2 (g5494));
AN2X1 gate6459(.O (g7002), .I1 (g6770), .I2 (g5054));
AN2X1 gate6460(.O (g6996), .I1 (g3678), .I2 (g6552));
AN2X1 gate6461(.O (g5066), .I1 (g395), .I2 (g3978));
AN2X1 gate6462(.O (g8860), .I1 (g527), .I2 (g8585));
AN2X1 gate6463(.O (g8341), .I1 (g501), .I2 (g7966));
AN2X1 gate6464(.O (g8710), .I1 (g2790), .I2 (g8421));
AN2X1 gate6465(.O (g9384), .I1 (g9383), .I2 (g6245));
AN2X1 gate6466(.O (g8645), .I1 (g550), .I2 (g8094));
AN3X1 gate6467(.O (I8209), .I1 (g2298), .I2 (g2316), .I3 (g2334));
AN2X1 gate6468(.O (g7657), .I1 (g7367), .I2 (g4201));
AN2X1 gate6469(.O (g8691), .I1 (g3805), .I2 (g8342));
AN2X1 gate6470(.O (g5048), .I1 (g394), .I2 (g3966));
AN2X1 gate6471(.O (g9024), .I1 (g8884), .I2 (g5317));
AN2X1 gate6472(.O (g8879), .I1 (g8782), .I2 (g6108));
AN2X1 gate6473(.O (g8607), .I1 (g8154), .I2 (g5616));
AN2X1 gate6474(.O (g8962), .I1 (g8890), .I2 (g5317));
AN2X1 gate6475(.O (g6611), .I1 (g3390), .I2 (g6249));
AN2X1 gate6476(.O (g1739), .I1 (g803), .I2 (g799));
AN2X1 gate6477(.O (g8275), .I1 (g4581), .I2 (g7993));
AN2X1 gate6478(.O (g8311), .I1 (g4540), .I2 (g7905));
AN2X1 gate6479(.O (g4400), .I1 (g1138), .I2 (g3614));
AN2X1 gate6480(.O (g6541), .I1 (g6144), .I2 (g3510));
AN4X1 gate6481(.O (I8574), .I1 (g3316), .I2 (g2057), .I3 (g2020), .I4 (g3238));
AN2X1 gate6482(.O (g5018), .I1 (g232), .I2 (g3930));
AN2X1 gate6483(.O (g5067), .I1 (g454), .I2 (g3980));
AN2X1 gate6484(.O (g5093), .I1 (g477), .I2 (g4003));
AN2X1 gate6485(.O (g9273), .I1 (g4748), .I2 (g9252));
AN2X1 gate6486(.O (g7557), .I1 (g7367), .I2 (g4147));
AN2X1 gate6487(.O (g4383), .I1 (g222), .I2 (g3097));
AN4X1 gate6488(.O (g4220), .I1 (g3533), .I2 (g3549), .I3 (g3568), .I4 (g3583));
AN2X1 gate6489(.O (g8380), .I1 (g681), .I2 (g7887));
AN2X1 gate6490(.O (g8832), .I1 (g501), .I2 (g8585));
AN2X1 gate6491(.O (g7071), .I1 (g6639), .I2 (g1872));
AN2X1 gate6492(.O (g4779), .I1 (g4176), .I2 (g1760));
AN2X1 gate6493(.O (g7705), .I1 (g7367), .I2 (g4514));
AN2X1 gate6494(.O (g8853), .I1 (g365), .I2 (g8545));
AN2X1 gate6495(.O (g7242), .I1 (g7081), .I2 (g6899));
AN2X1 gate6496(.O (g4423), .I1 (g465), .I2 (g3192));
AN2X1 gate6497(.O (g3188), .I1 (g2298), .I2 (g2316));
AN2X1 gate6498(.O (g5700), .I1 (g1638), .I2 (g4969));
AN2X1 gate6499(.O (g4361), .I1 (g471), .I2 (g3192));
AN2X1 gate6500(.O (g8931), .I1 (g3867), .I2 (g8761));
AN2X1 gate6501(.O (g4127), .I1 (g2628), .I2 (g2618));
AN2X1 gate6502(.O (g4451), .I1 (g359), .I2 (g3131));
AN2X1 gate6503(.O (g4327), .I1 (g2959), .I2 (g1867));
AN2X1 gate6504(.O (g6574), .I1 (g1045), .I2 (g5984));
AN2X1 gate6505(.O (g7038), .I1 (g6466), .I2 (g4841));
AN2X1 gate6506(.O (g8628), .I1 (g753), .I2 (g8199));
AN2X1 gate6507(.O (g8300), .I1 (g126), .I2 (g8111));
AN2X1 gate6508(.O (g9014), .I1 (g8906), .I2 (g8239));
AN2X1 gate6509(.O (g7212), .I1 (g1053), .I2 (g7010));
AN2X1 gate6510(.O (g5817), .I1 (g5395), .I2 (g3091));
AN2X1 gate6511(.O (g4472), .I1 (g440), .I2 (g3160));
AN2X1 gate6512(.O (g3466), .I1 (g936), .I2 (g2557));
AN2X1 gate6513(.O (g8440), .I1 (g714), .I2 (g7937));
AN4X1 gate6514(.O (I8523), .I1 (g3430), .I2 (g3398), .I3 (g3359), .I4 (g3341));
AN2X1 gate6515(.O (g5585), .I1 (g4741), .I2 (g4841));
AN4X1 gate6516(.O (I8643), .I1 (g2074), .I2 (g3287), .I3 (g3264), .I4 (g1987));
AN4X1 gate6517(.O (I9535), .I1 (g3062), .I2 (g2712), .I3 (g4253), .I4 (g2752));
AN2X1 gate6518(.O (g6175), .I1 (g4332), .I2 (g5614));
AN2X1 gate6519(.O (g8323), .I1 (g524), .I2 (g7966));
AN2X1 gate6520(.O (g9335), .I1 (g9320), .I2 (g6206));
AN2X1 gate6521(.O (g5441), .I1 (g4870), .I2 (g3497));
AN2X1 gate6522(.O (g4434), .I1 (g356), .I2 (g3131));
AN3X1 gate6523(.O (I9261), .I1 (g3777), .I2 (g3764), .I3 (g3746));
AN2X1 gate6524(.O (g4147), .I1 (I8014), .I2 (I8015));
AN4X1 gate6525(.O (I8551), .I1 (g3430), .I2 (g3398), .I3 (g3359), .I4 (g2106));
AN2X1 gate6526(.O (g9022), .I1 (g8887), .I2 (g5317));
AN2X1 gate6527(.O (g4681), .I1 (g4255), .I2 (g3533));
AN2X1 gate6528(.O (g8151), .I1 (g849), .I2 (g7658));
AN2X1 gate6529(.O (g8648), .I1 (g588), .I2 (g8094));
AN2X1 gate6530(.O (g7837), .I1 (g6470), .I2 (g7610));
AN2X1 gate6531(.O (g5458), .I1 (g4686), .I2 (g1616));
AN2X1 gate6532(.O (g3509), .I1 (g1637), .I2 (g1616));
AN4X1 gate6533(.O (I8613), .I1 (g2074), .I2 (g3287), .I3 (g3264), .I4 (g1987));
AN2X1 gate6534(.O (g8839), .I1 (g4050), .I2 (g8581));
AN2X1 gate6535(.O (g9037), .I1 (g8965), .I2 (g5345));
AN2X1 gate6536(.O (g6643), .I1 (g1860), .I2 (g5868));
AN2X1 gate6537(.O (g4936), .I1 (g214), .I2 (g3888));
AN2X1 gate6538(.O (g4117), .I1 (g2626), .I2 (g2616));
AN4X1 gate6539(.O (g4317), .I1 (g878), .I2 (g3086), .I3 (g1857), .I4 (g3659));
AN2X1 gate6540(.O (g8278), .I1 (g4589), .I2 (g7993));
AN2X1 gate6541(.O (g7192), .I1 (g7026), .I2 (g3526));
AN2X1 gate6542(.O (g8282), .I1 (g179), .I2 (g8156));
AN2X1 gate6543(.O (g5080), .I1 (g396), .I2 (g3991));
AN2X1 gate6544(.O (g5573), .I1 (g3011), .I2 (g4841));
AN2X1 gate6545(.O (g8693), .I1 (g3798), .I2 (g8342));
AN2X1 gate6546(.O (g8334), .I1 (g264), .I2 (g7838));
AN4X1 gate6547(.O (I8014), .I1 (g3430), .I2 (g3398), .I3 (g3359), .I4 (g3341));
AN2X1 gate6548(.O (g1919), .I1 (g1098), .I2 (g1087));
AN2X1 gate6549(.O (g6044), .I1 (g1467), .I2 (g5584));
AN2X1 gate6550(.O (g7031), .I1 (g3390), .I2 (g6717));
AN2X1 gate6551(.O (g6444), .I1 (g1676), .I2 (g6125));
AN2X1 gate6552(.O (g7252), .I1 (g3591), .I2 (g6977));
AN2X1 gate6553(.O (g8621), .I1 (g734), .I2 (g7937));
AN2X1 gate6554(.O (g4937), .I1 (g3086), .I2 (g4309));
AN2X1 gate6555(.O (g8313), .I1 (g4542), .I2 (g7951));
AN2X1 gate6556(.O (g4840), .I1 (g4235), .I2 (g1980));
AN4X1 gate6557(.O (I8436), .I1 (g3430), .I2 (g3398), .I3 (g3359), .I4 (g2106));
AN2X1 gate6558(.O (g4190), .I1 (g1122), .I2 (g3527));
AN2X1 gate6559(.O (g4390), .I1 (g560), .I2 (g2845));
AN2X1 gate6560(.O (g5126), .I1 (g556), .I2 (g4037));
AN2X1 gate6561(.O (g9012), .I1 (g8908), .I2 (g8239));
AN3X1 gate6562(.O (I8288), .I1 (g3666), .I2 (g3684), .I3 (g3694));
AN2X1 gate6563(.O (g4356), .I1 (g468), .I2 (g3192));
AN2X1 gate6564(.O (g9371), .I1 (g9352), .I2 (g5917));
AN2X1 gate6565(.O (g6414), .I1 (g673), .I2 (g6025));
AN2X1 gate6566(.O (g8264), .I1 (g105), .I2 (g8131));
AN2X1 gate6567(.O (g4163), .I1 (I8040), .I2 (I8041));
AN2X1 gate6568(.O (g8933), .I1 (g4511), .I2 (g8765));
AN2X1 gate6569(.O (g7177), .I1 (g7016), .I2 (g5586));
AN2X1 gate6570(.O (g4053), .I1 (g1292), .I2 (g3523));
AN2X1 gate6571(.O (g5588), .I1 (g3028), .I2 (g4969));
AN2X1 gate6572(.O (g4453), .I1 (g495), .I2 (g3192));
AN4X1 gate6573(.O (I8495), .I1 (g3430), .I2 (g3398), .I3 (g3359), .I4 (g2106));
AN4X1 gate6574(.O (I8437), .I1 (g3316), .I2 (g3287), .I3 (g3264), .I4 (g1987));
AN2X1 gate6575(.O (g6182), .I1 (g1519), .I2 (g5199));
AN2X1 gate6576(.O (g8724), .I1 (g3822), .I2 (g8464));
AN2X1 gate6577(.O (g8379), .I1 (g691), .I2 (g7793));
AN2X1 gate6578(.O (g7199), .I1 (g1467), .I2 (g7003));
AN2X1 gate6579(.O (g6916), .I1 (g727), .I2 (g6515));
AN2X1 gate6580(.O (g6022), .I1 (g5595), .I2 (g2424));
AN2X1 gate6581(.O (g8878), .I1 (g8777), .I2 (g6106));
AN2X1 gate6582(.O (g6422), .I1 (g714), .I2 (g6033));
AN2X1 gate6583(.O (g8289), .I1 (g348), .I2 (g7870));
AN2X1 gate6584(.O (g8835), .I1 (g270), .I2 (g8524));
AN2X1 gate6585(.O (g8271), .I1 (g130), .I2 (g8111));
AN2X1 gate6586(.O (g8611), .I1 (g669), .I2 (g7887));
AN2X1 gate6587(.O (g5043), .I1 (g213), .I2 (g3958));
AN3X1 gate6588(.O (I8296), .I1 (g3666), .I2 (g3684), .I3 (g3707));
AN2X1 gate6589(.O (g6437), .I1 (g859), .I2 (g6050));
AN2X1 gate6590(.O (g5443), .I1 (g1549), .I2 (g4935));
AN2X1 gate6591(.O (g7694), .I1 (g7367), .I2 (g4448));
AN2X1 gate6592(.O (g5116), .I1 (g355), .I2 (g4021));
AN2X1 gate6593(.O (g8238), .I1 (g100), .I2 (g8131));
AN2X1 gate6594(.O (g5034), .I1 (g583), .I2 (g3956));
AN2X1 gate6595(.O (g8332), .I1 (g417), .I2 (g7920));
AN2X1 gate6596(.O (g7701), .I1 (g7367), .I2 (g4497));
AN2X1 gate6597(.O (g8153), .I1 (g852), .I2 (g7658));
AN2X1 gate6598(.O (g4778), .I1 (g4169), .I2 (g1760));
AN2X1 gate6599(.O (g8744), .I1 (g3802), .I2 (g8464));
AN2X1 gate6600(.O (g7215), .I1 (g6111), .I2 (g6984));
AN4X1 gate6601(.O (I8412), .I1 (g3430), .I2 (g3398), .I3 (g3359), .I4 (g3341));
AN2X1 gate6602(.O (g4782), .I1 (g4187), .I2 (g1760));
AN2X1 gate6603(.O (g6042), .I1 (g1041), .I2 (g5581));
AN4X1 gate6604(.O (I8029), .I1 (g2074), .I2 (g2057), .I3 (g3264), .I4 (g1987));
AN2X1 gate6605(.O (g8901), .I1 (g8804), .I2 (g5631));
AN2X1 gate6606(.O (g6054), .I1 (g1057), .I2 (g5611));
AN2X1 gate6607(.O (g4526), .I1 (g2642), .I2 (g741));
AN2X1 gate6608(.O (g7008), .I1 (g6615), .I2 (g5083));
AN2X1 gate6609(.O (g2889), .I1 (g1612), .I2 (g1077));
AN2X1 gate6610(.O (g7136), .I1 (g4057), .I2 (g6953));
AN2X1 gate6611(.O (g5117), .I1 (g435), .I2 (g4024));
AN2X1 gate6612(.O (g8714), .I1 (g2873), .I2 (g8407));
AN2X1 gate6613(.O (g9025), .I1 (g8889), .I2 (g5317));
AN4X1 gate6614(.O (I8109), .I1 (g2074), .I2 (g3287), .I3 (g3264), .I4 (g3238));
AN2X1 gate6615(.O (g4702), .I1 (g4243), .I2 (g1690));
AN2X1 gate6616(.O (g6412), .I1 (g158), .I2 (g6024));
AN2X1 gate6617(.O (g7228), .I1 (g6688), .I2 (g7090));
AN2X1 gate6618(.O (g6990), .I1 (g799), .I2 (g6517));
AN2X1 gate6619(.O (g8262), .I1 (g4554), .I2 (g7855));
AN2X1 gate6620(.O (g6171), .I1 (g5363), .I2 (g4841));
AN2X1 gate6621(.O (g8736), .I1 (g3771), .I2 (g8464));
AN2X1 gate6622(.O (g4276), .I1 (g2216), .I2 (g2618));
AN2X1 gate6623(.O (g6429), .I1 (g168), .I2 (g6035));
AN2X1 gate6624(.O (g7033), .I1 (g6716), .I2 (g5190));
AN2X1 gate6625(.O (g9131), .I1 (g9055), .I2 (g5345));
AN2X1 gate6626(.O (g8623), .I1 (g755), .I2 (g8199));
AN2X1 gate6627(.O (g8076), .I1 (g7690), .I2 (g3521));
AN2X1 gate6628(.O (g7096), .I1 (g6677), .I2 (g5101));
AN2X1 gate6629(.O (g8722), .I1 (g2787), .I2 (g8386));
AN2X1 gate6630(.O (g7195), .I1 (g6984), .I2 (g4226));
AN2X1 gate6631(.O (g1844), .I1 (g792), .I2 (g795));
AN2X1 gate6632(.O (g5937), .I1 (g5562), .I2 (g2407));
AN2X1 gate6633(.O (g5079), .I1 (g375), .I2 (g3990));
AN2X1 gate6634(.O (g4546), .I1 (g2643), .I2 (g746));
AN2X1 gate6635(.O (g5479), .I1 (g5141), .I2 (g5037));
AN2X1 gate6636(.O (g6745), .I1 (g1872), .I2 (g6198));
AN2X1 gate6637(.O (g8285), .I1 (g118), .I2 (g8111));
AN2X1 gate6638(.O (g9226), .I1 (g9220), .I2 (g5403));
AN2X1 gate6639(.O (g6109), .I1 (g5453), .I2 (g5335));
AN3X1 gate6640(.O (g4224), .I1 (g2680), .I2 (g2683), .I3 (I8127));
AN2X1 gate6641(.O (g8384), .I1 (g636), .I2 (g7793));
AN2X1 gate6642(.O (g8339), .I1 (g345), .I2 (g7870));
AN4X1 gate6643(.O (g4320), .I1 (g3728), .I2 (g3750), .I3 (g3768), .I4 (I8299));
AN2X1 gate6644(.O (g8838), .I1 (g504), .I2 (g8585));
AN4X1 gate6645(.O (I8019), .I1 (g3430), .I2 (g3398), .I3 (g3359), .I4 (g2106));
AN2X1 gate6646(.O (g8737), .I1 (g2992), .I2 (g8493));
AN4X1 gate6647(.O (I8052), .I1 (g2162), .I2 (g2149), .I3 (g2137), .I4 (g2106));
AN2X1 gate6648(.O (g4906), .I1 (g4320), .I2 (g2728));
AN2X1 gate6649(.O (g4789), .I1 (g2751), .I2 (g4202));
AN2X1 gate6650(.O (g6049), .I1 (g1045), .I2 (g5597));
AN2X1 gate6651(.O (g8077), .I1 (g859), .I2 (g7616));
AN2X1 gate6652(.O (g7692), .I1 (g7367), .I2 (g4430));
AN2X1 gate6653(.O (g8643), .I1 (g547), .I2 (g8094));
AN2X1 gate6654(.O (g6715), .I1 (g677), .I2 (g5843));
AN2X1 gate6655(.O (g6098), .I1 (g5681), .I2 (g1247));
AN2X1 gate6656(.O (g5032), .I1 (g313), .I2 (g3950));
AN2X1 gate6657(.O (g5432), .I1 (g1537), .I2 (g4921));
AN2X1 gate6658(.O (g4299), .I1 (g3233), .I2 (g3358));
AN2X1 gate6659(.O (g9015), .I1 (g8905), .I2 (g8239));
AN2X1 gate6660(.O (g8742), .I1 (g2973), .I2 (g8493));
AN2X1 gate6661(.O (g8304), .I1 (g4523), .I2 (g7905));
AN2X1 gate6662(.O (g8926), .I1 (g4593), .I2 (g8755));
AN2X1 gate6663(.O (g6162), .I1 (g1134), .I2 (g5724));
AN2X1 gate6664(.O (g6268), .I1 (g1092), .I2 (g5309));
AN2X1 gate6665(.O (g7001), .I1 (g3722), .I2 (g6562));
AN2X1 gate6666(.O (g8273), .I1 (g185), .I2 (g8156));
AN2X1 gate6667(.O (g6419), .I1 (g162), .I2 (g6032));
AN2X1 gate6668(.O (g7676), .I1 (g7367), .I2 (g4216));
AN2X1 gate6669(.O (g6052), .I1 (g1049), .I2 (g5604));
AN4X1 gate6670(.O (g4078), .I1 (g3753), .I2 (g3732), .I3 (g3712), .I4 (g3700));
AN2X1 gate6671(.O (g8269), .I1 (g4569), .I2 (g7951));
AN2X1 gate6672(.O (g4959), .I1 (g376), .I2 (g3898));
AN4X1 gate6673(.O (I8006), .I1 (g2074), .I2 (g3287), .I3 (g2020), .I4 (g3238));
AN2X1 gate6674(.O (g4435), .I1 (g414), .I2 (g3160));
AN2X1 gate6675(.O (g4517), .I1 (I8593), .I2 (I8594));
AN2X1 gate6676(.O (g4690), .I1 (g4081), .I2 (g3078));
AN2X1 gate6677(.O (g4082), .I1 (g1296), .I2 (g3604));
AN2X1 gate6678(.O (g8712), .I1 (g2804), .I2 (g8386));
AN2X1 gate6679(.O (g8543), .I1 (g706), .I2 (g7887));
AN2X1 gate6680(.O (g7703), .I1 (g7367), .I2 (g4504));
AN2X1 gate6681(.O (g8729), .I1 (g2999), .I2 (g8493));
AN2X1 gate6682(.O (g8961), .I1 (g8885), .I2 (g5317));
AN2X1 gate6683(.O (g9247), .I1 (g4748), .I2 (g9227));
AN2X1 gate6684(.O (g8927), .I1 (g4594), .I2 (g8756));
AN4X1 gate6685(.O (I8045), .I1 (g3430), .I2 (g3398), .I3 (g3359), .I4 (g2106));
AN2X1 gate6686(.O (g5894), .I1 (g1118), .I2 (g5552));
AN2X1 gate6687(.O (g8660), .I1 (g1069), .I2 (g8147));
AN2X1 gate6688(.O (g8946), .I1 (g4556), .I2 (g8786));
AN2X1 gate6689(.O (g7677), .I1 (g7503), .I2 (g5073));
AN4X1 gate6690(.O (I8491), .I1 (g3316), .I2 (g2057), .I3 (g3264), .I4 (g3238));
AN2X1 gate6691(.O (g6006), .I1 (g5575), .I2 (g2424));
AN2X1 gate6692(.O (g4236), .I1 (g3260), .I2 (g3221));
AN2X1 gate6693(.O (g8513), .I1 (g718), .I2 (g7937));
AN2X1 gate6694(.O (g6406), .I1 (g154), .I2 (g6018));
AN2X1 gate6695(.O (g5475), .I1 (g3801), .I2 (g5022));
AN2X1 gate6696(.O (g3190), .I1 (g1658), .I2 (g2424));
AN2X1 gate6697(.O (g6105), .I1 (g5618), .I2 (g2817));
AN4X1 gate6698(.O (g4877), .I1 (g3746), .I2 (g3723), .I3 (g4288), .I4 (g3764));
AN2X1 gate6699(.O (g8378), .I1 (g677), .I2 (g7887));
AN2X1 gate6700(.O (g6487), .I1 (g5750), .I2 (g4969));
AN2X1 gate6701(.O (g7699), .I1 (g7367), .I2 (g4486));
AN2X1 gate6702(.O (g8335), .I1 (g342), .I2 (g7870));
AN2X1 gate6703(.O (g8831), .I1 (g423), .I2 (g8564));
AN2X1 gate6704(.O (g8288), .I1 (g270), .I2 (g7838));
AN2X1 gate6705(.O (g8382), .I1 (g685), .I2 (g7887));
AN2X1 gate6706(.O (g5484), .I1 (g1037), .I2 (g5096));
AN4X1 gate6707(.O (I8015), .I1 (g2074), .I2 (g2057), .I3 (g3264), .I4 (g3238));
AN2X1 gate6708(.O (g8749), .I1 (g2989), .I2 (g8493));
AN2X1 gate6709(.O (g4785), .I1 (g1678), .I2 (g4202));
AN2X1 gate6710(.O (g6045), .I1 (g1472), .I2 (g5591));
AN2X1 gate6711(.O (g5583), .I1 (g1775), .I2 (g4969));
AN2X1 gate6712(.O (g6091), .I1 (g5712), .I2 (g5038));
AN2X1 gate6713(.O (g8947), .I1 (g4558), .I2 (g8787));
AN2X1 gate6714(.O (g6407), .I1 (g5956), .I2 (g5367));
AN2X1 gate6715(.O (g6578), .I1 (g6218), .I2 (g3913));
AN2X1 gate6716(.O (g4194), .I1 (I8089), .I2 (I8090));
AN2X1 gate6717(.O (g8653), .I1 (g573), .I2 (g8094));
AN2X1 gate6718(.O (g4394), .I1 (g381), .I2 (g3160));
AN2X1 gate6719(.O (g8302), .I1 (g4521), .I2 (g7855));
AN2X1 gate6720(.O (g7186), .I1 (g6600), .I2 (g7044));
AN2X1 gate6721(.O (g6582), .I1 (g1122), .I2 (g5894));
AN2X1 gate6722(.O (g1733), .I1 (g1489), .I2 (g1481));
AN2X1 gate6723(.O (g8719), .I1 (g2821), .I2 (g8443));
AN2X1 gate6724(.O (g4705), .I1 (g190), .I2 (g3986));
AN2X1 gate6725(.O (g6415), .I1 (g5988), .I2 (g5367));
AN2X1 gate6726(.O (g7614), .I1 (g7367), .I2 (g4176));
AN2X1 gate6727(.O (g5970), .I1 (g5605), .I2 (g2424));
AN4X1 gate6728(.O (I8028), .I1 (g3430), .I2 (g3398), .I3 (g3359), .I4 (g3341));
AN2X1 gate6729(.O (g8265), .I1 (g134), .I2 (g8111));
AN2X1 gate6730(.O (g4955), .I1 (g215), .I2 (g3891));
AN3X1 gate6731(.O (g4254), .I1 (g3583), .I2 (g3568), .I3 (g3549));
AN2X1 gate6732(.O (g4814), .I1 (g150), .I2 (g4265));
AN2X1 gate6733(.O (g4150), .I1 (I8019), .I2 (I8020));
AN2X1 gate6734(.O (g4038), .I1 (g825), .I2 (g2949));
AN2X1 gate6735(.O (g9021), .I1 (g8886), .I2 (g5317));
AN2X1 gate6736(.O (g8296), .I1 (g351), .I2 (g7870));
AN2X1 gate6737(.O (g4409), .I1 (g384), .I2 (g3160));
AN2X1 gate6738(.O (g8725), .I1 (g3008), .I2 (g8493));
AN4X1 gate6739(.O (I8108), .I1 (g2162), .I2 (g2149), .I3 (g2137), .I4 (g2106));
AN2X1 gate6740(.O (g6689), .I1 (g1519), .I2 (g6239));
AN2X1 gate6741(.O (g7027), .I1 (g3390), .I2 (g6698));
AN2X1 gate6742(.O (g5547), .I1 (g4814), .I2 (g1819));
AN2X1 gate6743(.O (g7427), .I1 (g1472), .I2 (g7199));
AN2X1 gate6744(.O (g1898), .I1 (g959), .I2 (g955));
AN4X1 gate6745(.O (I8589), .I1 (g2074), .I2 (g3287), .I3 (g3264), .I4 (g3238));
AN2X1 gate6746(.O (g6428), .I1 (g5874), .I2 (g5494));
AN2X1 gate6747(.O (g6430), .I1 (g5874), .I2 (g5384));
AN2X1 gate6748(.O (g7003), .I1 (g1462), .I2 (g6689));
AN4X1 gate6749(.O (I8455), .I1 (g3430), .I2 (g3398), .I3 (g3359), .I4 (g3341));
AN2X1 gate6750(.O (g7695), .I1 (g7367), .I2 (g4466));
AN2X1 gate6751(.O (g8281), .I1 (g168), .I2 (g8042));
AN2X1 gate6752(.O (g5078), .I1 (g316), .I2 (g3989));
AN2X1 gate6753(.O (g6638), .I1 (g174), .I2 (g5755));
AN2X1 gate6754(.O (g7536), .I1 (g4414), .I2 (g7367));
AN2X1 gate6755(.O (g8297), .I1 (g429), .I2 (g7920));
AN2X1 gate6756(.O (g5082), .I1 (g476), .I2 (g3994));
AN2X1 gate6757(.O (g8745), .I1 (g2982), .I2 (g8493));
AN3X1 gate6758(.O (g4837), .I1 (g2573), .I2 (g2562), .I3 (I9202));
AN2X1 gate6759(.O (g8338), .I1 (g570), .I2 (g8181));
AN2X1 gate6760(.O (g8963), .I1 (g8891), .I2 (g5317));
AN2X1 gate6761(.O (g4062), .I1 (g809), .I2 (g2986));
AN2X1 gate6762(.O (g7416), .I1 (g7140), .I2 (g4969));
AN2X1 gate6763(.O (g8309), .I1 (g550), .I2 (g8181));
AN4X1 gate6764(.O (I8418), .I1 (g3316), .I2 (g3287), .I3 (g3264), .I4 (g3238));
AN2X1 gate6765(.O (g6448), .I1 (g5918), .I2 (g5384));
AN2X1 gate6766(.O (g6055), .I1 (g5239), .I2 (g4202));
AN2X1 gate6767(.O (g7654), .I1 (g7367), .I2 (g4142));
AN2X1 gate6768(.O (g4192), .I1 (g1126), .I2 (g3531));
AN2X1 gate6769(.O (g4392), .I1 (g303), .I2 (g3131));
AN2X1 gate6770(.O (g6196), .I1 (g4927), .I2 (g5615));
AN2X1 gate6771(.O (g6396), .I1 (g661), .I2 (g6008));
AN2X1 gate6772(.O (g8715), .I1 (g2761), .I2 (g8386));
AN2X1 gate6773(.O (g7537), .I1 (g7363), .I2 (g7411));
AN2X1 gate6774(.O (g8833), .I1 (g4583), .I2 (g8562));
AN2X1 gate6775(.O (g7017), .I1 (g3390), .I2 (g6706));
AN2X1 gate6776(.O (g7417), .I1 (g7144), .I2 (g1616));
AN2X1 gate6777(.O (g8584), .I1 (g8146), .I2 (g7034));
AN2X1 gate6778(.O (g9080), .I1 (g9011), .I2 (g5598));
AN2X1 gate6779(.O (g6418), .I1 (g5897), .I2 (g5494));
AN2X1 gate6780(.O (g6994), .I1 (g3658), .I2 (g6538));
AN2X1 gate6781(.O (g7128), .I1 (g6926), .I2 (g3047));
AN2X1 gate6782(.O (g8268), .I1 (g4568), .I2 (g7905));
AN2X1 gate6783(.O (g5064), .I1 (g315), .I2 (g3975));
AN2X1 gate6784(.O (g8362), .I1 (g504), .I2 (g7966));
AN2X1 gate6785(.O (g4958), .I1 (g296), .I2 (g3897));
AN2X1 gate6786(.O (g4176), .I1 (I8063), .I2 (I8064));
AN2X1 gate6787(.O (g4376), .I1 (g243), .I2 (g3097));
AN2X1 gate6788(.O (g7554), .I1 (g7367), .I2 (g4139));
AN2X1 gate6789(.O (g5563), .I1 (g3390), .I2 (g5070));
AN2X1 gate6790(.O (g1913), .I1 (g1528), .I2 (g1532));
AN2X1 gate6791(.O (g6021), .I1 (g5594), .I2 (g2424));
AN2X1 gate6792(.O (g6421), .I1 (g5847), .I2 (g5384));
AN2X1 gate6793(.O (g8728), .I1 (g3815), .I2 (g8464));
AN2X1 gate6794(.O (g8730), .I1 (g2863), .I2 (g8407));
AN4X1 gate6795(.O (g4225), .I1 (g2686), .I2 (g2689), .I3 (g2692), .I4 (g2695));
AN2X1 gate6796(.O (g8385), .I1 (g695), .I2 (g7811));
AN4X1 gate6797(.O (I8041), .I1 (g2074), .I2 (g2057), .I3 (g2020), .I4 (g3238));
AN2X1 gate6798(.O (g4073), .I1 (g1300), .I2 (g3567));
AN2X1 gate6799(.O (g4796), .I1 (g950), .I2 (g4584));
AN2X1 gate6800(.O (g8070), .I1 (g863), .I2 (g7616));
AN2X1 gate6801(.O (g5089), .I1 (g273), .I2 (g3998));
AN2X1 gate6802(.O (g4473), .I1 (g518), .I2 (g3192));
AN2X1 gate6803(.O (g5489), .I1 (g4912), .I2 (g5053));
AN2X1 gate6804(.O (g4124), .I1 (g2641), .I2 (g2640));
AN2X1 gate6805(.O (g4469), .I1 (I8495), .I2 (I8496));
AN2X1 gate6806(.O (g4377), .I1 (g297), .I2 (g3131));
AN4X1 gate6807(.O (I8058), .I1 (g2074), .I2 (g2057), .I3 (g2020), .I4 (g1987));
AN2X1 gate6808(.O (g8331), .I1 (g339), .I2 (g7870));
AN2X1 gate6809(.O (g9023), .I1 (g8888), .I2 (g5317));
AN4X1 gate6810(.O (g4287), .I1 (g3563), .I2 (g2334), .I3 (g3579), .I4 (I8237));
AN2X1 gate6811(.O (g7698), .I1 (g7367), .I2 (g4483));
AN2X1 gate6812(.O (g8087), .I1 (g7471), .I2 (g7634));
AN2X1 gate6813(.O (g8305), .I1 (g362), .I2 (g7870));
AN2X1 gate6814(.O (g4199), .I1 (g93), .I2 (g2769));
AN2X1 gate6815(.O (g5438), .I1 (g1545), .I2 (g4932));
AN2X1 gate6816(.O (g4781), .I1 (g4182), .I2 (g1760));
AN2X1 gate6817(.O (g6041), .I1 (g5189), .I2 (g4969));
AN2X1 gate6818(.O (g8748), .I1 (g2721), .I2 (g8483));
AN2X1 gate6819(.O (g9327), .I1 (g9316), .I2 (g5757));
AN2X1 gate6820(.O (g4797), .I1 (g3893), .I2 (g1616));
AN2X1 gate6821(.O (g9146), .I1 (g9135), .I2 (g6101));
AN2X1 gate6822(.O (g9346), .I1 (g9331), .I2 (g6222));
AN2X1 gate6823(.O (g3002), .I1 (g871), .I2 (g1834));
AN4X1 gate6824(.O (I8573), .I1 (g3430), .I2 (g3398), .I3 (g3359), .I4 (g2106));
AN2X1 gate6825(.O (g6168), .I1 (g1138), .I2 (g5191));
AN2X1 gate6826(.O (g7652), .I1 (g7367), .I2 (g4194));
AN2X1 gate6827(.O (g6058), .I1 (g5561), .I2 (g3501));
AN2X1 gate6828(.O (g7193), .I1 (g6911), .I2 (g1616));
AN4X1 gate6829(.O (I8569), .I1 (g3316), .I2 (g2057), .I3 (g2020), .I4 (g1987));
AN2X1 gate6830(.O (g6743), .I1 (g730), .I2 (g5916));
AN3X1 gate6831(.O (g4819), .I1 (g2573), .I2 (g2562), .I3 (I9166));
AN2X1 gate6832(.O (g8283), .I1 (g267), .I2 (g7838));
AN2X1 gate6833(.O (g9240), .I1 (g9223), .I2 (g5261));
AN2X1 gate6834(.O (g8059), .I1 (g7682), .I2 (g7032));
AN2X1 gate6835(.O (g8920), .I1 (g4578), .I2 (g8746));
AN2X1 gate6836(.O (g8459), .I1 (g655), .I2 (g7793));
AN2X1 gate6837(.O (g6411), .I1 (g5918), .I2 (g5494));
AN2X1 gate6838(.O (g8718), .I1 (g2774), .I2 (g8386));
AN2X1 gate6839(.O (g7598), .I1 (g7483), .I2 (g3466));
AN2X1 gate6840(.O (g3222), .I1 (g1537), .I2 (g1913));
AN2X1 gate6841(.O (g8261), .I1 (g174), .I2 (g8042));
AN2X1 gate6842(.O (g6474), .I1 (g6203), .I2 (g2424));
AN2X1 gate6843(.O (g7625), .I1 (g7367), .I2 (g4182));
AN2X1 gate6844(.O (g8793), .I1 (g8637), .I2 (g5622));
AN2X1 gate6845(.O (g6992), .I1 (g6610), .I2 (g3519));
AN2X1 gate6846(.O (g7232), .I1 (g6694), .I2 (g7091));
AN4X1 gate6847(.O (I8000), .I1 (g3430), .I2 (g3398), .I3 (g3359), .I4 (g3341));
AN3X1 gate6848(.O (g4314), .I1 (g3694), .I2 (g3684), .I3 (g3666));
AN4X1 gate6849(.O (I8400), .I1 (g3430), .I2 (g3398), .I3 (g3359), .I4 (g3341));
AN2X1 gate6850(.O (g9147), .I1 (g9136), .I2 (g6103));
AN2X1 gate6851(.O (g5062), .I1 (g235), .I2 (g3973));
AN2X1 gate6852(.O (g9347), .I1 (g9332), .I2 (g6226));
AN2X1 gate6853(.O (g4825), .I1 (g4228), .I2 (g1964));
AN2X1 gate6854(.O (g8721), .I1 (g2703), .I2 (g8464));
AN2X1 gate6855(.O (g7552), .I1 (g7319), .I2 (g5749));
AN2X1 gate6856(.O (g7606), .I1 (g7471), .I2 (g3466));
AN2X1 gate6857(.O (g4408), .I1 (g330), .I2 (g3131));
AN2X1 gate6858(.O (g9013), .I1 (g8907), .I2 (g8239));
AN2X1 gate6859(.O (g5298), .I1 (g1912), .I2 (g4814));
AN2X1 gate6860(.O (g6976), .I1 (g4399), .I2 (g6508));
AN2X1 gate6861(.O (g8940), .I1 (g4543), .I2 (g8775));
AN4X1 gate6862(.O (I8588), .I1 (g3430), .I2 (g3398), .I3 (g3359), .I4 (g3341));
AN3X1 gate6863(.O (g4230), .I1 (g2683), .I2 (g3491), .I3 (I8143));
AN2X1 gate6864(.O (g6400), .I1 (g150), .I2 (g6011));
AN3X1 gate6865(.O (I8127), .I1 (g2699), .I2 (g2674), .I3 (g2677));
AN2X1 gate6866(.O (g4433), .I1 (g278), .I2 (g3097));
AN2X1 gate6867(.O (g7691), .I1 (g7367), .I2 (g4427));
AN2X1 gate6868(.O (g5031), .I1 (g292), .I2 (g3948));
AN2X1 gate6869(.O (g7607), .I1 (g7325), .I2 (g4969));
AN2X1 gate6870(.O (g8826), .I1 (g420), .I2 (g8564));
AN2X1 gate6871(.O (g4395), .I1 (g405), .I2 (g3160));
AN2X1 gate6872(.O (g8741), .I1 (g3787), .I2 (g8464));
AN3X1 gate6873(.O (g5005), .I1 (g2728), .I2 (g4320), .I3 (I9330));
AN2X1 gate6874(.O (g2827), .I1 (g1889), .I2 (g1690));
AN2X1 gate6875(.O (g6423), .I1 (g5897), .I2 (g5384));
AN2X1 gate6876(.O (g5765), .I1 (g1695), .I2 (g5428));
AN4X1 gate6877(.O (I8240), .I1 (g2298), .I2 (g2316), .I3 (g2334), .I4 (g2354));
AN4X1 gate6878(.O (I8072), .I1 (g3316), .I2 (g3287), .I3 (g2020), .I4 (g3238));
AN2X1 gate6879(.O (g8609), .I1 (g7828), .I2 (g4969));
AN2X1 gate6880(.O (g8308), .I1 (g510), .I2 (g7966));
AN2X1 gate6881(.O (g7615), .I1 (g7488), .I2 (g3466));
AN2X1 gate6882(.O (g3229), .I1 (g1728), .I2 (g2015));
AN2X1 gate6883(.O (g8066), .I1 (g7488), .I2 (g7634));
AN4X1 gate6884(.O (I8034), .I1 (g2074), .I2 (g2057), .I3 (g3264), .I4 (g3238));
AN2X1 gate6885(.O (g4142), .I1 (I8005), .I2 (I8006));
AN2X1 gate6886(.O (g4342), .I1 (g228), .I2 (g3097));
AN3X1 gate6887(.O (I9222), .I1 (g4041), .I2 (g4044), .I3 (g2584));
AN2X1 gate6888(.O (g6999), .I1 (g815), .I2 (g6556));
AN4X1 gate6889(.O (g4255), .I1 (g3605), .I2 (g3644), .I3 (g3635), .I4 (I8186));
AN2X1 gate6890(.O (g6633), .I1 (g5526), .I2 (g5987));
AN2X1 gate6891(.O (g8711), .I1 (g3542), .I2 (g8407));
AN2X1 gate6892(.O (g5069), .I1 (g566), .I2 (g3983));
AN2X1 gate6893(.O (g4097), .I1 (g2624), .I2 (g2614));
AN2X1 gate6894(.O (g7832), .I1 (g5343), .I2 (g7599));
AN2X1 gate6895(.O (g4497), .I1 (I8551), .I2 (I8552));
AN2X1 gate6896(.O (g8455), .I1 (g652), .I2 (g7793));
AN2X1 gate6897(.O (g4154), .I1 (g1098), .I2 (g3495));
AN2X1 gate6898(.O (g8827), .I1 (g498), .I2 (g8585));
AN2X1 gate6899(.O (g8333), .I1 (g563), .I2 (g8181));
AN2X1 gate6900(.O (g6732), .I1 (g5874), .I2 (g5367));
AN2X1 gate6901(.O (g8846), .I1 (g510), .I2 (g8585));
AN2X1 gate6902(.O (g6753), .I1 (g5939), .I2 (g5384));
AN2X1 gate6903(.O (g7559), .I1 (g7367), .I2 (g4155));
AN4X1 gate6904(.O (I8413), .I1 (g3316), .I2 (g3287), .I3 (g3264), .I4 (g1987));
AN2X1 gate6905(.O (g5287), .I1 (g786), .I2 (g4724));
AN2X1 gate6906(.O (g4783), .I1 (g948), .I2 (g4527));
AN2X1 gate6907(.O (g6043), .I1 (g1069), .I2 (g5582));
AN4X1 gate6908(.O (g4312), .I1 (g3666), .I2 (g3684), .I3 (g3694), .I4 (g3707));
AN2X1 gate6909(.O (g7628), .I1 (g7367), .I2 (g4532));
AN2X1 gate6910(.O (g6434), .I1 (g855), .I2 (g6048));
AN2X1 gate6911(.O (g8290), .I1 (g588), .I2 (g8181));
AN2X1 gate6912(.O (g4129), .I1 (g2629), .I2 (g2621));
AN2X1 gate6913(.O (g8256), .I1 (g95), .I2 (g8131));
AN2X1 gate6914(.O (g4830), .I1 (g4288), .I2 (g3723));
AN2X1 gate6915(.O (g8816), .I1 (g336), .I2 (g8545));
AN2X1 gate6916(.O (g6914), .I1 (g6483), .I2 (g5246));
AN4X1 gate6917(.O (I8460), .I1 (g3430), .I2 (g3398), .I3 (g3359), .I4 (g2106));
AN2X1 gate6918(.O (g6013), .I1 (g5589), .I2 (g2424));
AN2X1 gate6919(.O (g6413), .I1 (g5939), .I2 (g5367));
AN2X1 gate6920(.O (g8700), .I1 (g3784), .I2 (g8342));
AN2X1 gate6921(.O (g7323), .I1 (g4065), .I2 (g7171));
AN2X1 gate6922(.O (g8263), .I1 (g4555), .I2 (g7905));
AN2X1 gate6923(.O (g8950), .I1 (g4582), .I2 (g8791));
AN2X1 gate6924(.O (g4068), .I1 (g121), .I2 (g3540));
AN4X1 gate6925(.O (I8079), .I1 (g3316), .I2 (g3287), .I3 (g2020), .I4 (g1987));
AN2X1 gate6926(.O (g5314), .I1 (g1509), .I2 (g4729));
AN2X1 gate6927(.O (g8723), .I1 (g2706), .I2 (g8421));
AN2X1 gate6928(.O (g8257), .I1 (g146), .I2 (g8042));
AN2X1 gate6929(.O (g8817), .I1 (g4545), .I2 (g8482));
AN2X1 gate6930(.O (g8301), .I1 (g182), .I2 (g8156));
AN2X1 gate6931(.O (g7010), .I1 (g1049), .I2 (g6574));
AN2X1 gate6932(.O (g6060), .I1 (g1065), .I2 (g5623));
AN2X1 gate6933(.O (g4699), .I1 (g1557), .I2 (g4276));
AN2X1 gate6934(.O (g6460), .I1 (g6178), .I2 (g2424));
AN2X1 gate6935(.O (g4398), .I1 (g567), .I2 (g2845));
AN2X1 gate6936(.O (g5008), .I1 (g231), .I2 (g3920));
AN2X1 gate6937(.O (g7278), .I1 (g6965), .I2 (g1745));
AN2X1 gate6938(.O (g6995), .I1 (g6435), .I2 (g1616));
AN2X1 gate6939(.O (g8441), .I1 (g746), .I2 (g8018));
AN2X1 gate6940(.O (g7235), .I1 (g6699), .I2 (g7094));
AN4X1 gate6941(.O (I8432), .I1 (g3316), .I2 (g3287), .I3 (g2020), .I4 (g3238));
AN2X1 gate6942(.O (g9084), .I1 (g8964), .I2 (g5345));
AN4X1 gate6943(.O (I8053), .I1 (g3316), .I2 (g3287), .I3 (g3264), .I4 (g3238));
AN2X1 gate6944(.O (g7282), .I1 (g5830), .I2 (g6939));
AN2X1 gate6945(.O (g5065), .I1 (g374), .I2 (g3977));
AN2X1 gate6946(.O (g5122), .I1 (g436), .I2 (g4030));
AN4X1 gate6947(.O (g4319), .I1 (g3728), .I2 (g3694), .I3 (g3750), .I4 (I8296));
AN2X1 gate6948(.O (g7693), .I1 (g7367), .I2 (g4445));
AN4X1 gate6949(.O (I8568), .I1 (g3430), .I2 (g3398), .I3 (g3359), .I4 (g3341));
AN2X1 gate6950(.O (g4352), .I1 (g387), .I2 (g3160));
AN2X1 gate6951(.O (g5033), .I1 (g393), .I2 (g3953));
AN3X1 gate6952(.O (I8157), .I1 (g2686), .I2 (g2689), .I3 (g2692));
AN2X1 gate6953(.O (g8458), .I1 (g756), .I2 (g8199));
AN2X1 gate6954(.O (g5096), .I1 (g1149), .I2 (g4400));
AN2X1 gate6955(.O (g4186), .I1 (g1118), .I2 (g3520));
AN2X1 gate6956(.O (g9276), .I1 (g9244), .I2 (g5649));
AN2X1 gate6957(.O (g4386), .I1 (g324), .I2 (g3131));
AN2X1 gate6958(.O (g6954), .I1 (g5518), .I2 (g6601));
AN2X1 gate6959(.O (g8074), .I1 (g855), .I2 (g7616));
AN2X1 gate6960(.O (g6053), .I1 (g1053), .I2 (g5608));
AN2X1 gate6961(.O (g4083), .I1 (g125), .I2 (g3610));
AN2X1 gate6962(.O (g8080), .I1 (g7467), .I2 (g7634));
AN2X1 gate6963(.O (g4483), .I1 (I8523), .I2 (I8524));
AN2X1 gate6964(.O (g3259), .I1 (g1976), .I2 (g1960));
AN2X1 gate6965(.O (g8713), .I1 (g2777), .I2 (g8421));
AN2X1 gate6966(.O (g5142), .I1 (g1677), .I2 (g4202));
AN2X1 gate6967(.O (g6157), .I1 (g1130), .I2 (g5717));
AN2X1 gate6968(.O (g5081), .I1 (g455), .I2 (g3993));
AN2X1 gate6969(.O (g9120), .I1 (g9052), .I2 (g5345));
AN2X1 gate6970(.O (g4187), .I1 (I8078), .I2 (I8079));
AN2X1 gate6971(.O (g9277), .I1 (g9248), .I2 (g5654));
AN2X1 gate6972(.O (g4387), .I1 (g378), .I2 (g3160));
AN2X1 gate6973(.O (g8688), .I1 (g3812), .I2 (g8342));
AN2X1 gate6974(.O (g8857), .I1 (g446), .I2 (g8564));
AN2X1 gate6975(.O (g8976), .I1 (g8903), .I2 (g6588));
AN2X1 gate6976(.O (g4427), .I1 (I8431), .I2 (I8432));
AN2X1 gate6977(.O (g4514), .I1 (I8588), .I2 (I8589));
AN2X1 gate6978(.O (g5783), .I1 (g1897), .I2 (g5287));
AN2X1 gate6979(.O (g7724), .I1 (g7337), .I2 (g5938));
AN2X1 gate6980(.O (g7179), .I1 (g6121), .I2 (g7035));
AN2X1 gate6981(.O (g4403), .I1 (I8400), .I2 (I8401));
AN2X1 gate6982(.O (g8326), .I1 (g258), .I2 (g7838));
AN2X1 gate6983(.O (g4145), .I1 (g2639), .I2 (g2635));
AN2X1 gate6984(.O (g4391), .I1 (g249), .I2 (g3097));
AN2X1 gate6985(.O (g5001), .I1 (g458), .I2 (g3912));
AN2X1 gate6986(.O (g7658), .I1 (g7367), .I2 (g4150));
AN2X1 gate6987(.O (g4107), .I1 (g2625), .I2 (g2615));
AN2X1 gate6988(.O (g1834), .I1 (g933), .I2 (g929));
AN2X1 gate6989(.O (g7271), .I1 (g6436), .I2 (g6922));
AN2X1 gate6990(.O (g4159), .I1 (g1102), .I2 (g3498));
AN2X1 gate6991(.O (g8383), .I1 (g730), .I2 (g7937));
AN2X1 gate6992(.O (g8924), .I1 (g4588), .I2 (g8752));
AN2X1 gate6993(.O (g7611), .I1 (g7367), .I2 (g4507));
AN2X1 gate6994(.O (g8779), .I1 (g8634), .I2 (g7037));
AN2X1 gate6995(.O (g6949), .I1 (g5483), .I2 (g6589));
AN3X1 gate6996(.O (g4315), .I1 (g3707), .I2 (g3728), .I3 (I8288));
AN2X1 gate6997(.O (g4047), .I1 (g1272), .I2 (g3503));
AN2X1 gate6998(.O (g8361), .I1 (g426), .I2 (g7920));
AN2X1 gate6999(.O (g6998), .I1 (g4474), .I2 (g6555));
AN2X1 gate7000(.O (g7238), .I1 (g6707), .I2 (g7098));
AN2X1 gate7001(.O (g5624), .I1 (g5140), .I2 (g2794));
AN2X1 gate7002(.O (g7680), .I1 (g7367), .I2 (g4166));
AN2X1 gate7003(.O (g8327), .I1 (g336), .I2 (g7870));
AN2X1 gate7004(.O (g6039), .I1 (g1037), .I2 (g5574));
AN2X1 gate7005(.O (g5068), .I1 (g475), .I2 (g3982));
AN2X1 gate7006(.O (g6439), .I1 (g789), .I2 (g6150));
AN4X1 gate7007(.O (I8546), .I1 (g3430), .I2 (g3398), .I3 (g3359), .I4 (g3341));
AN2X1 gate7008(.O (g8303), .I1 (g284), .I2 (g7838));
AN2X1 gate7009(.O (g8696), .I1 (g3743), .I2 (g8342));
AN2X1 gate7010(.O (g8732), .I1 (g3808), .I2 (g8464));
AN2X1 gate7011(.O (g4272), .I1 (g3233), .I2 (g3286));
AN2X1 gate7012(.O (g8944), .I1 (g4539), .I2 (g8783));
AN2X1 gate7013(.O (g5699), .I1 (g1667), .I2 (g4841));
AN2X1 gate7014(.O (g4417), .I1 (I8417), .I2 (I8418));
AN4X1 gate7015(.O (I8617), .I1 (g3430), .I2 (g3398), .I3 (g3359), .I4 (g2106));
AN2X1 gate7016(.O (g7600), .I1 (g7460), .I2 (g3466));
AN2X1 gate7017(.O (g4128), .I1 (g98), .I2 (g3693));
AN2X1 gate7018(.O (g3081), .I1 (g1682), .I2 (g1616));
AN2X1 gate7019(.O (g8316), .I1 (g513), .I2 (g7966));
AN4X1 gate7020(.O (I8299), .I1 (g3666), .I2 (g3684), .I3 (g3694), .I4 (g3707));
AN4X1 gate7021(.O (I8547), .I1 (g3316), .I2 (g2057), .I3 (g2020), .I4 (g3238));
AN2X1 gate7022(.O (g6970), .I1 (g5035), .I2 (g6490));
AN2X1 gate7023(.O (g8147), .I1 (g1065), .I2 (g7683));
AN2X1 gate7024(.O (g5119), .I1 (g543), .I2 (g4027));
AN2X1 gate7025(.O (g8697), .I1 (g3761), .I2 (g8342));
AN2X1 gate7026(.O (g8914), .I1 (g8795), .I2 (g8239));
AN4X1 gate7027(.O (g4902), .I1 (g4304), .I2 (g2770), .I3 (g2746), .I4 (g2728));
AN4X1 gate7028(.O (I8078), .I1 (g2162), .I2 (g2149), .I3 (g2137), .I4 (g2106));
AN2X1 gate7029(.O (g7175), .I1 (g6893), .I2 (g4841));
AN2X1 gate7030(.O (g5599), .I1 (g4745), .I2 (g4969));
AN2X1 gate7031(.O (g4490), .I1 (g521), .I2 (g3192));
AN3X1 gate7032(.O (g4823), .I1 (g4238), .I2 (g4230), .I3 (g174));
AN2X1 gate7033(.O (g4166), .I1 (I8045), .I2 (I8046));
AN2X1 gate7034(.O (g8820), .I1 (g261), .I2 (g8524));
AN2X1 gate7035(.O (g4366), .I1 (g216), .I2 (g3097));
AN2X1 gate7036(.O (g8936), .I1 (g3875), .I2 (g8768));
AN2X1 gate7037(.O (g6771), .I1 (g146), .I2 (g6004));
AN2X1 gate7038(.O (g8317), .I1 (g547), .I2 (g8181));
AN2X1 gate7039(.O (g4529), .I1 (I8612), .I2 (I8613));
AN2X1 gate7040(.O (g5125), .I1 (g517), .I2 (g4036));
AN2X1 gate7041(.O (g7184), .I1 (g6138), .I2 (g7043));
AN2X1 gate7042(.O (g4155), .I1 (I8028), .I2 (I8029));
AN2X1 gate7043(.O (g5984), .I1 (g1041), .I2 (g5484));
AN2X1 gate7044(.O (g4355), .I1 (g390), .I2 (g3160));
AN2X1 gate7045(.O (g8922), .I1 (g4586), .I2 (g8750));
AN2X1 gate7046(.O (g6738), .I1 (g5847), .I2 (g5367));
AN2X1 gate7047(.O (g8060), .I1 (g7535), .I2 (g4841));
AN2X1 gate7048(.O (g5106), .I1 (g398), .I2 (g4015));
AN2X1 gate7049(.O (g6991), .I1 (g5689), .I2 (g6520));
AN2X1 gate7050(.O (g8460), .I1 (g757), .I2 (g8199));
AN2X1 gate7051(.O (g9038), .I1 (g8966), .I2 (g5345));
AN2X1 gate7052(.O (g8739), .I1 (g3780), .I2 (g8464));
AN2X1 gate7053(.O (g4720), .I1 (g190), .I2 (g4055));
AN2X1 gate7054(.O (g4118), .I1 (g995), .I2 (g3790));
AN2X1 gate7055(.O (g4167), .I1 (g2783), .I2 (g1616));
AN2X1 gate7056(.O (g4367), .I1 (g240), .I2 (g3097));
AN3X1 gate7057(.O (g4872), .I1 (g1924), .I2 (g4225), .I3 (g4224));
AN2X1 gate7058(.O (g7634), .I1 (g7367), .I2 (g4549));
AN2X1 gate7059(.O (g8937), .I1 (g4524), .I2 (g8770));
AN2X1 gate7060(.O (g8079), .I1 (g831), .I2 (g7658));
AN2X1 gate7061(.O (g8294), .I1 (g281), .I2 (g7838));
AN2X1 gate7062(.O (g5046), .I1 (g314), .I2 (g3962));
AN2X1 gate7063(.O (g8840), .I1 (g4590), .I2 (g8582));
AN2X1 gate7064(.O (g4193), .I1 (g145), .I2 (g2727));
AN2X1 gate7065(.O (g4393), .I1 (g327), .I2 (g3131));
AN2X1 gate7066(.O (g4549), .I1 (I8642), .I2 (I8643));
AN2X1 gate7067(.O (g6915), .I1 (g6493), .I2 (g5246));
AN4X1 gate7068(.O (I8064), .I1 (g3316), .I2 (g3287), .I3 (g3264), .I4 (g1987));
AN2X1 gate7069(.O (g8942), .I1 (g4522), .I2 (g8780));
AN2X1 gate7070(.O (g2912), .I1 (g1080), .I2 (g1945));
AN2X1 gate7071(.O (g5107), .I1 (g478), .I2 (g4016));
AN2X1 gate7072(.O (g8704), .I1 (g2829), .I2 (g8386));
AN2X1 gate7073(.O (g6002), .I1 (g5539), .I2 (g2407));
AN2X1 gate7074(.O (g6402), .I1 (g665), .I2 (g6012));
AN2X1 gate7075(.O (g8954), .I1 (g8763), .I2 (g6097));
AN3X1 gate7076(.O (I8237), .I1 (g2298), .I2 (g2316), .I3 (g2354));
AN2X1 gate7077(.O (g6762), .I1 (g5847), .I2 (g5412));
AN2X1 gate7078(.O (g4740), .I1 (g2242), .I2 (g4275));
AN4X1 gate7079(.O (g3258), .I1 (g2298), .I2 (g2316), .I3 (g2334), .I4 (g2354));
AN2X1 gate7080(.O (g5047), .I1 (g373), .I2 (g3964));
AN4X1 gate7081(.O (I8089), .I1 (g2162), .I2 (g2149), .I3 (g2137), .I4 (g2106));
AN2X1 gate7082(.O (g8912), .I1 (g8796), .I2 (g8239));
AN4X1 gate7083(.O (I8071), .I1 (g2162), .I2 (g2149), .I3 (g2137), .I4 (g2106));
AN2X1 gate7084(.O (g6464), .I1 (g6177), .I2 (g2424));
AN2X1 gate7085(.O (g8929), .I1 (g3865), .I2 (g8759));
AN2X1 gate7086(.O (g3614), .I1 (g1134), .I2 (g2386));
AN2X1 gate7087(.O (g7036), .I1 (g6728), .I2 (g5197));
AN2X1 gate7088(.O (g7679), .I1 (g7447), .I2 (g5084));
AN2X1 gate7089(.O (g8626), .I1 (g752), .I2 (g8199));
AN2X1 gate7090(.O (g3984), .I1 (g2403), .I2 (g3085));
AN2X1 gate7091(.O (g5017), .I1 (g211), .I2 (g3928));
AN2X1 gate7092(.O (g4691), .I1 (g4219), .I2 (g1690));
AN2X1 gate7093(.O (g2949), .I1 (g822), .I2 (g1753));
AN2X1 gate7094(.O (g7182), .I1 (g6902), .I2 (g4969));
AN2X1 gate7095(.O (g6394), .I1 (g5988), .I2 (g5494));
AN2X1 gate7096(.O (g4962), .I1 (g457), .I2 (g3905));
AN2X1 gate7097(.O (g4158), .I1 (I8033), .I2 (I8034));
AN2X1 gate7098(.O (g6966), .I1 (g6580), .I2 (g5580));
AN2X1 gate7099(.O (g8735), .I1 (g2807), .I2 (g8443));
AN2X1 gate7100(.O (g8075), .I1 (g7460), .I2 (g7634));
AN2X1 gate7101(.O (g8949), .I1 (g4572), .I2 (g8790));
AN2X1 gate7102(.O (g7632), .I1 (g7445), .I2 (g3548));
AN2X1 gate7103(.O (g7653), .I1 (g7480), .I2 (g5754));
AN2X1 gate7104(.O (g8292), .I1 (g181), .I2 (g8156));
AN2X1 gate7105(.O (g2952), .I1 (g2474), .I2 (g2215));
AN2X1 gate7106(.O (g6438), .I1 (g4829), .I2 (g6051));
AN2X1 gate7107(.O (g4284), .I1 (g3260), .I2 (g3314));
AN2X1 gate7108(.O (g4239), .I1 (g1541), .I2 (g3222));
AN2X1 gate7109(.O (g5090), .I1 (g317), .I2 (g4000));
AN2X1 gate7110(.O (g8646), .I1 (g553), .I2 (g8094));
AN2X1 gate7111(.O (g6409), .I1 (g706), .I2 (g6020));
AN2X1 gate7112(.O (g4180), .I1 (g1114), .I2 (g3511));
AN2X1 gate7113(.O (g9270), .I1 (g4748), .I2 (g9241));
AN2X1 gate7114(.O (g4380), .I1 (g584), .I2 (g2845));
AN2X1 gate7115(.O (g4832), .I1 (g1110), .I2 (g4246));
AN2X1 gate7116(.O (g8439), .I1 (g699), .I2 (g7811));
AN2X1 gate7117(.O (g2986), .I1 (g806), .I2 (g1739));
AN2X1 gate7118(.O (g4420), .I1 (g275), .I2 (g3097));
AN2X1 gate7119(.O (g4507), .I1 (I8573), .I2 (I8574));
AN2X1 gate7120(.O (g4794), .I1 (g954), .I2 (g4574));
AN2X1 gate7121(.O (g8702), .I1 (g2837), .I2 (g8386));
AN2X1 gate7122(.O (g8919), .I1 (g4567), .I2 (g8743));
AN2X1 gate7123(.O (g8952), .I1 (g8788), .I2 (g6075));
AN2X1 gate7124(.O (g8276), .I1 (g150), .I2 (g8042));
AN2X1 gate7125(.O (g5063), .I1 (g294), .I2 (g3974));
AN2X1 gate7126(.O (g4100), .I1 (g113), .I2 (g3648));
AN2X1 gate7127(.O (g7553), .I1 (g7367), .I2 (g4135));
AN2X1 gate7128(.O (g8404), .I1 (g710), .I2 (g7937));
AN2X1 gate7129(.O (g5118), .I1 (g479), .I2 (g4026));
AN2X1 gate7130(.O (g8764), .I1 (g8231), .I2 (g4969));
OR4X1 gate7131(.O (g5057), .I1 (g3939), .I2 (g3925), .I3 (g3915), .I4 (g3907));
OR4X1 gate7132(.O (I14941), .I1 (g8275), .I2 (g8323), .I3 (g8459), .I4 (g8380));
OR2X1 gate7133(.O (g5193), .I1 (g5017), .I2 (g4366));
OR2X1 gate7134(.O (g9291), .I1 (g9273), .I2 (g6216));
OR2X1 gate7135(.O (g5549), .I1 (g2935), .I2 (g4712));
OR2X1 gate7136(.O (g7029), .I1 (g6433), .I2 (g5765));
OR2X1 gate7137(.O (g7787), .I1 (g4791), .I2 (g7602));
OR2X1 gate7138(.O (g6249), .I1 (g4066), .I2 (g5313));
OR3X1 gate7139(.O (g8906), .I1 (g8088), .I2 (g8062), .I3 (g8699));
OR2X1 gate7140(.O (g5232), .I1 (g5082), .I2 (g4412));
OR2X1 gate7141(.O (g8987), .I1 (g8927), .I2 (g8826));
OR2X1 gate7142(.O (g5253), .I1 (g5116), .I2 (g4451));
OR2X1 gate7143(.O (g7791), .I1 (g4796), .I2 (g7606));
OR4X1 gate7144(.O (I8225), .I1 (g3062), .I2 (g2712), .I3 (g2734), .I4 (g2752));
OR4X1 gate7145(.O (I15250), .I1 (g8238), .I2 (g8265), .I3 (g8272), .I4 (g8292));
OR2X1 gate7146(.O (g8991), .I1 (g8931), .I2 (g8831));
OR4X1 gate7147(.O (I9107), .I1 (g4133), .I2 (g4145), .I3 (g4138), .I4 (g4132));
OR2X1 gate7148(.O (g9008), .I1 (g8948), .I2 (g8857));
OR4X1 gate7149(.O (g2214), .I1 (g1376), .I2 (g1377), .I3 (g1378), .I4 (g1379));
OR2X1 gate7150(.O (g7575), .I1 (g7323), .I2 (g7142));
OR2X1 gate7151(.O (g9136), .I1 (g8952), .I2 (g9131));
OR3X1 gate7152(.O (g8907), .I1 (g8081), .I2 (g8064), .I3 (g8707));
OR3X1 gate7153(.O (g8082), .I1 (g7654), .I2 (g7628), .I3 (g7611));
OR2X1 gate7154(.O (g5710), .I1 (g4958), .I2 (g4351));
OR3X1 gate7155(.O (I9047), .I1 (g4155), .I2 (g4147), .I3 (g4139));
OR2X1 gate7156(.O (g9122), .I1 (g8953), .I2 (g9084));
OR3X1 gate7157(.O (g6270), .I1 (g1000), .I2 (g5335), .I3 (g1909));
OR2X1 gate7158(.O (g6610), .I1 (g4180), .I2 (g6061));
OR2X1 gate7159(.O (g6124), .I1 (g5432), .I2 (g4789));
OR2X1 gate7160(.O (g6980), .I1 (g6745), .I2 (g6028));
OR4X1 gate7161(.O (I14484), .I1 (g7993), .I2 (g7966), .I3 (g7793), .I4 (g7811));
OR2X1 gate7162(.O (g9137), .I1 (g8877), .I2 (g9118));
OR2X1 gate7163(.O (g9337), .I1 (g9240), .I2 (g9327));
OR2X1 gate7164(.O (g7086), .I1 (g4101), .I2 (g6464));
OR4X1 gate7165(.O (I15055), .I1 (I15051), .I2 (I15052), .I3 (I15053), .I4 (I15054));
OR4X1 gate7166(.O (I15111), .I1 (g7951), .I2 (g7920), .I3 (g7983), .I4 (g8181));
OR2X1 gate7167(.O (g5545), .I1 (g3617), .I2 (g4824));
OR2X1 gate7168(.O (g7025), .I1 (g6541), .I2 (g3095));
OR2X1 gate7169(.O (g4264), .I1 (g2490), .I2 (g3315));
OR2X1 gate7170(.O (g8899), .I1 (g8839), .I2 (g8652));
OR3X1 gate7171(.O (g8785), .I1 (g8623), .I2 (g8656), .I3 (I14985));
OR4X1 gate7172(.O (I15019), .I1 (g7951), .I2 (g7920), .I3 (g7983), .I4 (g8181));
OR2X1 gate7173(.O (g6144), .I1 (g4175), .I2 (g5458));
OR2X1 gate7174(.O (g9154), .I1 (g9142), .I2 (g9021));
OR2X1 gate7175(.O (g9354), .I1 (g9275), .I2 (g9344));
OR4X1 gate7176(.O (I15018), .I1 (g7855), .I2 (g7838), .I3 (g7905), .I4 (g7870));
OR2X1 gate7177(.O (g4179), .I1 (g207), .I2 (g3083));
OR2X1 gate7178(.O (g7682), .I1 (g6044), .I2 (g7412));
OR2X1 gate7179(.O (g6694), .I1 (g6151), .I2 (g5573));
OR2X1 gate7180(.O (g5204), .I1 (g5033), .I2 (g4379));
OR2X1 gate7181(.O (g9267), .I1 (g9251), .I2 (g6225));
OR2X1 gate7182(.O (g9001), .I1 (g8941), .I2 (g8846));
OR4X1 gate7183(.O (g8966), .I1 (g8741), .I2 (g8745), .I3 (g8912), .I4 (g8850));
OR2X1 gate7184(.O (g7445), .I1 (g4192), .I2 (g7193));
OR4X1 gate7185(.O (g5040), .I1 (g3900), .I2 (g3895), .I3 (g3890), .I4 (g4363));
OR2X1 gate7186(.O (g5440), .I1 (g4790), .I2 (g4786));
OR4X1 gate7187(.O (I15102), .I1 (I15098), .I2 (I15099), .I3 (I15100), .I4 (I15101));
OR4X1 gate7188(.O (g2229), .I1 (g1371), .I2 (g1372), .I3 (g1373), .I4 (g1374));
OR4X1 gate7189(.O (I14771), .I1 (g7993), .I2 (g7966), .I3 (g7793), .I4 (g7811));
OR4X1 gate7190(.O (I15231), .I1 (g8701), .I2 (g8715), .I3 (g8730), .I4 (g8720));
OR2X1 gate7191(.O (g8773), .I1 (I14959), .I2 (I14960));
OR4X1 gate7192(.O (g8009), .I1 (g3591), .I2 (g7406), .I3 (g7566), .I4 (I14302));
OR2X1 gate7193(.O (g8769), .I1 (I14951), .I2 (I14952));
OR2X1 gate7194(.O (g7227), .I1 (g6992), .I2 (g3128));
OR2X1 gate7195(.O (g6934), .I1 (g6422), .I2 (g6430));
OR2X1 gate7196(.O (g8993), .I1 (g8933), .I2 (g8835));
OR2X1 gate7197(.O (g6913), .I1 (g6733), .I2 (g6738));
OR2X1 gate7198(.O (g5235), .I1 (g5091), .I2 (g4422));
OR2X1 gate7199(.O (g5343), .I1 (g4690), .I2 (g2862));
OR4X1 gate7200(.O (I15085), .I1 (g8363), .I2 (g8342), .I3 (g8407), .I4 (g8386));
OR2X1 gate7201(.O (g5566), .I1 (g3617), .I2 (g4810));
OR4X1 gate7202(.O (I14759), .I1 (g7937), .I2 (g7887), .I3 (g8029), .I4 (g8018));
OR4X1 gate7203(.O (I15054), .I1 (g8363), .I2 (g8342), .I3 (g8407), .I4 (g8386));
OR4X1 gate7204(.O (I15243), .I1 (I15239), .I2 (I15240), .I3 (I15241), .I4 (I15242));
OR4X1 gate7205(.O (I14758), .I1 (g7993), .I2 (g7966), .I3 (g7793), .I4 (g7811));
OR3X1 gate7206(.O (g4736), .I1 (g4532), .I2 (g4517), .I3 (I9044));
OR2X1 gate7207(.O (g8895), .I1 (g8823), .I2 (g8646));
OR2X1 gate7208(.O (g7428), .I1 (g6040), .I2 (g7175));
OR2X1 gate7209(.O (g9352), .I1 (g9343), .I2 (g4526));
OR2X1 gate7210(.O (g7826), .I1 (g4804), .I2 (g7626));
OR3X1 gate7211(.O (g8788), .I1 (g8620), .I2 (g8658), .I3 (I14990));
OR2X1 gate7212(.O (g5202), .I1 (g5031), .I2 (g4377));
OR2X1 gate7213(.O (g5518), .I1 (g4744), .I2 (g4118));
OR4X1 gate7214(.O (g4737), .I1 (g4135), .I2 (g4529), .I3 (g4514), .I4 (I9047));
OR2X1 gate7215(.O (g7165), .I1 (g6434), .I2 (g6908));
OR2X1 gate7216(.O (g5264), .I1 (g5125), .I2 (g4490));
OR4X1 gate7217(.O (g8176), .I1 (g7566), .I2 (g1030), .I3 (g6664), .I4 (g6452));
OR2X1 gate7218(.O (g9387), .I1 (g9349), .I2 (g9384));
OR4X1 gate7219(.O (g2206), .I1 (g1363), .I2 (g1364), .I3 (g1365), .I4 (g1366));
OR4X1 gate7220(.O (I14951), .I1 (g8328), .I2 (g8316), .I3 (g8455), .I4 (g8378));
OR4X1 gate7221(.O (g9046), .I1 (g8744), .I2 (g8749), .I3 (g9016), .I4 (g8862));
OR2X1 gate7222(.O (g6932), .I1 (g6417), .I2 (g6423));
OR3X1 gate7223(.O (I15169), .I1 (g8483), .I2 (g8464), .I3 (g8514));
OR2X1 gate7224(.O (g9003), .I1 (g8943), .I2 (g8849));
OR4X1 gate7225(.O (g8796), .I1 (g8150), .I2 (g8078), .I3 (g8070), .I4 (g8360));
OR2X1 gate7226(.O (g8980), .I1 (g8920), .I2 (g8815));
OR2X1 gate7227(.O (g6716), .I1 (g6162), .I2 (g5588));
OR2X1 gate7228(.O (g7421), .I1 (g6745), .I2 (g7202));
OR2X1 gate7229(.O (g6699), .I1 (g6154), .I2 (g5579));
OR2X1 gate7230(.O (g5238), .I1 (g5094), .I2 (g4425));
OR2X1 gate7231(.O (g4927), .I1 (g4318), .I2 (g1590));
OR2X1 gate7232(.O (g5209), .I1 (g5044), .I2 (g4384));
OR4X1 gate7233(.O (I15084), .I1 (g7951), .I2 (g7920), .I3 (g7983), .I4 (g8181));
OR4X1 gate7234(.O (I15110), .I1 (g7855), .I2 (g7838), .I3 (g7905), .I4 (g7870));
OR2X1 gate7235(.O (g8900), .I1 (g8840), .I2 (g8653));
OR2X1 gate7236(.O (g5511), .I1 (g4743), .I2 (g4109));
OR2X1 gate7237(.O (g6717), .I1 (g4082), .I2 (g6005));
OR2X1 gate7238(.O (g3160), .I1 (g1751), .I2 (g449));
OR3X1 gate7239(.O (g8886), .I1 (g8727), .I2 (g8812), .I3 (I15254));
OR4X1 gate7240(.O (g2230), .I1 (g1380), .I2 (g1381), .I3 (g1382), .I4 (g1383));
OR4X1 gate7241(.O (I15242), .I1 (g8697), .I2 (g8714), .I3 (g8718), .I4 (g8719));
OR2X1 gate7242(.O (g5722), .I1 (g5001), .I2 (g4361));
OR2X1 gate7243(.O (g2845), .I1 (g1877), .I2 (g576));
OR4X1 gate7244(.O (I15230), .I1 (g8274), .I2 (g8321), .I3 (g8298), .I4 (g8696));
OR4X1 gate7245(.O (I15265), .I1 (I15261), .I2 (I15262), .I3 (I15263), .I4 (I15264));
OR4X1 gate7246(.O (g4786), .I1 (g4107), .I2 (g4097), .I3 (g4124), .I4 (I9099));
OR3X1 gate7247(.O (I13553), .I1 (g1166), .I2 (g1167), .I3 (g1170));
OR2X1 gate7248(.O (g8887), .I1 (I15265), .I2 (g8819));
OR2X1 gate7249(.O (g7080), .I1 (g4086), .I2 (g6462));
OR2X1 gate7250(.O (g4364), .I1 (g2952), .I2 (g1725));
OR2X1 gate7251(.O (g9148), .I1 (g9143), .I2 (g9024));
OR4X1 gate7252(.O (I14767), .I1 (g7937), .I2 (g7887), .I3 (g8029), .I4 (g8018));
OR2X1 gate7253(.O (g9355), .I1 (g9276), .I2 (g9345));
OR2X1 gate7254(.O (g3541), .I1 (g1663), .I2 (g1421));
OR3X1 gate7255(.O (I14990), .I1 (g8337), .I2 (g8379), .I3 (g8543));
OR2X1 gate7256(.O (g5231), .I1 (g5081), .I2 (g4411));
OR2X1 gate7257(.O (g5205), .I1 (g5034), .I2 (g4380));
OR4X1 gate7258(.O (g8891), .I1 (g8705), .I2 (g8811), .I3 (I15297), .I4 (I15298));
OR4X1 gate7259(.O (I15041), .I1 (g7855), .I2 (g7838), .I3 (g7905), .I4 (g7870));
OR2X1 gate7260(.O (g6115), .I1 (g3617), .I2 (g5558));
OR4X1 gate7261(.O (I15275), .I1 (g8693), .I2 (g8703), .I3 (g8712), .I4 (g8717));
OR2X1 gate7262(.O (g4297), .I1 (g3617), .I2 (g3602));
OR2X1 gate7263(.O (g7220), .I1 (g1304), .I2 (g7062));
OR2X1 gate7264(.O (g5572), .I1 (g5051), .I2 (g1236));
OR2X1 gate7265(.O (g8154), .I1 (g6054), .I2 (g7607));
OR4X1 gate7266(.O (I14766), .I1 (g7993), .I2 (g7966), .I3 (g7793), .I4 (g7811));
OR2X1 gate7267(.O (g6935), .I1 (g6429), .I2 (g6431));
OR3X1 gate7268(.O (I15165), .I1 (g8483), .I2 (g8464), .I3 (g8514));
OR2X1 gate7269(.O (g8979), .I1 (g8919), .I2 (g8813));
OR2X1 gate7270(.O (g5036), .I1 (g4047), .I2 (g2972));
OR2X1 gate7271(.O (g3339), .I1 (g1424), .I2 (g2014));
OR4X1 gate7272(.O (I15253), .I1 (g8698), .I2 (g8711), .I3 (g8722), .I4 (g8716));
OR2X1 gate7273(.O (g7443), .I1 (g7192), .I2 (g3158));
OR4X1 gate7274(.O (I14754), .I1 (g7937), .I2 (g7887), .I3 (g8029), .I4 (g8018));
OR3X1 gate7275(.O (I15175), .I1 (g8483), .I2 (g8464), .I3 (g8514));
OR4X1 gate7276(.O (I15264), .I1 (g8700), .I2 (g8708), .I3 (g8726), .I4 (g8731));
OR2X1 gate7277(.O (g9358), .I1 (g9279), .I2 (g9348));
OR2X1 gate7278(.O (g7697), .I1 (g7419), .I2 (g3187));
OR2X1 gate7279(.O (g6698), .I1 (g4073), .I2 (g6001));
OR2X1 gate7280(.O (g6964), .I1 (g6447), .I2 (g6448));
OR2X1 gate7281(.O (g5208), .I1 (g5043), .I2 (g4383));
OR2X1 gate7282(.O (g9174), .I1 (g9147), .I2 (g8963));
OR4X1 gate7283(.O (I15021), .I1 (I15017), .I2 (I15018), .I3 (I15019), .I4 (I15020));
OR2X1 gate7284(.O (g9239), .I1 (g7653), .I2 (g9226));
OR2X1 gate7285(.O (g5265), .I1 (g5126), .I2 (g4491));
OR4X1 gate7286(.O (I15073), .I1 (g7951), .I2 (g7920), .I3 (g7983), .I4 (g8181));
OR4X1 gate7287(.O (I15274), .I1 (g8306), .I2 (g8361), .I3 (g8299), .I4 (g8687));
OR3X1 gate7288(.O (g6457), .I1 (g6196), .I2 (g6209), .I3 (g4937));
OR2X1 gate7289(.O (g5233), .I1 (g5089), .I2 (g4420));
OR2X1 gate7290(.O (g6686), .I1 (g4068), .I2 (g5970));
OR3X1 gate7291(.O (I15292), .I1 (g8704), .I2 (g8710), .I3 (g8805));
OR2X1 gate7292(.O (g8893), .I1 (g8814), .I2 (g8643));
OR4X1 gate7293(.O (g7784), .I1 (g7406), .I2 (g6664), .I3 (g3492), .I4 (I14219));
OR2X1 gate7294(.O (g6121), .I1 (g5425), .I2 (g4785));
OR3X1 gate7295(.O (I14366), .I1 (g7566), .I2 (g1030), .I3 (g6664));
OR2X1 gate7296(.O (g5706), .I1 (g4955), .I2 (g4342));
OR2X1 gate7297(.O (g6740), .I1 (g4100), .I2 (g6022));
OR2X1 gate7298(.O (g4283), .I1 (g3587), .I2 (g2665));
OR2X1 gate7299(.O (g8984), .I1 (g8924), .I2 (g8822));
OR4X1 gate7300(.O (I15109), .I1 (g8131), .I2 (g8111), .I3 (g8042), .I4 (g8156));
OR2X1 gate7301(.O (g9123), .I1 (g8954), .I2 (g9037));
OR4X1 gate7302(.O (I15283), .I1 (g8291), .I2 (g8276), .I3 (g8325), .I4 (g8330));
OR2X1 gate7303(.O (g5138), .I1 (g4108), .I2 (g3049));
OR2X1 gate7304(.O (g7810), .I1 (g4799), .I2 (g7609));
OR2X1 gate7305(.O (g7363), .I1 (g7136), .I2 (g6903));
OR3X1 gate7306(.O (I9099), .I1 (g4127), .I2 (g4123), .I3 (g4117));
OR2X1 gate7307(.O (g9151), .I1 (g9144), .I2 (g8961));
OR2X1 gate7308(.O (g6525), .I1 (g6112), .I2 (g5547));
OR2X1 gate7309(.O (g6710), .I1 (g55), .I2 (g6264));
OR4X1 gate7310(.O (I6209), .I1 (g911), .I2 (g916), .I3 (g921), .I4 (g883));
OR3X1 gate7311(.O (g8904), .I1 (g8090), .I2 (g8080), .I3 (g8706));
OR2X1 gate7312(.O (g5707), .I1 (g4956), .I2 (g4343));
OR3X1 gate7313(.O (I14980), .I1 (g8362), .I2 (g8403), .I3 (g8610));
OR2X1 gate7314(.O (g9010), .I1 (g8950), .I2 (g8860));
OR2X1 gate7315(.O (g5201), .I1 (g5030), .I2 (g4376));
OR3X1 gate7316(.O (g8763), .I1 (g8232), .I2 (I14941), .I3 (I14942));
OR3X1 gate7317(.O (I9044), .I1 (g4150), .I2 (g4142), .I3 (g4549));
OR2X1 gate7318(.O (g8637), .I1 (g6057), .I2 (g8071));
OR2X1 gate7319(.O (g5715), .I1 (g4961), .I2 (g4355));
OR2X1 gate7320(.O (g9282), .I1 (g9270), .I2 (g6238));
OR4X1 gate7321(.O (I15040), .I1 (g8131), .I2 (g8111), .I3 (g8042), .I4 (g8156));
OR2X1 gate7322(.O (g5052), .I1 (g4049), .I2 (g4054));
OR4X1 gate7323(.O (I15252), .I1 (g8320), .I2 (g8307), .I3 (g8317), .I4 (g8692));
OR2X1 gate7324(.O (g7782), .I1 (g4783), .I2 (g7598));
OR2X1 gate7325(.O (g6931), .I1 (g6416), .I2 (g6421));
OR4X1 gate7326(.O (I14969), .I1 (g8315), .I2 (g8377), .I3 (g8359), .I4 (g8611));
OR2X1 gate7327(.O (g5070), .I1 (g4052), .I2 (g4058));
OR4X1 gate7328(.O (g2213), .I1 (g1367), .I2 (g1368), .I3 (g1369), .I4 (g1370));
OR2X1 gate7329(.O (g8982), .I1 (g8922), .I2 (g8820));
OR2X1 gate7330(.O (g4055), .I1 (g187), .I2 (g3012));
OR3X1 gate7331(.O (g8128), .I1 (g7566), .I2 (g6910), .I3 (g6452));
OR3X1 gate7332(.O (I11603), .I1 (g6193), .I2 (g6197), .I3 (g6175));
OR2X1 gate7333(.O (g9264), .I1 (g9247), .I2 (g6242));
OR2X1 gate7334(.O (g6440), .I1 (g6268), .I2 (g5700));
OR2X1 gate7335(.O (g6123), .I1 (g3617), .I2 (g5556));
OR4X1 gate7336(.O (I15051), .I1 (g8131), .I2 (g8111), .I3 (g8042), .I4 (g8156));
OR4X1 gate7337(.O (I15072), .I1 (g7855), .I2 (g7838), .I3 (g7905), .I4 (g7870));
OR4X1 gate7338(.O (I14496), .I1 (g7937), .I2 (g7887), .I3 (g8029), .I4 (g8018));
OR2X1 gate7339(.O (g8902), .I1 (g8844), .I2 (g8654));
OR3X1 gate7340(.O (I15152), .I1 (g8483), .I2 (g8464), .I3 (g8514));
OR2X1 gate7341(.O (g8155), .I1 (g7632), .I2 (g3219));
OR3X1 gate7342(.O (g8964), .I1 (g8915), .I2 (g8863), .I3 (I15400));
OR2X1 gate7343(.O (g5227), .I1 (g5077), .I2 (g4407));
OR4X1 gate7344(.O (I15020), .I1 (g8363), .I2 (g8342), .I3 (g8407), .I4 (g8386));
OR2X1 gate7345(.O (g5203), .I1 (g5032), .I2 (g4378));
OR3X1 gate7346(.O (I9029), .I1 (g4504), .I2 (g4494), .I3 (g4430));
OR2X1 gate7347(.O (g8989), .I1 (g8929), .I2 (g8829));
OR4X1 gate7348(.O (I15113), .I1 (I15109), .I2 (I15110), .I3 (I15111), .I4 (I15112));
OR2X1 gate7349(.O (g8834), .I1 (g7096), .I2 (g8229));
OR2X1 gate7350(.O (g5188), .I1 (g5008), .I2 (g4365));
OR2X1 gate7351(.O (g7435), .I1 (g6052), .I2 (g7182));
OR2X1 gate7352(.O (g7690), .I1 (g4181), .I2 (g7417));
OR2X1 gate7353(.O (g5216), .I1 (g5062), .I2 (g4391));
OR2X1 gate7354(.O (g3131), .I1 (g1749), .I2 (g368));
OR2X1 gate7355(.O (g8909), .I1 (g6043), .I2 (g8764));
OR3X1 gate7356(.O (g4734), .I1 (g4469), .I2 (g4448), .I3 (I9038));
OR2X1 gate7357(.O (g6933), .I1 (g6419), .I2 (g6428));
OR4X1 gate7358(.O (I14480), .I1 (g7937), .I2 (g7887), .I3 (g8029), .I4 (g8018));
OR2X1 gate7359(.O (g9285), .I1 (g9271), .I2 (g6221));
OR4X1 gate7360(.O (I6208), .I1 (g891), .I2 (g896), .I3 (g901), .I4 (g906));
OR2X1 gate7361(.O (g5217), .I1 (g5063), .I2 (g4392));
OR2X1 gate7362(.O (g9139), .I1 (g8879), .I2 (g9120));
OR2X1 gate7363(.O (g9339), .I1 (g9259), .I2 (g9335));
OR2X1 gate7364(.O (g5711), .I1 (g4959), .I2 (g4352));
OR2X1 gate7365(.O (g7222), .I1 (g6049), .I2 (g6971));
OR4X1 gate7366(.O (I14942), .I1 (g8439), .I2 (g8440), .I3 (g8405), .I4 (g8460));
OR2X1 gate7367(.O (g4688), .I1 (g4193), .I2 (g3190));
OR2X1 gate7368(.O (g5196), .I1 (g5020), .I2 (g4369));
OR2X1 gate7369(.O (g6132), .I1 (g5436), .I2 (g4793));
OR2X1 gate7370(.O (g8985), .I1 (g8925), .I2 (g8824));
OR2X1 gate7371(.O (g7089), .I1 (g4128), .I2 (g6474));
OR2X1 gate7372(.O (g5256), .I1 (g5119), .I2 (g4454));
OR4X1 gate7373(.O (I14468), .I1 (g7937), .I2 (g7887), .I3 (g8029), .I4 (g8018));
OR4X1 gate7374(.O (g8794), .I1 (g8153), .I2 (g8074), .I3 (g8069), .I4 (g8523));
OR2X1 gate7375(.O (g5021), .I1 (g943), .I2 (g4501));
OR2X1 gate7376(.O (g7254), .I1 (g6923), .I2 (g5298));
OR2X1 gate7377(.O (g6600), .I1 (g5443), .I2 (g6055));
OR3X1 gate7378(.O (g8905), .I1 (g8089), .I2 (g8087), .I3 (g8694));
OR2X1 gate7379(.O (g7438), .I1 (g7184), .I2 (g6978));
OR2X1 gate7380(.O (g6580), .I1 (g6039), .I2 (g6041));
OR2X1 gate7381(.O (g6262), .I1 (g4074), .I2 (g5334));
OR4X1 gate7382(.O (I15229), .I1 (g8262), .I2 (g8303), .I3 (g8268), .I4 (g8312));
OR4X1 gate7383(.O (I14479), .I1 (g7993), .I2 (g7966), .I3 (g7793), .I4 (g7811));
OR4X1 gate7384(.O (I15228), .I1 (g8270), .I2 (g8258), .I3 (g8281), .I4 (g8273));
OR2X1 gate7385(.O (g4072), .I1 (g196), .I2 (g2995));
OR2X1 gate7386(.O (g9135), .I1 (g8951), .I2 (g9130));
OR2X1 gate7387(.O (g9288), .I1 (g9272), .I2 (g6235));
OR4X1 gate7388(.O (I15112), .I1 (g8363), .I2 (g8342), .I3 (g8407), .I4 (g8386));
OR2X1 gate7389(.O (g5673), .I1 (g4823), .I2 (g4872));
OR2X1 gate7390(.O (g7062), .I1 (g4048), .I2 (g6456));
OR2X1 gate7391(.O (g4413), .I1 (g2371), .I2 (g3285));
OR3X1 gate7392(.O (g8884), .I1 (g8735), .I2 (g8818), .I3 (I15232));
OR2X1 gate7393(.O (g7788), .I1 (g4794), .I2 (g7604));
OR2X1 gate7394(.O (g8988), .I1 (g8928), .I2 (g8827));
OR2X1 gate7395(.O (g6926), .I1 (g6406), .I2 (g6411));
OR2X1 gate7396(.O (g8804), .I1 (g6060), .I2 (g8609));
OR4X1 gate7397(.O (g9054), .I1 (g8724), .I2 (g8729), .I3 (g9013), .I4 (g8680));
OR4X1 gate7398(.O (I15298), .I1 (g8332), .I2 (g8333), .I3 (g8686), .I4 (g8702));
OR2X1 gate7399(.O (g6543), .I1 (g6125), .I2 (g1553));
OR3X1 gate7400(.O (g8908), .I1 (g8079), .I2 (g8066), .I3 (g8855));
OR4X1 gate7401(.O (I14772), .I1 (g7937), .I2 (g7887), .I3 (g8029), .I4 (g8018));
OR4X1 gate7402(.O (I15232), .I1 (I15228), .I2 (I15229), .I3 (I15230), .I4 (I15231));
OR4X1 gate7403(.O (I15261), .I1 (g8256), .I2 (g8271), .I3 (g8267), .I4 (g8286));
OR2X1 gate7404(.O (g6927), .I1 (g6408), .I2 (g6413));
OR2X1 gate7405(.O (g9171), .I1 (g9146), .I2 (g8962));
OR4X1 gate7406(.O (g8965), .I1 (g8739), .I2 (g8742), .I3 (g8914), .I4 (g8847));
OR2X1 gate7407(.O (g5220), .I1 (g5066), .I2 (g4395));
OR2X1 gate7408(.O (g6436), .I1 (g6266), .I2 (g5699));
OR2X1 gate7409(.O (g8996), .I1 (g8936), .I2 (g8838));
OR2X1 gate7410(.O (g9138), .I1 (g8878), .I2 (g9119));
OR2X1 gate7411(.O (g9338), .I1 (g9258), .I2 (g9334));
OR2X1 gate7412(.O (g8777), .I1 (I14969), .I2 (I14970));
OR4X1 gate7413(.O (g9049), .I1 (g8732), .I2 (g8737), .I3 (g9015), .I4 (g8861));
OR4X1 gate7414(.O (I15031), .I1 (g7951), .I2 (g7920), .I3 (g7983), .I4 (g8181));
OR2X1 gate7415(.O (g8981), .I1 (g8921), .I2 (g8816));
OR3X1 gate7416(.O (g1690), .I1 (g1021), .I2 (g1025), .I3 (g1018));
OR2X1 gate7417(.O (g8997), .I1 (g8937), .I2 (g8841));
OR2X1 gate7418(.O (g6579), .I1 (g6098), .I2 (g1975));
OR2X1 gate7419(.O (g7088), .I1 (g6638), .I2 (g6641));
OR2X1 gate7420(.O (g6719), .I1 (g6166), .I2 (g6171));
OR2X1 gate7421(.O (g6917), .I1 (g6743), .I2 (g6753));
OR2X1 gate7422(.O (g9162), .I1 (g9158), .I2 (g9022));
OR4X1 gate7423(.O (g4735), .I1 (g4427), .I2 (g4414), .I3 (g4403), .I4 (I9041));
OR4X1 gate7424(.O (g9052), .I1 (g8728), .I2 (g8733), .I3 (g9014), .I4 (g8679));
OR2X1 gate7425(.O (g5210), .I1 (g5045), .I2 (g4385));
OR4X1 gate7426(.O (g2262), .I1 (g1384), .I2 (g1385), .I3 (g1386), .I4 (g1387));
OR4X1 gate7427(.O (I15043), .I1 (g8363), .I2 (g8342), .I3 (g8407), .I4 (g8386));
OR2X1 gate7428(.O (g7825), .I1 (g4801), .I2 (g7615));
OR2X1 gate7429(.O (g3760), .I1 (I7232), .I2 (I7233));
OR3X1 gate7430(.O (I9041), .I1 (g4483), .I2 (g4466), .I3 (g4445));
OR3X1 gate7431(.O (g5317), .I1 (g4727), .I2 (g4737), .I3 (g4735));
OR4X1 gate7432(.O (I14952), .I1 (g8456), .I2 (g8513), .I3 (g8458), .I4 (g8236));
OR2X1 gate7433(.O (g6706), .I1 (g4077), .I2 (g6002));
OR2X1 gate7434(.O (g7230), .I1 (g4190), .I2 (g6995));
OR2X1 gate7435(.O (g9006), .I1 (g8946), .I2 (g8853));
OR3X1 gate7436(.O (g8889), .I1 (I15283), .I2 (I15284), .I3 (I15285));
OR3X1 gate7437(.O (I14834), .I1 (g8483), .I2 (g8464), .I3 (g8514));
OR2X1 gate7438(.O (g7337), .I1 (g7278), .I2 (g4546));
OR2X1 gate7439(.O (g6138), .I1 (g5438), .I2 (g5442));
OR4X1 gate7440(.O (I15086), .I1 (I15082), .I2 (I15083), .I3 (I15084), .I4 (I15085));
OR2X1 gate7441(.O (g6707), .I1 (g6160), .I2 (g5585));
OR4X1 gate7442(.O (g8795), .I1 (g8151), .I2 (g8077), .I3 (g8075), .I4 (g8279));
OR2X1 gate7443(.O (g7248), .I1 (g7079), .I2 (g5652));
OR2X1 gate7444(.O (g1955), .I1 (g1189), .I2 (g16));
OR2X1 gate7445(.O (g5704), .I1 (g4936), .I2 (g4334));
OR2X1 gate7446(.O (g9007), .I1 (g8947), .I2 (g8854));
OR2X1 gate7447(.O (g7081), .I1 (g6172), .I2 (g6629));
OR2X1 gate7448(.O (g9261), .I1 (g9238), .I2 (g6227));
OR2X1 gate7449(.O (g8634), .I1 (g6047), .I2 (g8060));
OR4X1 gate7450(.O (I15017), .I1 (g8131), .I2 (g8111), .I3 (g8042), .I4 (g8156));
OR2X1 gate7451(.O (g7783), .I1 (g4787), .I2 (g7600));
OR2X1 gate7452(.O (g8613), .I1 (g8082), .I2 (g7616));
OR2X1 gate7453(.O (g8983), .I1 (g8923), .I2 (g8821));
OR2X1 gate7454(.O (g4876), .I1 (g4159), .I2 (g4167));
OR2X1 gate7455(.O (g6728), .I1 (g6168), .I2 (g5593));
OR2X1 gate7456(.O (g6470), .I1 (g5817), .I2 (g2934));
OR3X1 gate7457(.O (g8885), .I1 (g8723), .I2 (g8806), .I3 (I15243));
OR4X1 gate7458(.O (I7232), .I1 (g2367), .I2 (g2352), .I3 (g2378), .I4 (g2330));
OR2X1 gate7459(.O (g9165), .I1 (g9159), .I2 (g9023));
OR4X1 gate7460(.O (I15042), .I1 (g7951), .I2 (g7920), .I3 (g7983), .I4 (g8181));
OR4X1 gate7461(.O (g9055), .I1 (g8721), .I2 (g8725), .I3 (g9012), .I4 (g8859));
OR2X1 gate7462(.O (g6445), .I1 (g6105), .I2 (g6107));
OR3X1 gate7463(.O (g7258), .I1 (g7083), .I2 (g5403), .I3 (I13220));
OR2X1 gate7464(.O (g6602), .I1 (g6058), .I2 (g3092));
OR2X1 gate7465(.O (g4295), .I1 (g2828), .I2 (g2668));
OR4X1 gate7466(.O (I15030), .I1 (g7855), .I2 (g7838), .I3 (g7905), .I4 (g7870));
OR2X1 gate7467(.O (g6920), .I1 (g6395), .I2 (g6399));
OR2X1 gate7468(.O (g5561), .I1 (g4168), .I2 (g4797));
OR3X1 gate7469(.O (g6459), .I1 (g6259), .I2 (g6185), .I3 (I11603));
OR2X1 gate7470(.O (g6718), .I1 (g4083), .I2 (g6006));
OR2X1 gate7471(.O (g7026), .I1 (g4186), .I2 (g6554));
OR4X1 gate7472(.O (I14933), .I1 (g8385), .I2 (g8404), .I3 (g8441), .I4 (g8462));
OR3X1 gate7473(.O (g7426), .I1 (g1173), .I2 (g7217), .I3 (I13553));
OR2X1 gate7474(.O (g7170), .I1 (g6916), .I2 (g6444));
OR3X1 gate7475(.O (g7083), .I1 (g5448), .I2 (g6267), .I3 (g6710));
OR4X1 gate7476(.O (I15075), .I1 (I15071), .I2 (I15072), .I3 (I15073), .I4 (I15074));
OR2X1 gate7477(.O (g8990), .I1 (g8930), .I2 (g8830));
OR2X1 gate7478(.O (g8888), .I1 (I15276), .I2 (g8807));
OR2X1 gate7479(.O (g7191), .I1 (g7071), .I2 (g6980));
OR2X1 gate7480(.O (g5244), .I1 (g5107), .I2 (g4436));
OR2X1 gate7481(.O (g5140), .I1 (g4333), .I2 (g3509));
OR2X1 gate7482(.O (g7016), .I1 (g6042), .I2 (g6487));
OR2X1 gate7483(.O (g9168), .I1 (g9160), .I2 (g9025));
OR4X1 gate7484(.O (I15276), .I1 (I15272), .I2 (I15273), .I3 (I15274), .I4 (I15275));
OR3X1 gate7485(.O (I15285), .I1 (g8709), .I2 (g8713), .I3 (g8803));
OR2X1 gate7486(.O (g5214), .I1 (g5049), .I2 (g4389));
OR4X1 gate7487(.O (I15053), .I1 (g7951), .I2 (g7920), .I3 (g7983), .I4 (g8181));
OR4X1 gate7488(.O (I15254), .I1 (I15250), .I2 (I15251), .I3 (I15252), .I4 (I15253));
OR2X1 gate7489(.O (g4249), .I1 (g3617), .I2 (g1639));
OR2X1 gate7490(.O (g3986), .I1 (g202), .I2 (g3129));
OR3X1 gate7491(.O (I14302), .I1 (g6664), .I2 (g3492), .I3 (g979));
OR2X1 gate7492(.O (g9011), .I1 (g6046), .I2 (g8892));
OR4X1 gate7493(.O (I15101), .I1 (g8363), .I2 (g8342), .I3 (g8407), .I4 (g8386));
OR2X1 gate7494(.O (g5236), .I1 (g5092), .I2 (g4423));
OR2X1 gate7495(.O (g7272), .I1 (g6182), .I2 (g7038));
OR2X1 gate7496(.O (g8896), .I1 (g8828), .I2 (g8648));
OR2X1 gate7497(.O (g5222), .I1 (g5068), .I2 (g4397));
OR2X1 gate7498(.O (g4812), .I1 (g2490), .I2 (g4237));
OR2X1 gate7499(.O (g4829), .I1 (g863), .I2 (g4051));
OR2X1 gate7500(.O (g6685), .I1 (g4067), .I2 (g5969));
OR2X1 gate7501(.O (g5237), .I1 (g5093), .I2 (g4424));
OR4X1 gate7502(.O (I15074), .I1 (g8363), .I2 (g8342), .I3 (g8407), .I4 (g8386));
OR4X1 gate7503(.O (I15239), .I1 (g8264), .I2 (g8260), .I3 (g8277), .I4 (g8301));
OR2X1 gate7504(.O (g5194), .I1 (g5018), .I2 (g4367));
OR2X1 gate7505(.O (g9000), .I1 (g8940), .I2 (g8845));
OR2X1 gate7506(.O (g8897), .I1 (g8833), .I2 (g8650));
OR2X1 gate7507(.O (g7166), .I1 (g6437), .I2 (g6914));
OR2X1 gate7508(.O (g5242), .I1 (g5105), .I2 (g4434));
OR2X1 gate7509(.O (g5254), .I1 (g5117), .I2 (g4452));
OR4X1 gate7510(.O (I14932), .I1 (g8278), .I2 (g8329), .I3 (g8461), .I4 (g8382));
OR2X1 gate7511(.O (g6585), .I1 (g3617), .I2 (g6119));
OR2X1 gate7512(.O (g6673), .I1 (g4053), .I2 (g5937));
OR2X1 gate7513(.O (g5212), .I1 (g5047), .I2 (g4387));
OR2X1 gate7514(.O (g7167), .I1 (g6438), .I2 (g6915));
OR3X1 gate7515(.O (g8091), .I1 (g7215), .I2 (g6452), .I3 (I14366));
OR4X1 gate7516(.O (I15083), .I1 (g7855), .I2 (g7838), .I3 (g7905), .I4 (g7870));
OR2X1 gate7517(.O (g5229), .I1 (g5079), .I2 (g4409));
OR4X1 gate7518(.O (I15284), .I1 (g8335), .I2 (g8340), .I3 (g8290), .I4 (g8691));
OR4X1 gate7519(.O (g6458), .I1 (g6184), .I2 (g6259), .I3 (g6174), .I4 (g6214));
OR2X1 gate7520(.O (g7834), .I1 (g7724), .I2 (g6762));
OR2X1 gate7521(.O (g6734), .I1 (g6176), .I2 (g5599));
OR2X1 gate7522(.O (g4870), .I1 (g4154), .I2 (g3081));
OR2X1 gate7523(.O (g7687), .I1 (g6053), .I2 (g7416));
OR2X1 gate7524(.O (g6688), .I1 (g6145), .I2 (g5570));
OR4X1 gate7525(.O (I15052), .I1 (g7855), .I2 (g7838), .I3 (g7905), .I4 (g7870));
OR4X1 gate7526(.O (I14959), .I1 (g8322), .I2 (g8308), .I3 (g8438), .I4 (g8612));
OR2X1 gate7527(.O (g5708), .I1 (g2889), .I2 (g4699));
OR2X1 gate7528(.O (g5219), .I1 (g5065), .I2 (g4394));
OR2X1 gate7529(.O (g6924), .I1 (g6400), .I2 (g6405));
OR3X1 gate7530(.O (I15400), .I1 (g8736), .I2 (g8748), .I3 (g8740));
OR2X1 gate7531(.O (g9294), .I1 (g9274), .I2 (g6230));
OR3X1 gate7532(.O (g8758), .I1 (g8655), .I2 (I14932), .I3 (I14933));
OR2X1 gate7533(.O (g9356), .I1 (g9277), .I2 (g9346));
OR2X1 gate7534(.O (g7020), .I1 (g3617), .I2 (g6578));
OR4X1 gate7535(.O (I15241), .I1 (g8269), .I2 (g8314), .I3 (g8309), .I4 (g8695));
OR4X1 gate7536(.O (I15100), .I1 (g7951), .I2 (g7920), .I3 (g7983), .I4 (g8181));
OR2X1 gate7537(.O (g9363), .I1 (g9359), .I2 (g6210));
OR2X1 gate7538(.O (g6116), .I1 (g5546), .I2 (g4681));
OR3X1 gate7539(.O (g6565), .I1 (g2396), .I2 (g6131), .I3 (g1603));
OR2X1 gate7540(.O (g8994), .I1 (g8934), .I2 (g8836));
OR2X1 gate7541(.O (g5245), .I1 (g5108), .I2 (g4437));
OR2X1 gate7542(.O (g9357), .I1 (g9278), .I2 (g9347));
OR2X1 gate7543(.O (g3192), .I1 (g1756), .I2 (g530));
OR4X1 gate7544(.O (g4727), .I1 (g4417), .I2 (g4172), .I3 (g4163), .I4 (I9029));
OR2X1 gate7545(.O (g7040), .I1 (g6439), .I2 (g5783));
OR2X1 gate7546(.O (g5259), .I1 (g5122), .I2 (g4472));
OR3X1 gate7547(.O (I14831), .I1 (g8483), .I2 (g8464), .I3 (g8514));
OR3X1 gate7548(.O (I9038), .I1 (g4507), .I2 (g4497), .I3 (g4486));
OR4X1 gate7549(.O (I15082), .I1 (g8131), .I2 (g8111), .I3 (g8042), .I4 (g8156));
OR2X1 gate7550(.O (g5215), .I1 (g5050), .I2 (g4390));
OR4X1 gate7551(.O (I14753), .I1 (g7993), .I2 (g7966), .I3 (g7793), .I4 (g7811));
OR2X1 gate7552(.O (g2368), .I1 (I6208), .I2 (I6209));
OR2X1 gate7553(.O (g4747), .I1 (g3984), .I2 (g2912));
OR3X1 gate7554(.O (I13220), .I1 (g58), .I2 (g6258), .I3 (g5418));
OR4X1 gate7555(.O (I15263), .I1 (g8313), .I2 (g8297), .I3 (g8310), .I4 (g8690));
OR2X1 gate7556(.O (g6739), .I1 (g4099), .I2 (g6021));
OR4X1 gate7557(.O (I5757), .I1 (g969), .I2 (g970), .I3 (g966), .I4 (g963));
OR3X1 gate7558(.O (I8363), .I1 (g2655), .I2 (g1163), .I3 (g1160));
OR4X1 gate7559(.O (I14960), .I1 (g8621), .I2 (g8622), .I3 (g8628), .I4 (g8230));
OR2X1 gate7560(.O (g5228), .I1 (g5078), .I2 (g4408));
OR2X1 gate7561(.O (g5230), .I1 (g5080), .I2 (g4410));
OR3X1 gate7562(.O (g8890), .I1 (I15290), .I2 (I15291), .I3 (I15292));
OR4X1 gate7563(.O (I15273), .I1 (g8287), .I2 (g8334), .I3 (g8295), .I4 (g8339));
OR2X1 gate7564(.O (g5195), .I1 (g5019), .I2 (g4368));
OR2X1 gate7565(.O (g9004), .I1 (g8944), .I2 (g8851));
OR2X1 gate7566(.O (g7202), .I1 (g6028), .I2 (g7071));
OR4X1 gate7567(.O (I15033), .I1 (I15029), .I2 (I15030), .I3 (I15031), .I4 (I15032));
OR2X1 gate7568(.O (g8992), .I1 (g8932), .I2 (g8832));
OR4X1 gate7569(.O (I14970), .I1 (g8457), .I2 (g8383), .I3 (g8626), .I4 (g8233));
OR2X1 gate7570(.O (g4280), .I1 (I8224), .I2 (I8225));
OR2X1 gate7571(.O (g6912), .I1 (g4199), .I2 (g6567));
OR2X1 gate7572(.O (g5255), .I1 (g5118), .I2 (g4453));
OR4X1 gate7573(.O (g4790), .I1 (g4185), .I2 (g4131), .I3 (g4129), .I4 (I9107));
OR2X1 gate7574(.O (g6929), .I1 (g6412), .I2 (g6418));
OR2X1 gate7575(.O (g7450), .I1 (g6090), .I2 (g7195));
OR4X1 gate7576(.O (g1872), .I1 (g971), .I2 (g962), .I3 (g972), .I4 (I5757));
OR2X1 gate7577(.O (g5218), .I1 (g5064), .I2 (g4393));
OR2X1 gate7578(.O (g6735), .I1 (g4091), .I2 (g6013));
OR2X1 gate7579(.O (g5830), .I1 (g5714), .I2 (g5142));
OR4X1 gate7580(.O (I15291), .I1 (g8331), .I2 (g8336), .I3 (g8338), .I4 (g8688));
OR4X1 gate7581(.O (I7233), .I1 (g2315), .I2 (g2385), .I3 (g2294), .I4 (g2395));
OR2X1 gate7582(.O (g5221), .I1 (g5067), .I2 (g4396));
OR4X1 gate7583(.O (I15029), .I1 (g8131), .I2 (g8111), .I3 (g8042), .I4 (g8156));
OR2X1 gate7584(.O (g2043), .I1 (g1263), .I2 (g1257));
OR2X1 gate7585(.O (g8999), .I1 (g8939), .I2 (g8843));
OR2X1 gate7586(.O (g8146), .I1 (g6045), .I2 (g7597));
OR4X1 gate7587(.O (I8224), .I1 (g3019), .I2 (g3029), .I3 (g3038), .I4 (g3052));
OR2X1 gate7588(.O (g5716), .I1 (g4962), .I2 (g4356));
OR2X1 gate7589(.O (g6919), .I1 (g6771), .I2 (g6394));
OR2X1 gate7590(.O (g9002), .I1 (g8942), .I2 (g8848));
OR2X1 gate7591(.O (g6952), .I1 (g6633), .I2 (g6204));
OR4X1 gate7592(.O (I15240), .I1 (g8259), .I2 (g8294), .I3 (g8263), .I4 (g8305));
OR4X1 gate7593(.O (I14495), .I1 (g7993), .I2 (g7966), .I3 (g7793), .I4 (g7811));
OR2X1 gate7594(.O (g5241), .I1 (g5104), .I2 (g4433));
OR3X1 gate7595(.O (I14985), .I1 (g8341), .I2 (g8384), .I3 (g8542));
OR2X1 gate7596(.O (g3097), .I1 (g1746), .I2 (g287));
OR4X1 gate7597(.O (I15262), .I1 (g8293), .I2 (g8283), .I3 (g8304), .I4 (g8289));
OR2X1 gate7598(.O (g6925), .I1 (g6402), .I2 (g6407));
OR2X1 gate7599(.O (g6120), .I1 (g3617), .I2 (g5555));
OR2X1 gate7600(.O (g5211), .I1 (g5046), .I2 (g4386));
OR2X1 gate7601(.O (g6906), .I1 (g6715), .I2 (g6726));
OR4X1 gate7602(.O (I15099), .I1 (g7855), .I2 (g7838), .I3 (g7905), .I4 (g7870));
OR4X1 gate7603(.O (I15098), .I1 (g8131), .I2 (g8111), .I3 (g8042), .I4 (g8156));
OR4X1 gate7604(.O (I15251), .I1 (g8302), .I2 (g8288), .I3 (g8311), .I4 (g8296));
OR4X1 gate7605(.O (I15272), .I1 (g8237), .I2 (g8300), .I3 (g8261), .I4 (g8282));
OR2X1 gate7606(.O (g5483), .I1 (g4740), .I2 (g4098));
OR4X1 gate7607(.O (I15032), .I1 (g8363), .I2 (g8342), .I3 (g8407), .I4 (g8386));
OR2X1 gate7608(.O (g6907), .I1 (g6727), .I2 (g6732));
OR2X1 gate7609(.O (g9009), .I1 (g8949), .I2 (g8858));
OR2X1 gate7610(.O (g8995), .I1 (g8935), .I2 (g8837));
OR3X1 gate7611(.O (I14219), .I1 (g979), .I2 (g7566), .I3 (g1865));
OR2X1 gate7612(.O (g5200), .I1 (g5029), .I2 (g4375));
OR2X1 gate7613(.O (g5345), .I1 (g4736), .I2 (g4734));
OR2X1 gate7614(.O (g5223), .I1 (g5069), .I2 (g4398));
OR4X1 gate7615(.O (I15071), .I1 (g8131), .I2 (g8111), .I3 (g8042), .I4 (g8156));
OR4X1 gate7616(.O (I14467), .I1 (g7993), .I2 (g7966), .I3 (g7793), .I4 (g7811));
OR3X1 gate7617(.O (I15147), .I1 (g8483), .I2 (g8464), .I3 (g8514));
OR2X1 gate7618(.O (g6590), .I1 (g3617), .I2 (g6153));
OR3X1 gate7619(.O (I15172), .I1 (g8483), .I2 (g8464), .I3 (g8514));
OR2X1 gate7620(.O (g6928), .I1 (g6409), .I2 (g6415));
OR2X1 gate7621(.O (g6930), .I1 (g6414), .I2 (g6420));
OR2X1 gate7622(.O (g5537), .I1 (g3617), .I2 (g4835));
OR2X1 gate7623(.O (g7436), .I1 (g7183), .I2 (g6975));
OR2X1 gate7624(.O (g5243), .I1 (g5106), .I2 (g4435));
OR2X1 gate7625(.O (g5234), .I1 (g5090), .I2 (g4421));
OR4X1 gate7626(.O (I15044), .I1 (I15040), .I2 (I15041), .I3 (I15042), .I4 (I15043));
OR2X1 gate7627(.O (g6705), .I1 (g6157), .I2 (g5583));
OR2X1 gate7628(.O (g8894), .I1 (g8817), .I2 (g8645));
OR3X1 gate7629(.O (g8782), .I1 (g8624), .I2 (g8659), .I3 (I14980));
OR2X1 gate7630(.O (g9005), .I1 (g8945), .I2 (g8852));
OR2X1 gate7631(.O (g5213), .I1 (g5048), .I2 (g4388));
OR4X1 gate7632(.O (I15290), .I1 (g8285), .I2 (g8266), .I3 (g8318), .I4 (g8326));
OR4X1 gate7633(.O (g4374), .I1 (g1182), .I2 (g1186), .I3 (g1179), .I4 (I8363));
OR2X1 gate7634(.O (g8998), .I1 (g8938), .I2 (g8842));
OR2X1 gate7635(.O (g9124), .I1 (g8876), .I2 (g9038));
OR2X1 gate7636(.O (g5698), .I1 (g5057), .I2 (g5040));
OR4X1 gate7637(.O (I14485), .I1 (g7937), .I2 (g7887), .I3 (g8029), .I4 (g8018));
OR2X1 gate7638(.O (g5260), .I1 (g5123), .I2 (g4473));
OR2X1 gate7639(.O (g9377), .I1 (g9371), .I2 (g6757));
OR2X1 gate7640(.O (g6921), .I1 (g6396), .I2 (g6401));
OR2X1 gate7641(.O (g8986), .I1 (g8926), .I2 (g8825));
OR4X1 gate7642(.O (I15297), .I1 (g8280), .I2 (g8257), .I3 (g8319), .I4 (g8327));
ND2X1 gate7643(.O (I15888), .I1 (g9192), .I2 (I15887));
ND2X1 gate7644(.O (I7466), .I1 (g2982), .I2 (g1704));
ND2X1 gate7645(.O (I10092), .I1 (g4881), .I2 (g2177));
ND2X1 gate7646(.O (g5686), .I1 (g5132), .I2 (g1263));
ND2X1 gate7647(.O (I5521), .I1 (g1098), .I2 (I5519));
ND2X1 gate7648(.O (g4528), .I1 (I8606), .I2 (I8607));
ND2X1 gate7649(.O (g5625), .I1 (g2044), .I2 (g4957));
ND2X1 gate7650(.O (I7538), .I1 (g2996), .I2 (g1715));
ND2X1 gate7651(.O (I11143), .I1 (g5493), .I2 (I11142));
ND2X1 gate7652(.O (I7467), .I1 (g2982), .I2 (I7466));
ND2X1 gate7653(.O (g4839), .I1 (g1879), .I2 (g4269));
ND2X1 gate7654(.O (I10906), .I1 (g5492), .I2 (g2605));
ND2X1 gate7655(.O (I12575), .I1 (g6574), .I2 (g1049));
ND2X1 gate7656(.O (I7181), .I1 (g795), .I2 (I7179));
ND2X1 gate7657(.O (g4235), .I1 (g1415), .I2 (g2668));
ND2X1 gate7658(.O (g6286), .I1 (I11178), .I2 (I11179));
ND2X1 gate7659(.O (I7421), .I1 (g2525), .I2 (g2703));
ND2X1 gate7660(.O (g5141), .I1 (I9548), .I2 (I9549));
ND2X1 gate7661(.O (g6911), .I1 (I12597), .I2 (I12598));
ND2X1 gate7662(.O (g4548), .I1 (I8636), .I2 (I8637));
ND2X1 gate7663(.O (I15855), .I1 (g9168), .I2 (g9165));
ND2X1 gate7664(.O (I11110), .I1 (g2734), .I2 (I11108));
ND2X1 gate7665(.O (I11179), .I1 (g3019), .I2 (I11177));
ND2X1 gate7666(.O (g6473), .I1 (g5269), .I2 (g5988));
ND2X1 gate7667(.O (I6524), .I1 (g1102), .I2 (I6522));
ND2X1 gate7668(.O (I11178), .I1 (g5466), .I2 (I11177));
ND2X1 gate7669(.O (I8510), .I1 (g2517), .I2 (g2807));
ND2X1 gate7670(.O (I8245), .I1 (g3506), .I2 (I8243));
ND2X1 gate7671(.O (g4313), .I1 (g3712), .I2 (g3700));
ND2X1 gate7672(.O (I11186), .I1 (g3029), .I2 (I11184));
ND2X1 gate7673(.O (g6469), .I1 (g5918), .I2 (g5278));
ND2X1 gate7674(.O (I13685), .I1 (g1977), .I2 (g7237));
ND2X1 gate7675(.O (I6258), .I1 (g837), .I2 (I6257));
ND2X1 gate7676(.O (g6177), .I1 (I10889), .I2 (I10890));
ND2X1 gate7677(.O (I13800), .I1 (g7429), .I2 (g1061));
ND2X1 gate7678(.O (I15819), .I1 (g9148), .I2 (I15817));
ND2X1 gate7679(.O (I15818), .I1 (g9151), .I2 (I15817));
ND2X1 gate7680(.O (I5600), .I1 (g1489), .I2 (I5598));
ND2X1 gate7681(.O (g6287), .I1 (I11185), .I2 (I11186));
ND2X1 gate7682(.O (I9978), .I1 (g4880), .I2 (g2092));
ND2X1 gate7683(.O (I9243), .I1 (g4305), .I2 (I9241));
ND2X1 gate7684(.O (I6274), .I1 (g840), .I2 (I6273));
ND3X1 gate7685(.O (g5284), .I1 (g4344), .I2 (g4335), .I3 (g4963));
ND2X1 gate7686(.O (I10745), .I1 (g2100), .I2 (I10743));
ND2X1 gate7687(.O (g5239), .I1 (I9746), .I2 (I9747));
ND2X1 gate7688(.O (I9234), .I1 (g4310), .I2 (I9233));
ND2X1 gate7689(.O (I6170), .I1 (g843), .I2 (g911));
ND2X1 gate7690(.O (I13587), .I1 (g2556), .I2 (g7234));
ND2X1 gate7691(.O (g6510), .I1 (g5278), .I2 (g5874));
ND2X1 gate7692(.O (I6939), .I1 (g2161), .I2 (g2051));
ND2X1 gate7693(.O (I11117), .I1 (g3062), .I2 (I11115));
ND2X1 gate7694(.O (g5559), .I1 (g5132), .I2 (g1257));
ND2X1 gate7695(.O (g3232), .I1 (g2298), .I2 (g2276));
ND2X1 gate7696(.O (I7531), .I1 (g2487), .I2 (g3787));
ND2X1 gate7697(.O (g3938), .I1 (I7610), .I2 (I7611));
ND2X1 gate7698(.O (I7505), .I1 (g3802), .I2 (I7503));
ND2X1 gate7699(.O (I7011), .I1 (g2333), .I2 (I7009));
ND2X1 gate7700(.O (I11123), .I1 (g5517), .I2 (I11122));
ND2X1 gate7701(.O (I11751), .I1 (g6112), .I2 (I11750));
ND2X1 gate7702(.O (g6701), .I1 (I12032), .I2 (I12033));
ND2X1 gate7703(.O (g4835), .I1 (I9195), .I2 (I9196));
ND2X1 gate7704(.O (I13639), .I1 (g7257), .I2 (I13638));
ND2X1 gate7705(.O (I10329), .I1 (g2562), .I2 (I10327));
ND2X1 gate7706(.O (g6215), .I1 (I10981), .I2 (I10982));
ND2X1 gate7707(.O (I6904), .I1 (g2105), .I2 (g1838));
ND2X1 gate7708(.O (I13638), .I1 (g7257), .I2 (g7069));
ND2X1 gate7709(.O (I10328), .I1 (g5467), .I2 (I10327));
ND2X1 gate7710(.O (g5750), .I1 (I10314), .I2 (I10315));
ND2X1 gate7711(.O (I7480), .I1 (g3808), .I2 (I7478));
ND2X1 gate7712(.O (I11841), .I1 (g2548), .I2 (g6158));
ND2X1 gate7713(.O (I7569), .I1 (g3780), .I2 (I7567));
ND2X1 gate7714(.O (I9964), .I1 (g1938), .I2 (I9963));
ND2X1 gate7715(.O (g3525), .I1 (I7010), .I2 (I7011));
ND2X1 gate7716(.O (g4332), .I1 (g3681), .I2 (g2368));
ND2X1 gate7717(.O (g7535), .I1 (I13786), .I2 (I13787));
ND2X1 gate7718(.O (I6757), .I1 (g186), .I2 (g1983));
ND2X1 gate7719(.O (I12051), .I1 (g5956), .I2 (g5939));
ND2X1 gate7720(.O (g3358), .I1 (I6940), .I2 (I6941));
ND2X1 gate7721(.O (I11116), .I1 (g5481), .I2 (I11115));
ND2X1 gate7722(.O (I11615), .I1 (g6239), .I2 (I11614));
ND2X1 gate7723(.O (I6522), .I1 (g1919), .I2 (g1102));
ND2X1 gate7724(.O (I9057), .I1 (g4059), .I2 (g1504));
ND2X1 gate7725(.O (I10991), .I1 (g5632), .I2 (g2389));
ND2X1 gate7726(.O (I9549), .I1 (g4307), .I2 (I9547));
ND2X1 gate7727(.O (I8255), .I1 (g3825), .I2 (I8253));
ND2X1 gate7728(.O (g4492), .I1 (I8537), .I2 (I8538));
ND3X1 gate7729(.O (g4714), .I1 (g4344), .I2 (g4335), .I3 (g4328));
ND2X1 gate7730(.O (I11142), .I1 (g5493), .I2 (g3062));
ND2X1 gate7731(.O (I7423), .I1 (g2703), .I2 (I7421));
ND2X1 gate7732(.O (I11165), .I1 (g3029), .I2 (I11163));
ND2X1 gate7733(.O (I6234), .I1 (g896), .I2 (I6232));
ND2X1 gate7734(.O (I10744), .I1 (g5550), .I2 (I10743));
ND2X1 gate7735(.O (g5555), .I1 (I9979), .I2 (I9980));
ND2X1 gate7736(.O (I10849), .I1 (g2595), .I2 (I10847));
ND2X1 gate7737(.O (g4889), .I1 (I9242), .I2 (I9243));
ND2X1 gate7738(.O (g4476), .I1 (I8511), .I2 (I8512));
ND2X1 gate7739(.O (g6142), .I1 (I10790), .I2 (I10791));
ND2X1 gate7740(.O (I10848), .I1 (g5490), .I2 (I10847));
ND4X1 gate7741(.O (g4871), .I1 (g3635), .I2 (g3605), .I3 (g4220), .I4 (g3644));
ND2X1 gate7742(.O (g6497), .I1 (g5278), .I2 (g5847));
ND2X1 gate7743(.O (I7240), .I1 (g1658), .I2 (I7239));
ND2X1 gate7744(.O (g5567), .I1 (g1879), .I2 (g4883));
ND2X1 gate7745(.O (I10361), .I1 (g1118), .I2 (I10359));
ND2X1 gate7746(.O (I7443), .I1 (g2973), .I2 (g1701));
ND2X1 gate7747(.O (I13600), .I1 (g7244), .I2 (I13598));
ND2X1 gate7748(.O (I9691), .I1 (g5096), .I2 (g1037));
ND2X1 gate7749(.O (g6218), .I1 (I10992), .I2 (I10993));
ND2X1 gate7750(.O (g4231), .I1 (g2276), .I2 (g3258));
ND2X1 gate7751(.O (I11137), .I1 (g3052), .I2 (I11135));
ND2X1 gate7752(.O (I7533), .I1 (g3787), .I2 (I7531));
ND2X1 gate7753(.O (I11873), .I1 (g2543), .I2 (g6187));
ND2X1 gate7754(.O (I12552), .I1 (g1462), .I2 (I12550));
ND2X1 gate7755(.O (I9985), .I1 (g4836), .I2 (g2096));
ND2X1 gate7756(.O (I11614), .I1 (g6239), .I2 (g1519));
ND2X1 gate7757(.O (g7093), .I1 (I12870), .I2 (I12871));
ND2X1 gate7758(.O (g9191), .I1 (I15856), .I2 (I15857));
ND2X1 gate7759(.O (I6843), .I1 (g205), .I2 (I6842));
ND2X1 gate7760(.O (I8119), .I1 (g1904), .I2 (g3220));
ND2X1 gate7761(.O (I11122), .I1 (g5517), .I2 (g2712));
ND2X1 gate7762(.O (I8152), .I1 (g38), .I2 (I8150));
ND2X1 gate7763(.O (I7460), .I1 (g2506), .I2 (I7459));
ND2X1 gate7764(.O (I14473), .I1 (g8147), .I2 (I14472));
ND2X1 gate7765(.O (I10789), .I1 (g5512), .I2 (g2170));
ND2X1 gate7766(.O (I7937), .I1 (g3614), .I2 (g1138));
ND2X1 gate7767(.O (I11136), .I1 (g5476), .I2 (I11135));
ND2X1 gate7768(.O (I6232), .I1 (g834), .I2 (g896));
ND2X1 gate7769(.O (I7479), .I1 (g2502), .I2 (I7478));
ND2X1 gate7770(.O (I10359), .I1 (g5552), .I2 (g1118));
ND2X1 gate7771(.O (I6813), .I1 (g210), .I2 (g2052));
ND2X1 gate7772(.O (g1759), .I1 (I5599), .I2 (I5600));
ND2X1 gate7773(.O (g5558), .I1 (I10000), .I2 (I10001));
ND2X1 gate7774(.O (I6740), .I1 (g195), .I2 (I6739));
ND2X1 gate7775(.O (g4513), .I1 (I8582), .I2 (I8583));
ND2X1 gate7776(.O (I11164), .I1 (g5469), .I2 (I11163));
ND2X1 gate7777(.O (I8939), .I1 (g4239), .I2 (I8938));
ND2X1 gate7778(.O (g6119), .I1 (I10744), .I2 (I10745));
ND2X1 gate7779(.O (g7257), .I1 (I13214), .I2 (I13215));
ND2X1 gate7780(.O (I7156), .I1 (g2331), .I2 (g929));
ND2X1 gate7781(.O (g4679), .I1 (I8939), .I2 (I8940));
ND2X1 gate7782(.O (I11575), .I1 (g5894), .I2 (I11574));
ND2X1 gate7783(.O (g3518), .I1 (I6997), .I2 (I6998));
ND2X1 gate7784(.O (I8636), .I1 (g2481), .I2 (I8635));
ND3X1 gate7785(.O (g4831), .I1 (g3635), .I2 (g3605), .I3 (g4220));
ND2X1 gate7786(.O (I11109), .I1 (g5522), .I2 (I11108));
ND2X1 gate7787(.O (g6893), .I1 (I12551), .I2 (I12552));
ND2X1 gate7788(.O (I11108), .I1 (g5522), .I2 (g2734));
ND2X1 gate7789(.O (g6274), .I1 (I11102), .I2 (I11103));
ND2X1 gate7790(.O (I9151), .I1 (g3883), .I2 (g1649));
ND2X1 gate7791(.O (I7453), .I1 (g3226), .I2 (I7452));
ND2X1 gate7792(.O (g6170), .I1 (I10874), .I2 (I10875));
ND2X1 gate7793(.O (I11750), .I1 (g6112), .I2 (g1486));
ND2X1 gate7794(.O (I7568), .I1 (g2481), .I2 (I7567));
ND2X1 gate7795(.O (g6280), .I1 (I11136), .I2 (I11137));
ND2X1 gate7796(.O (I7157), .I1 (g2331), .I2 (I7156));
ND2X1 gate7797(.O (I8637), .I1 (g2743), .I2 (I8635));
ND2X1 gate7798(.O (g4869), .I1 (g4254), .I2 (g3533));
ND2X1 gate7799(.O (I8536), .I1 (g2506), .I2 (g2798));
ND2X1 gate7800(.O (I9278), .I1 (g4313), .I2 (I9276));
ND2X1 gate7801(.O (g3658), .I1 (I7149), .I2 (I7150));
ND3X1 gate7802(.O (g6187), .I1 (g5633), .I2 (g3735), .I3 (g3716));
ND2X1 gate7803(.O (I6275), .I1 (g906), .I2 (I6273));
ND2X1 gate7804(.O (I9235), .I1 (g2180), .I2 (I9233));
ND2X1 gate7805(.O (I10981), .I1 (g5625), .I2 (I10980));
ND2X1 gate7806(.O (g2395), .I1 (I6274), .I2 (I6275));
ND2X1 gate7807(.O (I9693), .I1 (g1037), .I2 (I9691));
ND2X1 gate7808(.O (I9548), .I1 (g1952), .I2 (I9547));
ND2X1 gate7809(.O (g7480), .I1 (I13639), .I2 (I13640));
ND2X1 gate7810(.O (I10899), .I1 (g5520), .I2 (g2752));
ND2X1 gate7811(.O (g1678), .I1 (I5506), .I2 (I5507));
ND2X1 gate7812(.O (I11757), .I1 (g1758), .I2 (g6118));
ND3X1 gate7813(.O (g5672), .I1 (g5056), .I2 (g5039), .I3 (g5023));
ND2X1 gate7814(.O (g6695), .I1 (I12016), .I2 (I12017));
ND2X1 gate7815(.O (g3680), .I1 (I7187), .I2 (I7188));
ND2X1 gate7816(.O (g1682), .I1 (I5520), .I2 (I5521));
ND2X1 gate7817(.O (g6159), .I1 (I10835), .I2 (I10836));
ND2X1 gate7818(.O (I8537), .I1 (g2506), .I2 (I8536));
ND2X1 gate7819(.O (I13397), .I1 (g1057), .I2 (I13395));
ND2X1 gate7820(.O (I6905), .I1 (g2105), .I2 (I6904));
ND2X1 gate7821(.O (I8243), .I1 (g2011), .I2 (g3506));
ND2X1 gate7822(.O (I8328), .I1 (g2721), .I2 (I8326));
ND2X1 gate7823(.O (g2783), .I1 (I6523), .I2 (I6524));
ND2X1 gate7824(.O (I9965), .I1 (g4869), .I2 (I9963));
ND2X1 gate7825(.O (I6750), .I1 (g1733), .I2 (g1494));
ND2X1 gate7826(.O (I13213), .I1 (g7065), .I2 (g7082));
ND2X1 gate7827(.O (g5712), .I1 (I10224), .I2 (I10225));
ND2X1 gate7828(.O (g4745), .I1 (I9070), .I2 (I9071));
ND2X1 gate7829(.O (I11574), .I1 (g5894), .I2 (g1122));
ND3X1 gate7830(.O (g4309), .I1 (g3002), .I2 (g3124), .I3 (g3659));
ND2X1 gate7831(.O (I10061), .I1 (g4910), .I2 (I10060));
ND2X1 gate7832(.O (I7616), .I1 (g3008), .I2 (g1721));
ND2X1 gate7833(.O (I8512), .I1 (g2807), .I2 (I8510));
ND2X1 gate7834(.O (g3889), .I1 (I7437), .I2 (I7438));
ND2X1 gate7835(.O (I10360), .I1 (g5552), .I2 (I10359));
ND2X1 gate7836(.O (I8166), .I1 (g3231), .I2 (I8164));
ND2X1 gate7837(.O (I7503), .I1 (g2498), .I2 (g3802));
ND2X1 gate7838(.O (g3722), .I1 (I7215), .I2 (I7216));
ND2X1 gate7839(.O (g4575), .I1 (I8679), .I2 (I8680));
ND2X1 gate7840(.O (I15863), .I1 (g9174), .I2 (I15862));
ND2X1 gate7841(.O (I13396), .I1 (g7212), .I2 (I13395));
ND2X1 gate7842(.O (I14472), .I1 (g8147), .I2 (g1069));
ND2X1 gate7843(.O (I14246), .I1 (g1065), .I2 (I14244));
ND2X1 gate7844(.O (I7277), .I1 (g2497), .I2 (g1898));
ND2X1 gate7845(.O (I10071), .I1 (g4954), .I2 (g2253));
ND2X1 gate7846(.O (I6172), .I1 (g911), .I2 (I6170));
ND2X1 gate7847(.O (I7617), .I1 (g3008), .I2 (I7616));
ND2X1 gate7848(.O (g6902), .I1 (I12576), .I2 (I12577));
ND2X1 gate7849(.O (I9153), .I1 (g1649), .I2 (I9151));
ND2X1 gate7850(.O (g7316), .I1 (I13377), .I2 (I13378));
ND2X1 gate7851(.O (g3231), .I1 (g1889), .I2 (g1904));
ND2X1 gate7852(.O (I6134), .I1 (g846), .I2 (I6133));
ND2X1 gate7853(.O (I12080), .I1 (g5971), .I2 (I12078));
ND2X1 gate7854(.O (I7892), .I1 (g2979), .I2 (I7891));
ND2X1 gate7855(.O (I8393), .I1 (g2949), .I2 (I8392));
ND2X1 gate7856(.O (g1910), .I1 (g1435), .I2 (g1439));
ND2X1 gate7857(.O (I13787), .I1 (g1477), .I2 (I13785));
ND2X1 gate7858(.O (I12031), .I1 (g5918), .I2 (g5897));
ND2X1 gate7859(.O (g5632), .I1 (g2276), .I2 (g4901));
ND2X1 gate7860(.O (g5095), .I1 (I9476), .I2 (I9477));
ND2X1 gate7861(.O (g4881), .I1 (g2460), .I2 (g4315));
ND2X1 gate7862(.O (g2352), .I1 (I6171), .I2 (I6172));
ND2X1 gate7863(.O (I7140), .I1 (g2397), .I2 (I7138));
ND2X1 gate7864(.O (g6463), .I1 (g5918), .I2 (g5278));
ND2X1 gate7865(.O (I7478), .I1 (g2502), .I2 (g3808));
ND2X1 gate7866(.O (I8121), .I1 (g3220), .I2 (I8119));
ND2X1 gate7867(.O (I6202), .I1 (g831), .I2 (I6201));
ND2X1 gate7868(.O (I13640), .I1 (g7069), .I2 (I13638));
ND2X1 gate7869(.O (g3613), .I1 (I7086), .I2 (I7087));
ND2X1 gate7870(.O (g5752), .I1 (I10328), .I2 (I10329));
ND2X1 gate7871(.O (I12869), .I1 (g2536), .I2 (g6618));
ND2X1 gate7872(.O (I8253), .I1 (g2454), .I2 (g3825));
ND2X1 gate7873(.O (I8938), .I1 (g4239), .I2 (g1545));
ND2X1 gate7874(.O (I6776), .I1 (g1134), .I2 (I6774));
ND2X1 gate7875(.O (I8606), .I1 (g2487), .I2 (I8605));
ND2X1 gate7876(.O (I7214), .I1 (g815), .I2 (g2091));
ND3X1 gate7877(.O (g4305), .I1 (g3712), .I2 (g3700), .I3 (g3732));
ND2X1 gate7878(.O (I9476), .I1 (g4038), .I2 (I9475));
ND2X1 gate7879(.O (I13003), .I1 (g7010), .I2 (I13002));
ND2X1 gate7880(.O (I6996), .I1 (g2275), .I2 (g2242));
ND2X1 gate7881(.O (g5189), .I1 (I9692), .I2 (I9693));
ND2X1 gate7882(.O (I13786), .I1 (g7427), .I2 (I13785));
ND2X1 gate7883(.O (I6878), .I1 (g1910), .I2 (I6876));
ND2X1 gate7884(.O (g3679), .I1 (I7180), .I2 (I7181));
ND2X1 gate7885(.O (I8607), .I1 (g2764), .I2 (I8605));
ND2X1 gate7886(.O (I8659), .I1 (g2471), .I2 (I8658));
ND2X1 gate7887(.O (I9477), .I1 (g1942), .I2 (I9475));
ND2X1 gate7888(.O (g4227), .I1 (I8133), .I2 (I8134));
ND2X1 gate7889(.O (I6997), .I1 (g2275), .I2 (I6996));
ND2X1 gate7890(.O (I12079), .I1 (g5988), .I2 (I12078));
ND2X1 gate7891(.O (g6570), .I1 (I11751), .I2 (I11752));
ND2X1 gate7892(.O (I12078), .I1 (g5988), .I2 (g5971));
ND2X1 gate7893(.O (I12598), .I1 (g1126), .I2 (I12596));
ND2X1 gate7894(.O (I10889), .I1 (g5590), .I2 (I10888));
ND2X1 gate7895(.O (I10980), .I1 (g5625), .I2 (g2210));
ND2X1 gate7896(.O (I10888), .I1 (g5590), .I2 (g2259));
ND2X1 gate7897(.O (g2315), .I1 (I6103), .I2 (I6104));
ND2X1 gate7898(.O (g4502), .I1 (I8559), .I2 (I8560));
ND4X1 gate7899(.O (g6158), .I1 (g3735), .I2 (g3716), .I3 (g5633), .I4 (g3754));
ND2X1 gate7900(.O (g5575), .I1 (I10039), .I2 (I10040));
ND2X1 gate7901(.O (I11149), .I1 (g5473), .I2 (g3038));
ND2X1 gate7902(.O (I8559), .I1 (g2502), .I2 (I8558));
ND2X1 gate7903(.O (g6275), .I1 (I11109), .I2 (I11110));
ND2X1 gate7904(.O (g6615), .I1 (I11842), .I2 (I11843));
ND2X1 gate7905(.O (I7150), .I1 (g1974), .I2 (I7148));
ND2X1 gate7906(.O (g5539), .I1 (I9947), .I2 (I9948));
ND2X1 gate7907(.O (I7438), .I1 (g3822), .I2 (I7436));
ND2X1 gate7908(.O (I7009), .I1 (g2295), .I2 (g2333));
ND2X1 gate7909(.O (I15862), .I1 (g9174), .I2 (g9171));
ND2X1 gate7910(.O (I12017), .I1 (g5847), .I2 (I12015));
ND2X1 gate7911(.O (g6284), .I1 (I11164), .I2 (I11165));
ND2X1 gate7912(.O (g6180), .I1 (I10900), .I2 (I10901));
ND2X1 gate7913(.O (g4741), .I1 (I9058), .I2 (I9059));
ND2X1 gate7914(.O (I9946), .I1 (g2128), .I2 (g4905));
ND2X1 gate7915(.O (g4910), .I1 (g2460), .I2 (g4314));
ND2X1 gate7916(.O (I10625), .I1 (g5314), .I2 (g1514));
ND2X1 gate7917(.O (g2330), .I1 (I6134), .I2 (I6135));
ND2X1 gate7918(.O (g6559), .I1 (g5814), .I2 (g6109));
ND2X1 gate7919(.O (g3012), .I1 (I6758), .I2 (I6759));
ND2X1 gate7920(.O (g9202), .I1 (I15881), .I2 (I15882));
ND2X1 gate7921(.O (g3706), .I1 (g1556), .I2 (g2510));
ND2X1 gate7922(.O (I9182), .I1 (g4231), .I2 (I9181));
ND2X1 gate7923(.O (I9382), .I1 (g4062), .I2 (I9381));
ND2X1 gate7924(.O (I10060), .I1 (g4910), .I2 (g2226));
ND2X1 gate7925(.O (I10197), .I1 (g4724), .I2 (I10196));
ND2X1 gate7926(.O (I6500), .I1 (g1913), .I2 (I6499));
ND2X1 gate7927(.O (I10855), .I1 (g5521), .I2 (I10854));
ND2X1 gate7928(.O (I8151), .I1 (g3229), .I2 (I8150));
ND2X1 gate7929(.O (I13378), .I1 (g1472), .I2 (I13376));
ND2X1 gate7930(.O (I9947), .I1 (g2128), .I2 (I9946));
ND2X1 gate7931(.O (I11096), .I1 (g2734), .I2 (I11094));
ND2X1 gate7932(.O (I10867), .I1 (g5480), .I2 (I10866));
ND2X1 gate7933(.O (I5505), .I1 (g1532), .I2 (g1528));
ND2X1 gate7934(.O (I13802), .I1 (g1061), .I2 (I13800));
ND2X1 gate7935(.O (I10315), .I1 (g1041), .I2 (I10313));
ND3X1 gate7936(.O (g5305), .I1 (g5009), .I2 (g4335), .I3 (g4328));
ND2X1 gate7937(.O (I6523), .I1 (g1919), .I2 (I6522));
ND2X1 gate7938(.O (I10819), .I1 (g5567), .I2 (I10818));
ND2X1 gate7939(.O (I12016), .I1 (g5874), .I2 (I12015));
ND2X1 gate7940(.O (I10818), .I1 (g5567), .I2 (g2039));
ND2X1 gate7941(.O (g5748), .I1 (I10306), .I2 (I10307));
ND2X1 gate7942(.O (I11549), .I1 (g5984), .I2 (g1045));
ND2X1 gate7943(.O (g9179), .I1 (I15818), .I2 (I15819));
ND2X1 gate7944(.O (I7085), .I1 (g1753), .I2 (g1918));
ND2X1 gate7945(.O (I7485), .I1 (g2989), .I2 (g1708));
ND2X1 gate7946(.O (I6104), .I1 (g921), .I2 (I6102));
ND2X1 gate7947(.O (I6499), .I1 (g1913), .I2 (g1537));
ND2X1 gate7948(.O (g4256), .I1 (g3233), .I2 (g1444));
ND2X1 gate7949(.O (I8134), .I1 (g1646), .I2 (I8132));
ND2X1 gate7950(.O (g7503), .I1 (I13686), .I2 (I13687));
ND2X1 gate7951(.O (I10094), .I1 (g2177), .I2 (I10092));
ND2X1 gate7952(.O (I6273), .I1 (g840), .I2 (g906));
ND2X1 gate7953(.O (g2367), .I1 (I6202), .I2 (I6203));
ND2X1 gate7954(.O (g4700), .I1 (g2460), .I2 (g4271));
ND2X1 gate7955(.O (I13002), .I1 (g7010), .I2 (g1053));
ND2X1 gate7956(.O (I9233), .I1 (g4310), .I2 (g2180));
ND2X1 gate7957(.O (I10019), .I1 (g2174), .I2 (I10017));
ND2X1 gate7958(.O (g4263), .I1 (g3260), .I2 (g1435));
ND2X1 gate7959(.O (I10196), .I1 (g4724), .I2 (g1958));
ND2X1 gate7960(.O (I10018), .I1 (g4700), .I2 (I10017));
ND2X1 gate7961(.O (g6282), .I1 (I11150), .I2 (I11151));
ND2X1 gate7962(.O (I10866), .I1 (g5480), .I2 (g2605));
ND2X1 gate7963(.O (I7270), .I1 (g955), .I2 (I7268));
ND2X1 gate7964(.O (I10001), .I1 (g1929), .I2 (I9999));
ND2X1 gate7965(.O (I7610), .I1 (g2471), .I2 (I7609));
ND2X1 gate7966(.O (I9171), .I1 (g4244), .I2 (I9169));
ND2X1 gate7967(.O (I10923), .I1 (g5525), .I2 (g2752));
ND2X1 gate7968(.O (I7069), .I1 (g1639), .I2 (I7068));
ND2X1 gate7969(.O (I10300), .I1 (g2562), .I2 (I10298));
ND3X1 gate7970(.O (g7244), .I1 (g7050), .I2 (g3757), .I3 (g3739));
ND2X1 gate7971(.O (I7540), .I1 (g1715), .I2 (I7538));
ND2X1 gate7972(.O (g7140), .I1 (I13003), .I2 (I13004));
ND2X1 gate7973(.O (g5689), .I1 (I10197), .I2 (I10198));
ND2X1 gate7974(.O (I9745), .I1 (g4826), .I2 (g1549));
ND2X1 gate7975(.O (I9963), .I1 (g1938), .I2 (g4869));
ND2X1 gate7976(.O (g7082), .I1 (I12853), .I2 (I12854));
ND2X1 gate7977(.O (I6135), .I1 (g916), .I2 (I6133));
ND2X1 gate7978(.O (g3678), .I1 (I7173), .I2 (I7174));
ND2X1 gate7979(.O (I15881), .I1 (g9190), .I2 (I15880));
ND2X1 gate7980(.O (I11080), .I1 (g2511), .I2 (I11078));
ND2X1 gate7981(.O (I10854), .I1 (g5521), .I2 (g2584));
ND2X1 gate7982(.O (I6916), .I1 (g2360), .I2 (g1732));
ND2X1 gate7983(.O (g5564), .I1 (I10018), .I2 (I10019));
ND2X1 gate7984(.O (I8658), .I1 (g2471), .I2 (g2724));
ND2X1 gate7985(.O (I5696), .I1 (g1513), .I2 (I5695));
ND2X1 gate7986(.O (I7510), .I1 (g2992), .I2 (g1711));
ND2X1 gate7987(.O (I12853), .I1 (g6701), .I2 (I12852));
ND2X1 gate7988(.O (g4474), .I1 (I8503), .I2 (I8504));
ND2X1 gate7989(.O (I10314), .I1 (g5484), .I2 (I10313));
ND2X1 gate7990(.O (I6102), .I1 (g849), .I2 (g921));
ND2X1 gate7991(.O (I11843), .I1 (g6158), .I2 (I11841));
ND2X1 gate7992(.O (I10307), .I1 (g3019), .I2 (I10305));
ND2X1 gate7993(.O (g5589), .I1 (I10061), .I2 (I10062));
ND2X1 gate7994(.O (I8132), .I1 (g3232), .I2 (g1646));
ND2X1 gate7995(.O (I8680), .I1 (g2706), .I2 (I8678));
ND2X1 gate7996(.O (g3602), .I1 (I7069), .I2 (I7070));
ND2X1 gate7997(.O (I6752), .I1 (g1494), .I2 (I6750));
ND2X1 gate7998(.O (I6917), .I1 (g2360), .I2 (I6916));
ND2X1 gate7999(.O (g1775), .I1 (I5620), .I2 (I5621));
ND2X1 gate8000(.O (I7215), .I1 (g815), .I2 (I7214));
ND2X1 gate8001(.O (g3767), .I1 (I7240), .I2 (I7241));
ND2X1 gate8002(.O (I5697), .I1 (g1524), .I2 (I5695));
ND2X1 gate8003(.O (I8558), .I1 (g2502), .I2 (g2790));
ND2X1 gate8004(.O (I12053), .I1 (g5939), .I2 (I12051));
ND2X1 gate8005(.O (I6233), .I1 (g834), .I2 (I6232));
ND2X1 gate8006(.O (I10335), .I1 (g5462), .I2 (I10334));
ND2X1 gate8007(.O (g9205), .I1 (I15898), .I2 (I15899));
ND2X1 gate8008(.O (I8511), .I1 (g2517), .I2 (I8510));
ND2X1 gate8009(.O (I10993), .I1 (g2389), .I2 (I10991));
ND2X1 gate8010(.O (I14839), .I1 (g1073), .I2 (I14837));
ND2X1 gate8011(.O (g5538), .I1 (g5132), .I2 (g1266));
ND2X1 gate8012(.O (I15897), .I1 (g9202), .I2 (g9203));
ND2X1 gate8013(.O (I14838), .I1 (g8660), .I2 (I14837));
ND2X1 gate8014(.O (g7237), .I1 (g7050), .I2 (g3739));
ND2X1 gate8015(.O (I9070), .I1 (g4400), .I2 (I9069));
ND2X1 gate8016(.O (g6153), .I1 (I10819), .I2 (I10820));
ND2X1 gate8017(.O (g6680), .I1 (g5403), .I2 (g6252));
ND2X1 gate8018(.O (g8239), .I1 (g8073), .I2 (g8092));
ND2X1 gate8019(.O (I11171), .I1 (g5477), .I2 (I11170));
ND2X1 gate8020(.O (I6171), .I1 (g843), .I2 (I6170));
ND2X1 gate8021(.O (I10039), .I1 (g4893), .I2 (I10038));
ND2X1 gate8022(.O (I10306), .I1 (g5470), .I2 (I10305));
ND2X1 gate8023(.O (I10038), .I1 (g4893), .I2 (g2202));
ND2X1 gate8024(.O (g3028), .I1 (I6775), .I2 (I6776));
ND2X1 gate8025(.O (I11079), .I1 (g5697), .I2 (I11078));
ND2X1 gate8026(.O (I7891), .I1 (g2979), .I2 (g1499));
ND2X1 gate8027(.O (I10143), .I1 (g4707), .I2 (I10142));
ND2X1 gate8028(.O (I13599), .I1 (g2551), .I2 (I13598));
ND2X1 gate8029(.O (I11078), .I1 (g5697), .I2 (g2511));
ND2X1 gate8030(.O (I13598), .I1 (g2551), .I2 (g7244));
ND2X1 gate8031(.O (g5562), .I1 (I10010), .I2 (I10011));
ND2X1 gate8032(.O (I10791), .I1 (g2170), .I2 (I10789));
ND2X1 gate8033(.O (I15850), .I1 (g9154), .I2 (I15848));
ND2X1 gate8034(.O (I8339), .I1 (g2966), .I2 (I8338));
ND2X1 gate8035(.O (g5257), .I1 (I9768), .I2 (I9769));
ND2X1 gate8036(.O (I6759), .I1 (g1983), .I2 (I6757));
ND2X1 gate8037(.O (g5605), .I1 (I10093), .I2 (I10094));
ND2X1 gate8038(.O (g3883), .I1 (g2276), .I2 (g3188));
ND2X1 gate8039(.O (I11158), .I1 (g3052), .I2 (I11156));
ND2X1 gate8040(.O (I6201), .I1 (g831), .I2 (g891));
ND2X1 gate8041(.O (I9169), .I1 (g1935), .I2 (g4244));
ND2X1 gate8042(.O (g5751), .I1 (I10321), .I2 (I10322));
ND2X1 gate8043(.O (I9059), .I1 (g1504), .I2 (I9057));
ND2X1 gate8044(.O (g6476), .I1 (g5939), .I2 (g5269));
ND2X1 gate8045(.O (I11144), .I1 (g3062), .I2 (I11142));
ND2X1 gate8046(.O (I9767), .I1 (g4832), .I2 (g1114));
ND2X1 gate8047(.O (g6722), .I1 (I12079), .I2 (I12080));
ND2X1 gate8048(.O (I10223), .I1 (g2522), .I2 (g4895));
ND2X1 gate8049(.O (g6285), .I1 (I11171), .I2 (I11172));
ND2X1 gate8050(.O (I12577), .I1 (g1049), .I2 (I12575));
ND2X1 gate8051(.O (I6539), .I1 (g2555), .I2 (I6538));
ND2X1 gate8052(.O (I10321), .I1 (g5459), .I2 (I10320));
ND2X1 gate8053(.O (I13017), .I1 (g6941), .I2 (I13016));
ND2X1 gate8054(.O (g6424), .I1 (I11550), .I2 (I11551));
ND2X1 gate8055(.O (I10953), .I1 (g5565), .I2 (I10952));
ND2X1 gate8056(.O (I15857), .I1 (g9165), .I2 (I15855));
ND2X1 gate8057(.O (g6477), .I1 (g5269), .I2 (g5918));
ND2X1 gate8058(.O (g4820), .I1 (I9170), .I2 (I9171));
ND2X1 gate8059(.O (I10334), .I1 (g5462), .I2 (g2573));
ND2X1 gate8060(.O (I13687), .I1 (g7237), .I2 (I13685));
ND2X1 gate8061(.O (I11752), .I1 (g1486), .I2 (I11750));
ND2X1 gate8062(.O (I7068), .I1 (g1639), .I2 (g1643));
ND2X1 gate8063(.O (I12852), .I1 (g6701), .I2 (g6695));
ND2X1 gate8064(.O (I7468), .I1 (g1704), .I2 (I7466));
ND2X1 gate8065(.O (g6273), .I1 (I11095), .I2 (I11096));
ND2X1 gate8066(.O (I9826), .I1 (g4729), .I2 (g1509));
ND2X1 gate8067(.O (I8660), .I1 (g2724), .I2 (I8658));
ND2X1 gate8068(.O (I10000), .I1 (g4839), .I2 (I9999));
ND2X1 gate8069(.O (I10908), .I1 (g2605), .I2 (I10906));
ND2X1 gate8070(.O (I11842), .I1 (g2548), .I2 (I11841));
ND2X1 gate8071(.O (I7576), .I1 (g1718), .I2 (I7574));
ND2X1 gate8072(.O (I7149), .I1 (g799), .I2 (I7148));
ND2X1 gate8073(.O (I12576), .I1 (g6574), .I2 (I12575));
ND2X1 gate8074(.O (I13016), .I1 (g6941), .I2 (g1142));
ND2X1 gate8075(.O (g4294), .I1 (I8244), .I2 (I8245));
ND2X1 gate8076(.O (I8679), .I1 (g2467), .I2 (I8678));
ND2X1 gate8077(.O (I7241), .I1 (g2134), .I2 (I7239));
ND2X1 gate8078(.O (I12052), .I1 (g5956), .I2 (I12051));
ND2X1 gate8079(.O (I15856), .I1 (g9168), .I2 (I15855));
ND2X1 gate8080(.O (I15880), .I1 (g9190), .I2 (g9179));
ND2X1 gate8081(.O (I10992), .I1 (g5632), .I2 (I10991));
ND2X1 gate8082(.O (I9827), .I1 (g4729), .I2 (I9826));
ND2X1 gate8083(.O (g7069), .I1 (g5435), .I2 (g6680));
ND2X1 gate8084(.O (I11124), .I1 (g2712), .I2 (I11122));
ND2X1 gate8085(.O (I8560), .I1 (g2790), .I2 (I8558));
ND2X1 gate8086(.O (g4954), .I1 (g4319), .I2 (g2460));
ND2X1 gate8087(.O (g4810), .I1 (I9152), .I2 (I9153));
ND2X1 gate8088(.O (g7540), .I1 (I13801), .I2 (I13802));
ND2X1 gate8089(.O (g4363), .I1 (I8339), .I2 (I8340));
ND2X1 gate8090(.O (I13686), .I1 (g1977), .I2 (I13685));
ND2X1 gate8091(.O (I9196), .I1 (g1652), .I2 (I9194));
ND2X1 gate8092(.O (I10835), .I1 (g5514), .I2 (I10834));
ND2X1 gate8093(.O (g6178), .I1 (g2205), .I2 (g5568));
ND2X1 gate8094(.O (I7893), .I1 (g1499), .I2 (I7891));
ND2X1 gate8095(.O (I7186), .I1 (g2353), .I2 (g1834));
ND2X1 gate8096(.O (I11875), .I1 (g6187), .I2 (I11873));
ND2X1 gate8097(.O (g4912), .I1 (I9277), .I2 (I9278));
ND2X1 gate8098(.O (g3890), .I1 (I7444), .I2 (I7445));
ND2X1 gate8099(.O (I9994), .I1 (g4871), .I2 (I9992));
ND2X1 gate8100(.O (g3011), .I1 (I6751), .I2 (I6752));
ND2X1 gate8101(.O (I7939), .I1 (g1138), .I2 (I7937));
ND2X1 gate8102(.O (I6203), .I1 (g891), .I2 (I6201));
ND2X1 gate8103(.O (I9181), .I1 (g4231), .I2 (g2007));
ND2X1 gate8104(.O (g5753), .I1 (I10335), .I2 (I10336));
ND2X1 gate8105(.O (I8164), .I1 (g1943), .I2 (g3231));
ND2X1 gate8106(.O (I9381), .I1 (g4062), .I2 (g1908));
ND2X1 gate8107(.O (I15887), .I1 (g9192), .I2 (g9191));
ND2X1 gate8108(.O (g7144), .I1 (I13017), .I2 (I13018));
ND2X1 gate8109(.O (I10142), .I1 (g4707), .I2 (g1916));
ND2X1 gate8110(.O (I6940), .I1 (g2161), .I2 (I6939));
ND2X1 gate8111(.O (I7187), .I1 (g2353), .I2 (I7186));
ND2X1 gate8112(.O (I7461), .I1 (g3815), .I2 (I7459));
ND2X1 gate8113(.O (g5565), .I1 (g2044), .I2 (g4933));
ND2X1 gate8114(.O (g5681), .I1 (g5132), .I2 (g2043));
ND2X1 gate8115(.O (g6265), .I1 (I11079), .I2 (I11080));
ND2X1 gate8116(.O (g5697), .I1 (g2044), .I2 (g5005));
ND2X1 gate8117(.O (I11170), .I1 (g5477), .I2 (g3038));
ND2X1 gate8118(.O (g6164), .I1 (I10848), .I2 (I10849));
ND2X1 gate8119(.O (I8956), .I1 (g4246), .I2 (I8955));
ND2X1 gate8120(.O (I6741), .I1 (g1970), .I2 (I6739));
ND2X1 gate8121(.O (g6770), .I1 (I12180), .I2 (I12181));
ND2X1 gate8122(.O (I13589), .I1 (g7234), .I2 (I13587));
ND2X1 gate8123(.O (I13588), .I1 (g2556), .I2 (I13587));
ND2X1 gate8124(.O (I8338), .I1 (g2966), .I2 (g1698));
ND2X1 gate8125(.O (g3924), .I1 (I7568), .I2 (I7569));
ND2X1 gate8126(.O (I10952), .I1 (g5565), .I2 (g2340));
ND2X1 gate8127(.O (I6758), .I1 (g186), .I2 (I6757));
ND2X1 gate8128(.O (I6066), .I1 (g883), .I2 (I6064));
ND2X1 gate8129(.O (g7065), .I1 (I12833), .I2 (I12834));
ND2X1 gate8130(.O (I11616), .I1 (g1519), .I2 (I11614));
ND2X1 gate8131(.O (I10790), .I1 (g5512), .I2 (I10789));
ND2X1 gate8132(.O (I9058), .I1 (g4059), .I2 (I9057));
ND2X1 gate8133(.O (I10873), .I1 (g5516), .I2 (g2595));
ND2X1 gate8134(.O (I8957), .I1 (g1110), .I2 (I8955));
ND2X1 gate8135(.O (g3665), .I1 (I7157), .I2 (I7158));
ND2X1 gate8136(.O (I6133), .I1 (g846), .I2 (g916));
ND2X1 gate8137(.O (g6281), .I1 (I11143), .I2 (I11144));
ND2X1 gate8138(.O (I6774), .I1 (g2386), .I2 (g1134));
ND2X1 gate8139(.O (I11101), .I1 (g5491), .I2 (g2712));
ND2X1 gate8140(.O (I11177), .I1 (g5466), .I2 (g3019));
ND2X1 gate8141(.O (I10834), .I1 (g5514), .I2 (g2584));
ND2X1 gate8142(.O (I6538), .I1 (g2555), .I2 (g2557));
ND2X1 gate8143(.O (I9992), .I1 (g2145), .I2 (g4871));
ND2X1 gate8144(.O (I11874), .I1 (g2543), .I2 (I11873));
ND2X1 gate8145(.O (I15817), .I1 (g9151), .I2 (g9148));
ND2X1 gate8146(.O (I12833), .I1 (g6722), .I2 (I12832));
ND2X1 gate8147(.O (I10320), .I1 (g5459), .I2 (g2573));
ND2X1 gate8148(.O (I10073), .I1 (g2253), .I2 (I10071));
ND2X1 gate8149(.O (g8231), .I1 (I14473), .I2 (I14474));
ND2X1 gate8150(.O (g5363), .I1 (I9827), .I2 (I9828));
ND2X1 gate8151(.O (g3681), .I1 (g866), .I2 (g2368));
ND2X1 gate8152(.O (I8504), .I1 (g2038), .I2 (I8502));
ND2X1 gate8153(.O (g3914), .I1 (I7532), .I2 (I7533));
ND2X1 gate8154(.O (I12951), .I1 (g7003), .I2 (g1467));
ND3X1 gate8155(.O (g5568), .I1 (g2044), .I2 (g4902), .I3 (g4320));
ND2X1 gate8156(.O (I12033), .I1 (g5897), .I2 (I12031));
ND2X1 gate8157(.O (I8470), .I1 (g2525), .I2 (g2821));
ND2X1 gate8158(.O (I7512), .I1 (g1711), .I2 (I7510));
ND2X1 gate8159(.O (g9203), .I1 (I15888), .I2 (I15889));
ND2X1 gate8160(.O (I11185), .I1 (g5474), .I2 (I11184));
ND2X1 gate8161(.O (g4244), .I1 (g3549), .I2 (g3533));
ND2X1 gate8162(.O (I6257), .I1 (g837), .I2 (g901));
ND2X1 gate8163(.O (I7148), .I1 (g799), .I2 (g1974));
ND2X1 gate8164(.O (I9183), .I1 (g2007), .I2 (I9181));
ND2X1 gate8165(.O (I9383), .I1 (g1908), .I2 (I9381));
ND2X1 gate8166(.O (I14474), .I1 (g1069), .I2 (I14472));
ND2X1 gate8167(.O (I8678), .I1 (g2467), .I2 (g2706));
ND2X1 gate8168(.O (I10327), .I1 (g5467), .I2 (g2562));
ND2X1 gate8169(.O (g7828), .I1 (I14245), .I2 (I14246));
ND2X1 gate8170(.O (I8635), .I1 (g2481), .I2 (g2743));
ND2X1 gate8171(.O (I6751), .I1 (g1733), .I2 (I6750));
ND2X1 gate8172(.O (g6504), .I1 (g5269), .I2 (g5874));
ND2X1 gate8173(.O (I13215), .I1 (g7082), .I2 (I13213));
ND2X1 gate8174(.O (g2378), .I1 (I6233), .I2 (I6234));
ND2X1 gate8175(.O (I10982), .I1 (g2210), .I2 (I10980));
ND2X1 gate8176(.O (I7279), .I1 (g1898), .I2 (I7277));
ND2X1 gate8177(.O (I9999), .I1 (g4839), .I2 (g1929));
ND2X1 gate8178(.O (g4110), .I1 (I7938), .I2 (I7939));
ND2X1 gate8179(.O (g4310), .I1 (g3666), .I2 (g2460));
ND2X1 gate8180(.O (g4824), .I1 (I9182), .I2 (I9183));
ND2X1 gate8181(.O (g5661), .I1 (I10143), .I2 (I10144));
ND2X1 gate8182(.O (I8582), .I1 (g2498), .I2 (I8581));
ND2X1 gate8183(.O (I7938), .I1 (g3614), .I2 (I7937));
ND2X1 gate8184(.O (I5620), .I1 (g1092), .I2 (I5619));
ND2X1 gate8185(.O (I10040), .I1 (g2202), .I2 (I10038));
ND2X1 gate8186(.O (g8798), .I1 (g6984), .I2 (g8644));
ND2X1 gate8187(.O (g4563), .I1 (I8659), .I2 (I8660));
ND2X1 gate8188(.O (g6169), .I1 (I10867), .I2 (I10868));
ND2X1 gate8189(.O (g6283), .I1 (I11157), .I2 (I11158));
ND2X1 gate8190(.O (g4237), .I1 (I8151), .I2 (I8152));
ND2X1 gate8191(.O (I11576), .I1 (g1122), .I2 (I11574));
ND2X1 gate8192(.O (I8502), .I1 (g2986), .I2 (g2038));
ND2X1 gate8193(.O (I10847), .I1 (g5490), .I2 (g2595));
ND2X1 gate8194(.O (I8940), .I1 (g1545), .I2 (I8938));
ND2X1 gate8195(.O (I10062), .I1 (g2226), .I2 (I10060));
ND2X1 gate8196(.O (I11115), .I1 (g5481), .I2 (g3062));
ND2X1 gate8197(.O (g5546), .I1 (I9964), .I2 (I9965));
ND2X1 gate8198(.O (g7325), .I1 (I13396), .I2 (I13397));
ND2X1 gate8199(.O (I5520), .I1 (g1087), .I2 (I5519));
ND2X1 gate8200(.O (g6203), .I1 (I10953), .I2 (I10954));
ND2X1 gate8201(.O (I11184), .I1 (g5474), .I2 (g3029));
ND2X1 gate8202(.O (I7158), .I1 (g929), .I2 (I7156));
ND2X1 gate8203(.O (I6924), .I1 (g1728), .I2 (I6923));
ND2X1 gate8204(.O (I12832), .I1 (g6722), .I2 (g6709));
ND2X1 gate8205(.O (I10072), .I1 (g4954), .I2 (I10071));
ND2X1 gate8206(.O (g4836), .I1 (g4288), .I2 (g1879));
ND2X1 gate8207(.O (g3894), .I1 (I7460), .I2 (I7461));
ND2X1 gate8208(.O (g6188), .I1 (I10924), .I2 (I10925));
ND2X1 gate8209(.O (I7174), .I1 (g2006), .I2 (I7172));
ND2X1 gate8210(.O (I13214), .I1 (g7065), .I2 (I13213));
ND2X1 gate8211(.O (I10820), .I1 (g2039), .I2 (I10818));
ND2X1 gate8212(.O (I7239), .I1 (g1658), .I2 (g2134));
ND2X1 gate8213(.O (I8165), .I1 (g1943), .I2 (I8164));
ND2X1 gate8214(.O (I7180), .I1 (g2351), .I2 (I7179));
ND2X1 gate8215(.O (I6103), .I1 (g849), .I2 (I6102));
ND2X1 gate8216(.O (I8133), .I1 (g3232), .I2 (I8132));
ND2X1 gate8217(.O (g1819), .I1 (I5696), .I2 (I5697));
ND2X1 gate8218(.O (I12032), .I1 (g5918), .I2 (I12031));
ND2X1 gate8219(.O (g5035), .I1 (I9382), .I2 (I9383));
ND2X1 gate8220(.O (I9954), .I1 (g2131), .I2 (I9953));
ND2X1 gate8221(.O (I8538), .I1 (g2798), .I2 (I8536));
ND2X1 gate8222(.O (I15864), .I1 (g9171), .I2 (I15862));
ND2X1 gate8223(.O (I12871), .I1 (g6618), .I2 (I12869));
ND2X1 gate8224(.O (g6466), .I1 (I11615), .I2 (I11616));
ND2X1 gate8225(.O (g7447), .I1 (I13599), .I2 (I13600));
ND2X1 gate8226(.O (g6165), .I1 (I10855), .I2 (I10856));
ND2X1 gate8227(.O (g6571), .I1 (I11758), .I2 (I11759));
ND3X1 gate8228(.O (g5310), .I1 (g5009), .I2 (g4335), .I3 (g4963));
ND2X1 gate8229(.O (g4298), .I1 (I8254), .I2 (I8255));
ND2X1 gate8230(.O (I10743), .I1 (g5550), .I2 (g2100));
ND2X1 gate8231(.O (g5762), .I1 (I10360), .I2 (I10361));
ND2X1 gate8232(.O (g3925), .I1 (I7575), .I2 (I7576));
ND2X1 gate8233(.O (g5590), .I1 (g2044), .I2 (g4906));
ND2X1 gate8234(.O (I11759), .I1 (g6118), .I2 (I11757));
ND2X1 gate8235(.O (g5657), .I1 (g5021), .I2 (g4381));
ND2X1 gate8236(.O (I11758), .I1 (g1758), .I2 (I11757));
ND2X1 gate8237(.O (g6467), .I1 (g5956), .I2 (g5269));
ND2X1 gate8238(.O (g5556), .I1 (I9986), .I2 (I9987));
ND2X1 gate8239(.O (g4219), .I1 (I8120), .I2 (I8121));
ND2X1 gate8240(.O (g2385), .I1 (I6258), .I2 (I6259));
ND4X1 gate8241(.O (g7234), .I1 (g3757), .I2 (g3739), .I3 (g7050), .I4 (g3770));
ND2X1 gate8242(.O (g4252), .I1 (g2276), .I2 (g3313));
ND2X1 gate8243(.O (g3906), .I1 (I7504), .I2 (I7505));
ND2X1 gate8244(.O (I6775), .I1 (g2386), .I2 (I6774));
ND2X1 gate8245(.O (I7010), .I1 (g2295), .I2 (I7009));
ND2X1 gate8246(.O (I10890), .I1 (g2259), .I2 (I10888));
ND2X1 gate8247(.O (I8605), .I1 (g2487), .I2 (g2764));
ND2X1 gate8248(.O (g6181), .I1 (I10907), .I2 (I10908));
ND2X1 gate8249(.O (g4911), .I1 (g4320), .I2 (g2044));
ND2X1 gate8250(.O (I9475), .I1 (g4038), .I2 (g1942));
ND2X1 gate8251(.O (I6739), .I1 (g195), .I2 (g1970));
ND2X1 gate8252(.O (I7172), .I1 (g1739), .I2 (g2006));
ND2X1 gate8253(.O (I7278), .I1 (g2497), .I2 (I7277));
ND2X1 gate8254(.O (I11135), .I1 (g5476), .I2 (g3052));
ND2X1 gate8255(.O (I7618), .I1 (g1721), .I2 (I7616));
ND2X1 gate8256(.O (g2801), .I1 (I6539), .I2 (I6540));
ND2X1 gate8257(.O (g5557), .I1 (I9993), .I2 (I9994));
ND2X1 gate8258(.O (g3907), .I1 (I7511), .I2 (I7512));
ND2X1 gate8259(.O (I6501), .I1 (g1537), .I2 (I6499));
ND2X1 gate8260(.O (I13004), .I1 (g1053), .I2 (I13002));
ND2X1 gate8261(.O (I9276), .I1 (g2533), .I2 (g4313));
ND2X1 gate8262(.O (g3656), .I1 (I7139), .I2 (I7140));
ND2X1 gate8263(.O (g3915), .I1 (I7539), .I2 (I7540));
ND2X1 gate8264(.O (g4399), .I1 (I8393), .I2 (I8394));
ND2X1 gate8265(.O (I9986), .I1 (g4836), .I2 (I9985));
ND2X1 gate8266(.O (I7567), .I1 (g2481), .I2 (g3780));
ND2X1 gate8267(.O (I9277), .I1 (g2533), .I2 (I9276));
ND2X1 gate8268(.O (I11163), .I1 (g5469), .I2 (g3029));
ND2X1 gate8269(.O (I12551), .I1 (g6689), .I2 (I12550));
ND2X1 gate8270(.O (g7121), .I1 (I12952), .I2 (I12953));
ND2X1 gate8271(.O (I9987), .I1 (g2096), .I2 (I9985));
ND2X1 gate8272(.O (g3899), .I1 (I7479), .I2 (I7480));
ND2X1 gate8273(.O (I9547), .I1 (g1952), .I2 (g4307));
ND2X1 gate8274(.O (I7179), .I1 (g2351), .I2 (g795));
ND2X1 gate8275(.O (I8326), .I1 (g2011), .I2 (g2721));
ND2X1 gate8276(.O (I12181), .I1 (g6163), .I2 (I12179));
ND2X1 gate8277(.O (I10011), .I1 (g4821), .I2 (I10009));
ND2X1 gate8278(.O (I7611), .I1 (g3771), .I2 (I7609));
ND2X1 gate8279(.O (I10627), .I1 (g1514), .I2 (I10625));
ND2X1 gate8280(.O (g4887), .I1 (I9234), .I2 (I9235));
ND2X1 gate8281(.O (g4228), .I1 (g1408), .I2 (g2665));
ND2X1 gate8282(.O (I10925), .I1 (g2752), .I2 (I10923));
ND2X1 gate8283(.O (I6998), .I1 (g2242), .I2 (I6996));
ND2X1 gate8284(.O (I8327), .I1 (g2011), .I2 (I8326));
ND2X1 gate8285(.O (g6023), .I1 (I10626), .I2 (I10627));
ND2X1 gate8286(.O (I7511), .I1 (g2992), .I2 (I7510));
ND2X1 gate8287(.O (g2333), .I1 (g985), .I2 (g990));
ND2X1 gate8288(.O (I8472), .I1 (g2821), .I2 (I8470));
ND2X1 gate8289(.O (I7574), .I1 (g2999), .I2 (g1718));
ND2X1 gate8290(.O (g9190), .I1 (I15849), .I2 (I15850));
ND2X1 gate8291(.O (I12870), .I1 (g2536), .I2 (I12869));
ND2X1 gate8292(.O (I6925), .I1 (g33), .I2 (I6923));
ND2X1 gate8293(.O (I13395), .I1 (g7212), .I2 (g1057));
ND2X1 gate8294(.O (g5540), .I1 (I9954), .I2 (I9955));
ND2X1 gate8295(.O (I10626), .I1 (g5314), .I2 (I10625));
ND2X1 gate8296(.O (I14245), .I1 (g7683), .I2 (I14244));
ND2X1 gate8297(.O (I10299), .I1 (g5461), .I2 (I10298));
ND2X1 gate8298(.O (g3895), .I1 (I7467), .I2 (I7468));
ND2X1 gate8299(.O (I10298), .I1 (g5461), .I2 (g2562));
ND2X1 gate8300(.O (g6472), .I1 (g5971), .I2 (g5269));
ND2X1 gate8301(.O (I6906), .I1 (g1838), .I2 (I6904));
ND2X1 gate8302(.O (I5599), .I1 (g1481), .I2 (I5598));
ND2X1 gate8303(.O (I9194), .I1 (g4252), .I2 (g1652));
ND2X1 gate8304(.O (I10856), .I1 (g2584), .I2 (I10854));
ND2X1 gate8305(.O (I15882), .I1 (g9179), .I2 (I15880));
ND2X1 gate8306(.O (I7139), .I1 (g2404), .I2 (I7138));
ND2X1 gate8307(.O (I9071), .I1 (g1149), .I2 (I9069));
ND2X1 gate8308(.O (I9242), .I1 (g2540), .I2 (I9241));
ND3X1 gate8309(.O (g5291), .I1 (g4344), .I2 (g5002), .I3 (g4963));
ND2X1 gate8310(.O (I9948), .I1 (g4905), .I2 (I9946));
ND2X1 gate8311(.O (I8581), .I1 (g2498), .I2 (g2777));
ND2X1 gate8312(.O (I9955), .I1 (g4831), .I2 (I9953));
ND2X1 gate8313(.O (g2751), .I1 (I6500), .I2 (I6501));
ND2X1 gate8314(.O (I6876), .I1 (g1967), .I2 (g1910));
ND2X1 gate8315(.O (I9769), .I1 (g1114), .I2 (I9767));
ND2X1 gate8316(.O (I10080), .I1 (g2256), .I2 (I10078));
ND2X1 gate8317(.O (I10924), .I1 (g5525), .I2 (I10923));
ND2X1 gate8318(.O (I15849), .I1 (g9162), .I2 (I15848));
ND2X1 gate8319(.O (g3286), .I1 (I6905), .I2 (I6906));
ND2X1 gate8320(.O (I15848), .I1 (g9162), .I2 (g9154));
ND2X1 gate8321(.O (I9993), .I1 (g2145), .I2 (I9992));
ND2X1 gate8322(.O (I12597), .I1 (g6582), .I2 (I12596));
ND2X1 gate8323(.O (I5695), .I1 (g1513), .I2 (g1524));
ND2X1 gate8324(.O (I7444), .I1 (g2973), .I2 (I7443));
ND2X1 gate8325(.O (I7269), .I1 (g2486), .I2 (I7268));
ND2X1 gate8326(.O (I10198), .I1 (g1958), .I2 (I10196));
ND2X1 gate8327(.O (g5594), .I1 (I10072), .I2 (I10073));
ND2X1 gate8328(.O (I13785), .I1 (g7427), .I2 (g1477));
ND2X1 gate8329(.O (I6877), .I1 (g1967), .I2 (I6876));
ND2X1 gate8330(.O (I10868), .I1 (g2605), .I2 (I10866));
ND2X1 gate8331(.O (g2474), .I1 (g1405), .I2 (g1412));
ND2X1 gate8332(.O (I12854), .I1 (g6695), .I2 (I12852));
ND2X1 gate8333(.O (I10225), .I1 (g4895), .I2 (I10223));
ND2X1 gate8334(.O (I11151), .I1 (g3038), .I2 (I11149));
ND2X1 gate8335(.O (I11172), .I1 (g3038), .I2 (I11170));
ND2X1 gate8336(.O (I6064), .I1 (g852), .I2 (g883));
ND2X1 gate8337(.O (g4893), .I1 (g2460), .I2 (g4312));
ND2X1 gate8338(.O (g5550), .I1 (g1879), .I2 (g4830));
ND2X1 gate8339(.O (I14244), .I1 (g7683), .I2 (g1065));
ND2X1 gate8340(.O (g3900), .I1 (I7486), .I2 (I7487));
ND2X1 gate8341(.O (g6163), .I1 (g5633), .I2 (g3716));
ND2X1 gate8342(.O (I7436), .I1 (g2517), .I2 (g3822));
ND2X1 gate8343(.O (I12550), .I1 (g6689), .I2 (g1462));
ND2X1 gate8344(.O (g4821), .I1 (g4220), .I2 (g3605));
ND2X1 gate8345(.O (I6844), .I1 (g2016), .I2 (I6842));
ND2X1 gate8346(.O (I12596), .I1 (g6582), .I2 (g1126));
ND2X1 gate8347(.O (I7422), .I1 (g2525), .I2 (I7421));
ND2X1 gate8348(.O (I13377), .I1 (g7199), .I2 (I13376));
ND2X1 gate8349(.O (I12180), .I1 (g1961), .I2 (I12179));
ND2X1 gate8350(.O (I10010), .I1 (g1949), .I2 (I10009));
ND2X1 gate8351(.O (g3886), .I1 (I7422), .I2 (I7423));
ND2X1 gate8352(.O (I6814), .I1 (g210), .I2 (I6813));
ND2X1 gate8353(.O (I10079), .I1 (g4911), .I2 (I10078));
ND2X1 gate8354(.O (I7437), .I1 (g2517), .I2 (I7436));
ND2X1 gate8355(.O (g3314), .I1 (I6917), .I2 (I6918));
ND2X1 gate8356(.O (I10078), .I1 (g4911), .I2 (g2256));
ND3X1 gate8357(.O (g5312), .I1 (g5009), .I2 (g5002), .I3 (g4963));
ND2X1 gate8358(.O (I10322), .I1 (g2573), .I2 (I10320));
ND2X1 gate8359(.O (g2051), .I1 (g1444), .I2 (g1450));
ND2X1 gate8360(.O (I10901), .I1 (g2752), .I2 (I10899));
ND2X1 gate8361(.O (I6918), .I1 (g1732), .I2 (I6916));
ND2X1 gate8362(.O (I9980), .I1 (g2092), .I2 (I9978));
ND2X1 gate8363(.O (I9069), .I1 (g4400), .I2 (g1149));
ND2X1 gate8364(.O (I8583), .I1 (g2777), .I2 (I8581));
ND2X1 gate8365(.O (g4359), .I1 (I8327), .I2 (I8328));
ND2X1 gate8366(.O (I10144), .I1 (g1916), .I2 (I10142));
ND2X1 gate8367(.O (I11551), .I1 (g1045), .I2 (I11549));
ND2X1 gate8368(.O (g3887), .I1 (I7429), .I2 (I7430));
ND2X1 gate8369(.O (I7454), .I1 (g1106), .I2 (I7452));
ND2X1 gate8370(.O (I10336), .I1 (g2573), .I2 (I10334));
ND2X1 gate8371(.O (g6627), .I1 (I11874), .I2 (I11875));
ND2X1 gate8372(.O (I7532), .I1 (g2487), .I2 (I7531));
ND2X1 gate8373(.O (I10017), .I1 (g4700), .I2 (g2174));
ND2X1 gate8374(.O (I5619), .I1 (g1092), .I2 (g1130));
ND2X1 gate8375(.O (I13376), .I1 (g7199), .I2 (g1472));
ND2X1 gate8376(.O (I11103), .I1 (g2712), .I2 (I11101));
ND2X1 gate8377(.O (I11095), .I1 (g5515), .I2 (I11094));
ND2X1 gate8378(.O (g8633), .I1 (g8176), .I2 (g6232));
ND2X1 gate8379(.O (I8503), .I1 (g2986), .I2 (I8502));
ND2X1 gate8380(.O (g4880), .I1 (g4287), .I2 (g1879));
ND3X1 gate8381(.O (g5576), .I1 (g4894), .I2 (g4888), .I3 (g4884));
ND2X1 gate8382(.O (I10224), .I1 (g2522), .I2 (I10223));
ND2X1 gate8383(.O (I7429), .I1 (g3222), .I2 (I7428));
ND2X1 gate8384(.O (I8120), .I1 (g1904), .I2 (I8119));
ND2X1 gate8385(.O (I12015), .I1 (g5874), .I2 (g5847));
ND2X1 gate8386(.O (I5598), .I1 (g1481), .I2 (g1489));
ND2X1 gate8387(.O (g6276), .I1 (I11116), .I2 (I11117));
ND2X1 gate8388(.O (g4243), .I1 (I8165), .I2 (I8166));
ND2X1 gate8389(.O (g5747), .I1 (I10299), .I2 (I10300));
ND2X1 gate8390(.O (I6842), .I1 (g205), .I2 (g2016));
ND2X1 gate8391(.O (I7138), .I1 (g2404), .I2 (g2397));
ND2X1 gate8392(.O (I10954), .I1 (g2340), .I2 (I10952));
ND2X1 gate8393(.O (I6941), .I1 (g2051), .I2 (I6939));
ND2X1 gate8394(.O (g6503), .I1 (g5269), .I2 (g5897));
ND2X1 gate8395(.O (I5519), .I1 (g1087), .I2 (g1098));
ND2X1 gate8396(.O (I12179), .I1 (g1961), .I2 (g6163));
ND2X1 gate8397(.O (g8681), .I1 (I14838), .I2 (I14839));
ND2X1 gate8398(.O (I15899), .I1 (g9203), .I2 (I15897));
ND2X1 gate8399(.O (I15898), .I1 (g9202), .I2 (I15897));
ND2X1 gate8400(.O (I12953), .I1 (g1467), .I2 (I12951));
ND2X1 gate8401(.O (I8244), .I1 (g2011), .I2 (I8243));
ND2X1 gate8402(.O (g6277), .I1 (I11123), .I2 (I11124));
ND2X1 gate8403(.O (I7575), .I1 (g2999), .I2 (I7574));
ND2X1 gate8404(.O (I8340), .I1 (g1698), .I2 (I8338));
ND2X1 gate8405(.O (g4090), .I1 (I7892), .I2 (I7893));
ND2X1 gate8406(.O (I9768), .I1 (g4832), .I2 (I9767));
ND2X1 gate8407(.O (g6516), .I1 (g5897), .I2 (g5278));
ND2X1 gate8408(.O (g3129), .I1 (I6843), .I2 (I6844));
ND2X1 gate8409(.O (g4456), .I1 (I8471), .I2 (I8472));
ND2X1 gate8410(.O (I7539), .I1 (g2996), .I2 (I7538));
ND2X1 gate8411(.O (g2995), .I1 (I6740), .I2 (I6741));
ND2X1 gate8412(.O (g2294), .I1 (I6065), .I2 (I6066));
ND2X1 gate8413(.O (g3221), .I1 (I6877), .I2 (I6878));
ND2X1 gate8414(.O (I7268), .I1 (g2486), .I2 (g955));
ND2X1 gate8415(.O (I5506), .I1 (g1532), .I2 (I5505));
ND2X1 gate8416(.O (I7452), .I1 (g3226), .I2 (g1106));
ND2X1 gate8417(.O (g6709), .I1 (I12052), .I2 (I12053));
ND2X1 gate8418(.O (I6540), .I1 (g2557), .I2 (I6538));
ND2X1 gate8419(.O (I10093), .I1 (g4881), .I2 (I10092));
ND2X1 gate8420(.O (I9195), .I1 (g4252), .I2 (I9194));
ND2X1 gate8421(.O (I7086), .I1 (g1753), .I2 (I7085));
ND2X1 gate8422(.O (I7486), .I1 (g2989), .I2 (I7485));
ND2X1 gate8423(.O (g6435), .I1 (I11575), .I2 (I11576));
ND2X1 gate8424(.O (g6482), .I1 (g5269), .I2 (g5847));
ND2X1 gate8425(.O (I7504), .I1 (g2498), .I2 (I7503));
ND2X1 gate8426(.O (I10875), .I1 (g2595), .I2 (I10873));
ND2X1 gate8427(.O (I7070), .I1 (g1643), .I2 (I7068));
ND2X1 gate8428(.O (I14837), .I1 (g8660), .I2 (g1073));
ND2X1 gate8429(.O (g4686), .I1 (I8956), .I2 (I8957));
ND2X1 gate8430(.O (I11094), .I1 (g5515), .I2 (g2734));
ND2X1 gate8431(.O (I5507), .I1 (g1528), .I2 (I5505));
ND2X1 gate8432(.O (I11150), .I1 (g5473), .I2 (I11149));
ND2X1 gate8433(.O (I13801), .I1 (g7429), .I2 (I13800));
ND2X1 gate8434(.O (I9692), .I1 (g5096), .I2 (I9691));
ND2X1 gate8435(.O (g7444), .I1 (I13588), .I2 (I13589));
ND2X1 gate8436(.O (I13018), .I1 (g1142), .I2 (I13016));
ND2X1 gate8437(.O (I6259), .I1 (g901), .I2 (I6257));
ND2X1 gate8438(.O (I7087), .I1 (g1918), .I2 (I7085));
ND2X1 gate8439(.O (I7487), .I1 (g1708), .I2 (I7485));
ND2X1 gate8440(.O (I6923), .I1 (g1728), .I2 (g33));
ND2X1 gate8441(.O (g3818), .I1 (I7278), .I2 (I7279));
ND2X1 gate8442(.O (I8394), .I1 (g1925), .I2 (I8392));
ND2X1 gate8443(.O (I9979), .I1 (g4880), .I2 (I9978));
ND2X1 gate8444(.O (g3893), .I1 (I7453), .I2 (I7454));
ND2X1 gate8445(.O (I7445), .I1 (g1701), .I2 (I7443));
ND2X1 gate8446(.O (I7173), .I1 (g1739), .I2 (I7172));
ND2X1 gate8447(.O (I8471), .I1 (g2525), .I2 (I8470));
ND2X1 gate8448(.O (I9828), .I1 (g1509), .I2 (I9826));
ND2X1 gate8449(.O (g5595), .I1 (I10079), .I2 (I10080));
ND2X1 gate8450(.O (I8955), .I1 (g4246), .I2 (g1110));
ND2X1 gate8451(.O (g9192), .I1 (I15863), .I2 (I15864));
ND2X1 gate8452(.O (I8254), .I1 (g2454), .I2 (I8253));
ND2X1 gate8453(.O (I10836), .I1 (g2584), .I2 (I10834));
ND2X1 gate8454(.O (I9746), .I1 (g4826), .I2 (I9745));
ND2X1 gate8455(.O (I7459), .I1 (g2506), .I2 (g3815));
ND2X1 gate8456(.O (I11102), .I1 (g5491), .I2 (I11101));
ND2X1 gate8457(.O (I11157), .I1 (g5482), .I2 (I11156));
ND2X1 gate8458(.O (g3939), .I1 (I7617), .I2 (I7618));
ND2X1 gate8459(.O (I8150), .I1 (g3229), .I2 (g38));
ND2X1 gate8460(.O (g3083), .I1 (I6814), .I2 (I6815));
ND2X1 gate8461(.O (I9953), .I1 (g2131), .I2 (g4831));
ND4X1 gate8462(.O (g4879), .I1 (g2595), .I2 (g2584), .I3 (g4270), .I4 (g4281));
ND2X1 gate8463(.O (I10313), .I1 (g5484), .I2 (g1041));
ND2X1 gate8464(.O (I6065), .I1 (g852), .I2 (I6064));
ND2X1 gate8465(.O (I10305), .I1 (g5470), .I2 (g3019));
ND2X1 gate8466(.O (I10900), .I1 (g5520), .I2 (I10899));
ND2X1 gate8467(.O (I9747), .I1 (g1549), .I2 (I9745));
ND2X1 gate8468(.O (g8627), .I1 (g6232), .I2 (g8091));
ND2X1 gate8469(.O (I11550), .I1 (g5984), .I2 (I11549));
ND2X1 gate8470(.O (I9241), .I1 (g2540), .I2 (g4305));
ND2X1 gate8471(.O (g5512), .I1 (g1879), .I2 (g4877));
ND2X1 gate8472(.O (I7188), .I1 (g1834), .I2 (I7186));
ND2X1 gate8473(.O (I10874), .I1 (g5516), .I2 (I10873));
ND2X1 gate8474(.O (I7216), .I1 (g2091), .I2 (I7214));
ND2X1 gate8475(.O (I12952), .I1 (g7003), .I2 (I12951));
ND2X1 gate8476(.O (I7428), .I1 (g3222), .I2 (g1541));
ND2X1 gate8477(.O (I10009), .I1 (g1949), .I2 (g4821));
ND2X1 gate8478(.O (I7430), .I1 (g1541), .I2 (I7428));
ND2X1 gate8479(.O (I11156), .I1 (g5482), .I2 (g3052));
ND2X1 gate8480(.O (I9152), .I1 (g3883), .I2 (I9151));
ND2X1 gate8481(.O (I5621), .I1 (g1130), .I2 (I5619));
ND2X1 gate8482(.O (I6815), .I1 (g2052), .I2 (I6813));
ND2X1 gate8483(.O (g4905), .I1 (g4282), .I2 (g3533));
ND2X1 gate8484(.O (g3811), .I1 (I7269), .I2 (I7270));
ND2X1 gate8485(.O (g3315), .I1 (I6924), .I2 (I6925));
ND2X1 gate8486(.O (I10907), .I1 (g5492), .I2 (I10906));
ND2X1 gate8487(.O (I7609), .I1 (g2471), .I2 (g3771));
ND2X1 gate8488(.O (I12834), .I1 (g6709), .I2 (I12832));
ND2X1 gate8489(.O (I8392), .I1 (g2949), .I2 (g1925));
ND2X1 gate8490(.O (I9170), .I1 (g1935), .I2 (I9169));
ND2X1 gate8491(.O (I15889), .I1 (g9191), .I2 (I15887));
NR4X1 gate8492(.O (g4884), .I1 (g4492), .I2 (g4476), .I3 (g4456), .I4 (g4294));
NR3X1 gate8493(.O (g8656), .I1 (g8199), .I2 (I14758), .I3 (I14759));
NR2X1 gate8494(.O (g3260), .I1 (g1728), .I2 (g2490));
NR2X1 gate8495(.O (g5615), .I1 (g4714), .I2 (g3002));
NR3X1 gate8496(.O (g8236), .I1 (g8199), .I2 (I14495), .I3 (I14496));
NR2X1 gate8497(.O (g4160), .I1 (g1231), .I2 (g2834));
NR2X1 gate8498(.O (g7406), .I1 (g7191), .I2 (g1600));
NR2X1 gate8499(.O (g6259), .I1 (g3002), .I2 (g5312));
NR4X1 gate8500(.O (g6465), .I1 (g5403), .I2 (g5802), .I3 (g5769), .I4 (g5790));
NR4X1 gate8501(.O (g3515), .I1 (g1388), .I2 (g2262), .I3 (g2230), .I4 (g2214));
NR3X1 gate8502(.O (g8812), .I1 (g8443), .I2 (g8421), .I3 (I15086));
NR2X1 gate8503(.O (g3528), .I1 (g2343), .I2 (g1391));
NR2X1 gate8504(.O (g8073), .I1 (g7658), .I2 (g7654));
NR2X1 gate8505(.O (g3555), .I1 (g2359), .I2 (g1398));
NR3X1 gate8506(.O (g8819), .I1 (g8443), .I2 (g8421), .I3 (I15113));
NR3X1 gate8507(.O (g8694), .I1 (g7658), .I2 (g8613), .I3 (g7634));
NR3X1 gate8508(.O (g8806), .I1 (g8443), .I2 (g8421), .I3 (I15044));
NR3X1 gate8509(.O (g8230), .I1 (g8199), .I2 (I14467), .I3 (I14468));
NR3X1 gate8510(.O (g8807), .I1 (g8443), .I2 (g8421), .I3 (I15055));
NR4X1 gate8511(.O (g4888), .I1 (g4548), .I2 (g4528), .I3 (g4513), .I4 (g4502));
NR3X1 gate8512(.O (g8859), .I1 (g8493), .I2 (g8239), .I3 (I15165));
NR2X1 gate8513(.O (g7326), .I1 (g7194), .I2 (g6999));
NR3X1 gate8514(.O (g8699), .I1 (g7658), .I2 (g8613), .I3 (g7634));
NR3X1 gate8515(.O (g8855), .I1 (g7658), .I2 (g8613), .I3 (g7634));
NR2X1 gate8516(.O (g8644), .I1 (g4146), .I2 (g8128));
NR2X1 gate8517(.O (g6193), .I1 (g1926), .I2 (g5310));
NR3X1 gate8518(.O (g8818), .I1 (g8443), .I2 (g8421), .I3 (I15102));
NR2X1 gate8519(.O (g3885), .I1 (g3310), .I2 (g3466));
NR2X1 gate8520(.O (g6174), .I1 (g1855), .I2 (g5305));
NR2X1 gate8521(.O (g3233), .I1 (g1714), .I2 (g1459));
NR3X1 gate8522(.O (g8811), .I1 (g8443), .I2 (g8421), .I3 (I15075));
NR2X1 gate8523(.O (g8629), .I1 (g6270), .I2 (g8009));
NR4X1 gate8524(.O (g8279), .I1 (g7658), .I2 (g7616), .I3 (g8082), .I4 (g7634));
NR4X1 gate8525(.O (g3504), .I1 (g1375), .I2 (g2229), .I3 (g2213), .I4 (g2206));
NR4X1 gate8526(.O (g8625), .I1 (g1000), .I2 (g6573), .I3 (g1860), .I4 (g8009));
NR3X1 gate8527(.O (g8232), .I1 (g8199), .I2 (I14479), .I3 (I14480));
NR3X1 gate8528(.O (g8659), .I1 (g8199), .I2 (I14771), .I3 (I14772));
NR2X1 gate8529(.O (g6209), .I1 (g2332), .I2 (g5305));
NR4X1 gate8530(.O (g8630), .I1 (g6110), .I2 (g7784), .I3 (g3591), .I4 (g1864));
NR2X1 gate8531(.O (g6184), .I1 (g875), .I2 (g5291));
NR3X1 gate8532(.O (g8655), .I1 (g8199), .I2 (I14753), .I3 (I14754));
NR2X1 gate8533(.O (g5772), .I1 (g5428), .I2 (g1888));
NR2X1 gate8534(.O (g2521), .I1 (g65), .I2 (g62));
NR2X1 gate8535(.O (g7324), .I1 (g7189), .I2 (g6994));
NR4X1 gate8536(.O (g5023), .I1 (g3894), .I2 (g3889), .I3 (g3886), .I4 (g4359));
NR4X1 gate8537(.O (g8360), .I1 (g7658), .I2 (g7616), .I3 (g8082), .I4 (g7634));
NR4X1 gate8538(.O (g8641), .I1 (g6559), .I2 (g162), .I3 (g7784), .I4 (g3591));
NR2X1 gate8539(.O (g3505), .I1 (g2263), .I2 (g1395));
NR3X1 gate8540(.O (g8658), .I1 (g8199), .I2 (I14766), .I3 (I14767));
NR3X1 gate8541(.O (g8680), .I1 (g8493), .I2 (g8239), .I3 (I14834));
NR3X1 gate8542(.O (g4894), .I1 (g4298), .I2 (g4575), .I3 (g4563));
NR2X1 gate8543(.O (g7314), .I1 (g7180), .I2 (g6972));
NR4X1 gate8544(.O (g8092), .I1 (g7634), .I2 (g7628), .I3 (g7616), .I4 (g7611));
NR2X1 gate8545(.O (g7322), .I1 (g7188), .I2 (g6991));
NR4X1 gate8546(.O (g8523), .I1 (g7658), .I2 (g7616), .I3 (g8082), .I4 (g7634));
NR2X1 gate8547(.O (g7312), .I1 (g7178), .I2 (g6970));
NR2X1 gate8548(.O (g6452), .I1 (g6270), .I2 (g2245));
NR2X1 gate8549(.O (g2014), .I1 (g1421), .I2 (g1416));
NR3X1 gate8550(.O (g8862), .I1 (g8493), .I2 (g8239), .I3 (I15172));
NR2X1 gate8551(.O (g6185), .I1 (g5305), .I2 (g1590));
NR3X1 gate8552(.O (g8679), .I1 (g8493), .I2 (g8239), .I3 (I14831));
NR4X1 gate8553(.O (g5039), .I1 (g3924), .I2 (g3914), .I3 (g3906), .I4 (g3899));
NR3X1 gate8554(.O (g8805), .I1 (g8443), .I2 (g8421), .I3 (I15033));
NR3X1 gate8555(.O (g7152), .I1 (g6253), .I2 (g7083), .I3 (g5418));
NR3X1 gate8556(.O (g6664), .I1 (g5836), .I2 (g1901), .I3 (g1788));
NR2X1 gate8557(.O (g1980), .I1 (g1430), .I2 (g1431));
NR3X1 gate8558(.O (g8233), .I1 (g8199), .I2 (I14484), .I3 (I14485));
NR3X1 gate8559(.O (g8706), .I1 (g7658), .I2 (g8613), .I3 (g7634));
NR4X1 gate8560(.O (g6910), .I1 (g1011), .I2 (g1837), .I3 (g6559), .I4 (g1008));
NR3X1 gate8561(.O (g8707), .I1 (g7658), .I2 (g8613), .I3 (g7634));
NR2X1 gate8562(.O (g7328), .I1 (g7196), .I2 (g7001));
NR2X1 gate8563(.O (g3516), .I1 (g2282), .I2 (g1401));
NR4X1 gate8564(.O (g6197), .I1 (g875), .I2 (g866), .I3 (g1590), .I4 (g5291));
NR2X1 gate8565(.O (g8635), .I1 (g1034), .I2 (g8128));
NR2X1 gate8566(.O (g8801), .I1 (g8635), .I2 (g3790));
NR2X1 gate8567(.O (g3310), .I1 (g936), .I2 (g2557));
NR2X1 gate8568(.O (g7318), .I1 (g7185), .I2 (g6979));
NR2X1 gate8569(.O (g7321), .I1 (g7187), .I2 (g6990));
NR3X1 gate8570(.O (g3237), .I1 (g1444), .I2 (g1838), .I3 (g1454));
NR3X1 gate8571(.O (g8861), .I1 (g8493), .I2 (g8239), .I3 (I15169));
NR2X1 gate8572(.O (g4354), .I1 (g1424), .I2 (g3541));
NR3X1 gate8573(.O (g8803), .I1 (g8443), .I2 (g8421), .I3 (I15021));
NR2X1 gate8574(.O (g4676), .I1 (g3885), .I2 (g3094));
NR3X1 gate8575(.O (g8847), .I1 (g8493), .I2 (g8239), .I3 (I15147));
NR2X1 gate8576(.O (g4349), .I1 (g2496), .I2 (g3310));
NR3X1 gate8577(.O (g3225), .I1 (g1021), .I2 (g1025), .I3 (g1889));
NR2X1 gate8578(.O (g7566), .I1 (g7421), .I2 (g1597));
NR3X1 gate8579(.O (g8863), .I1 (g8493), .I2 (g8239), .I3 (I15175));
NR2X1 gate8580(.O (g1964), .I1 (g1428), .I2 (g1429));
NR3X1 gate8581(.O (g7209), .I1 (g1789), .I2 (g146), .I3 (g6984));
NR3X1 gate8582(.O (g5614), .I1 (g3002), .I2 (g1590), .I3 (g4714));
NR2X1 gate8583(.O (g4318), .I1 (g3681), .I2 (g1590));
NR2X1 gate8584(.O (g6214), .I1 (g878), .I2 (g5284));
NR2X1 gate8585(.O (g4232), .I1 (g1934), .I2 (g3591));
NR3X1 gate8586(.O (g6489), .I1 (g5802), .I2 (g5769), .I3 (g5790));
NR3X1 gate8587(.O (g3790), .I1 (g985), .I2 (g990), .I3 (g2295));
NR3X1 gate8588(.O (g5056), .I1 (g3556), .I2 (g2872), .I3 (g3938));
NR3X1 gate8589(.O (g8850), .I1 (g8493), .I2 (g8239), .I3 (I15152));
endmodule