module s38584(clk, g35, g36, g6744, g6745, g6746, g6747, g6748, g6749, g6750, g6751, g6752, g6753, g84, g120, g5, g113, g126, g99, g53, g116, g92, g56, g91, g44, g57, g100, g54, g124, g125, g114, g134, g72, g115, g135, g90, g127, g64, g73, g7243, g7245, g7257, g7260, g7540, g7916, g7946, g8132, g8178, g8215, g8235, g8277, g8279, g8283, g8291, g8342, g8344, g8353, g8358, g8398, g8403, g8416, g8475, g8719, g8783, g8784, g8785, g8786, g8787, g8788, g8789, g8839, g8870, g8915, g8916, g8917, g8918, g8919, g8920, g9019, g9048, g9251, g9497, g9553, g9555, g9615, g9617, g9680, g9682, g9741, g9743, g9817, g10122, g10306, g10500, g10527, g11349, g11388, g11418, g11447, g11678, g11770, g12184, g12238, g12300, g12350, g12368, g12422, g12470, g12832, g12919, g12923, g13039, g13049, g13068, g13085, g13099, g13259, g13272, g13865, g13881, g13895, g13906, g13926, g13966, g14096, g14125, g14147, g14167, g14189, g14201, g14217, g14421, g14451, g14518, g14597, g14635, g14662, g14673, g14694, g14705, g14738, g14749, g14779, g14828, g16603, g16624, g16627, g16656, g16659, g16686, g16693, g16718, g16722, g16744, g16748, g16775, g16874, g16924, g16955, g17291, g17316, g17320, g17400, g17404, g17423, g17519, g17577, g17580, g17604, g17607, g17639, g17646, g17649, g17674, g17678, g17685, g17688, g17711, g17715, g17722, g17739, g17743, g17760, g17764, g17778, g17787, g17813, g17819, g17845, g17871, g18092, g18094, g18095, g18096, g18097, g18098, g18099, g18100, g18101, g18881, g19334, g19357, g20049, g20557, g20652, g20654, g20763, g20899, g20901, g21176, g21245, g21270, g21292, g21698, g21727, g23002, g23190, g23612, g23652, g23683, g23759, g24151, g25114, g25167, g25219, g25259, g25582, g25583, g25584, g25585, g25586, g25587, g25588, g25589, g25590, g26801, g26875, g26876, g26877, g27831, g28030, g28041, g28042, g28753, g29210, g29211, g29212, g29213, g29214, g29215, g29216, g29217, g29218, g29219, g29220, g29221, g30327, g30329, g30330, g30331, g30332, g31521, g31656, g31665, g31793, g31860, g31861, g31862, g31863, g32185, g32429, g32454, g32975, g33079, g33435, g33533, g33636, g33659, g33874, g33894, g33935, g33945, g33946, g33947, g33948, g33949, g33950, g33959, g34201, g34221, g34232, g34233, g34234, g34235, g34236, g34237, g34238, g34239, g34240, g34383, g34425, g34435, g34436, g34437, g34597, g34788, g34839, g34913, g34915, g34917, g34919, g34921, g34923, g34925, g34927, g34956, g34972, g24168, g24178, g12833, g24174, g24181, g24172, g24161, g24177, g24171, g24163, g24170, g24185, g24164, g24173, g24162, g24179, g24180, g24175, g24183, g24166, g24176, g24184, g24169, g24182, g24165, g24167);
input clk, g35, g36, g6744, g6745, g6746, g6747, g6748, g6749, g6750, g6751, g6752, g6753, g84, g120, g5, g113, g126, g99, g53, g116, g92, g56, g91, g44, g57, g100, g54, g124, g125, g114, g134, g72, g115, g135, g90, g127, g64, g73;
output g7243, g7245, g7257, g7260, g7540, g7916, g7946, g8132, g8178, g8215, g8235, g8277, g8279, g8283, g8291, g8342, g8344, g8353, g8358, g8398, g8403, g8416, g8475, g8719, g8783, g8784, g8785, g8786, g8787, g8788, g8789, g8839, g8870, g8915, g8916, g8917, g8918, g8919, g8920, g9019, g9048, g9251, g9497, g9553, g9555, g9615, g9617, g9680, g9682, g9741, g9743, g9817, g10122, g10306, g10500, g10527, g11349, g11388, g11418, g11447, g11678, g11770, g12184, g12238, g12300, g12350, g12368, g12422, g12470, g12832, g12919, g12923, g13039, g13049, g13068, g13085, g13099, g13259, g13272, g13865, g13881, g13895, g13906, g13926, g13966, g14096, g14125, g14147, g14167, g14189, g14201, g14217, g14421, g14451, g14518, g14597, g14635, g14662, g14673, g14694, g14705, g14738, g14749, g14779, g14828, g16603, g16624, g16627, g16656, g16659, g16686, g16693, g16718, g16722, g16744, g16748, g16775, g16874, g16924, g16955, g17291, g17316, g17320, g17400, g17404, g17423, g17519, g17577, g17580, g17604, g17607, g17639, g17646, g17649, g17674, g17678, g17685, g17688, g17711, g17715, g17722, g17739, g17743, g17760, g17764, g17778, g17787, g17813, g17819, g17845, g17871, g18092, g18094, g18095, g18096, g18097, g18098, g18099, g18100, g18101, g18881, g19334, g19357, g20049, g20557, g20652, g20654, g20763, g20899, g20901, g21176, g21245, g21270, g21292, g21698, g21727, g23002, g23190, g23612, g23652, g23683, g23759, g24151, g25114, g25167, g25219, g25259, g25582, g25583, g25584, g25585, g25586, g25587, g25588, g25589, g25590, g26801, g26875, g26876, g26877, g27831, g28030, g28041, g28042, g28753, g29210, g29211, g29212, g29213, g29214, g29215, g29216, g29217, g29218, g29219, g29220, g29221, g30327, g30329, g30330, g30331, g30332, g31521, g31656, g31665, g31793, g31860, g31861, g31862, g31863, g32185, g32429, g32454, g32975, g33079, g33435, g33533, g33636, g33659, g33874, g33894, g33935, g33945, g33946, g33947, g33948, g33949, g33950, g33959, g34201, g34221, g34232, g34233, g34234, g34235, g34236, g34237, g34238, g34239, g34240, g34383, g34425, g34435, g34436, g34437, g34597, g34788, g34839, g34913, g34915, g34917, g34919, g34921, g34923, g34925, g34927, g34956, g34972, g24168, g24178, g12833, g24174, g24181, g24172, g24161, g24177, g24171, g24163, g24170, g24185, g24164, g24173, g24162, g24179, g24180, g24175, g24183, g24166, g24176, g24184, g24169, g24182, g24165, g24167;
wire clk, g35, g36, g6744, g6745, g6746, g6747, g6748, g6749, g6750, g6751, g6752, g6753, g84, g120, g5, g113, g126, g99, g53, g116, g92, g56, g91, g44, g57, g100, g54, g124, g125, g114, g134, g72, g115, g135, g90, g127, g64, g73;
wire g5057, g2771, g1882, g6462, g2299, g4040, g2547, g559, g3017, g3243, g452;
wire g464, g3542, g5232, g5813, g2907, g1744, g5909, g1802, g3554, g6219, g807;
wire g6031, g847, g976, g4172, g4372, g3512, g749, g3490, g6005, g4235, g1600;
wire g1714, g3649, g3155, g3355, g2236, g4555, g3698, g6073, g1736, g1968, g4621;
wire g5607, g2657, g5659, g490, g311, g6069, g772, g5587, g6177, g6377, g3167;
wire g5615, g4567, g3057, g3457, g6287, g1500, g2563, g4776, g4593, g6199, g2295;
wire g1384, g1339, g5180, g2844, g1024, g5591, g3598, g4264, g767, g5853, g3321;
wire g2089, g4933, g4521, g5507, g3625, g6291, g294, g5559, g5794, g6144, g3813;
wire g562, g608, g1205, g3909, g6259, g5905, g921, g2955, g203, g6088, g1099;
wire g4878, g5204, g5630, g3606, g1926, g6215, g3586, g291, g4674, g3570, g640;
wire g5969, g1862, g676, g843, g4132, g4332, g4153, g5666, g6336, g622, g3506;
wire g4558, g6065, g6322, g3111, g117, g2837, g939, g278, g4492, g4864, g1036;
wire g128, g1178, g3239, g718, g6195, g1135, g6137, g6395, g3380, g5343, g554;
wire g496, g3853, g5134, g1422, g3794, g2485, g925, g48, g5555, g878, g1798;
wire g4076, g2941, g3905, g763, g6255, g4375, g4871, g4722, g590, g6692, g1632;
wire g5313, g3100, g1495, g6497, g1437, g6154, g1579, g5567, g1752, g1917, g744;
wire g3040, g4737, g4809, g6267, g3440, g3969, g1442, g5965, g4477, g1233, g4643;
wire g5264, g6329, g2610, g5160, g5360, g5933, g1454, g753, g1296, g3151, g2980;
wire g6727, g3530, g4742, g4104, g1532, g4304, g2177, g3010, g52, g4754, g1189;
wire g2287, g4273, g1389, g1706, g5835, g1171, g4269, g2399, g3372, g4983, g5611;
wire g3618, g4572, g3143, g2898, g3343, g3235, g4543, g3566, g4534, g4961, g6398;
wire g4927, g2259, g2819, g4414, g5802, g2852, g417, g681, g437, g351, g5901;
wire g2886, g3494, g5511, g3518, g1604, g4135, g5092, g4831, g4382, g6386, g479;
wire g3965, g4749, g2008, g736, g3933, g222, g3050, g5736, g1052, g58, g5623;
wire g2122, g2465, g6483, g5889, g4495, g365, g4653, g3179, g1728, g2433, g3835;
wire g6187, g4917, g1070, g822, g6027, g914, g5339, g4164, g969, g2807, g5424;
wire g4054, g6191, g5077, g5523, g3680, g6637, g174, g1682, g355, g1087, g1105;
wire g2342, g6307, g3802, g6159, g2255, g2815, g911, g43, g4012, g1748, g5551;
wire g5742, g3558, g5499, g2960, g3901, g4888, g6251, g6315, g1373, g3092, g157;
wire g2783, g4281, g3574, g2112, g1283, g433, g4297, g5983, g1459, g758, g5712;
wire g4138, g4639, g6537, g5543, g1582, g3736, g5961, g6243, g632, g1227, g3889;
wire g3476, g1664, g1246, g6128, g6629, g246, g4049, g4449, g2932, g4575, g4098;
wire g4498, g528, g5436, g16, g3139, g102, g4584, g142, g5335, g5831, g239;
wire g1216, g2848, g5805, g5022, g4019, g1030, g3672, g3231, g6490, g1430, g4452;
wire g2241, g1564, g5798, g6148, g6649, g110, g884, g3742, g225, g4486, g4504;
wire g5873, g5037, g2319, g5495, g4185, g5208, g2152, g5579, g5869, g5719, g1589;
wire g5752, g6279, g5917, g2975, g6167, g3983, g2599, g1448, g881, g3712, g2370;
wire g5164, g1333, g153, g6549, g4087, g4801, g2984, g3961, g5770, g962, g101;
wire g4226, g6625, g51, g1018, g1418, g4045, g1467, g2461, g5706, g457, g2756;
wire g5990, g471, g1256, g5029, g6519, g4169, g1816, g4369, g3436, g5787, g4578;
wire g4459, g3831, g2514, g3288, g2403, g2145, g1700, g513, g2841, g5297, g3805;
wire g2763, g4793, g952, g1263, g1950, g5138, g2307, g5109, g5791, g3798, g4664;
wire g2223, g5808, g6645, g2016, g5759, g3873, g3632, g2315, g2811, g5957, g2047;
wire g3869, g6358, g3719, g5575, g46, g3752, g3917, g4188, g1585, g4388, g6275;
wire g6311, g4216, g1041, g2595, g2537, g136, g4430, g4564, g3454, g4826, g6239;
wire g3770, g232, g5268, g6545, g2417, g1772, g4741, g5052, g5452, g1890, g2629;
wire g572, g2130, g4108, g4308, g475, g990, g31, g3412, g45, g799, g3706;
wire g3990, g5385, g5881, g1992, g3029, g3171, g3787, g812, g832, g5897, g4165;
wire g4571, g3281, g4455, g2902, g333, g168, g2823, g3684, g3639, g5331, g3338;
wire g5406, g3791, g269, g401, g6040, g441, g5105, g3808, g9, g3759, g4467;
wire g3957, g4093, g1760, g6151, g6351, g160, g5445, g5373, g2279, g3498, g586;
wire g869, g2619, g1183, g1608, g4197, g5283, g1779, g2652, g5459, g2193, g2393;
wire g5767, g661, g4950, g5535, g2834, g1361, g3419, g6235, g1146, g2625, g150;
wire g1696, g6555, g859, g3385, g3881, g6621, g3470, g3897, g518, g3025, g538;
wire g2606, g1472, g6113, g542, g5188, g5689, g1116, g405, g5216, g6494, g4669;
wire g5428, g996, g4531, g2860, g4743, g6593, g2710, g215, g4411, g1413, g4474;
wire g5308, g6641, g3045, g6, g1936, g55, g504, g2587, g4480, g2311, g3602;
wire g5571, g3578, g468, g5448, g3767, g5827, g3582, g6271, g4688, g5774, g2380;
wire g5196, g5396, g3227, g2020, g4000, g1079, g6541, g3203, g1668, g4760, g262;
wire g1840, g70, g5467, g460, g6209, g74, g5290, g655, g3502, g2204, g5256;
wire g4608, g794, g4023, g4423, g3689, g5381, g5685, g703, g5421, g862, g3247;
wire g2040, g4999, g4146, g4633, g1157, g5723, g4732, g5101, g5817, g2151, g2351;
wire g2648, g6736, g4944, g4072, g344, g4443, g3466, g4116, g5041, g5441, g4434;
wire g3827, g6500, g5673, g3133, g3333, g979, g4681, g298, g3774, g2667, g3396;
wire g4210, g1894, g2988, g3538, g301, g341, g827, g1075, g6077, g2555, g5011;
wire g199, g6523, g1526, g4601, g854, g1484, g4922, g5080, g5863, g4581, g3021;
wire g2518, g2567, g568, g3263, g6613, g6044, g6444, g2965, g5857, g1616, g890;
wire g5976, g3562, g4294, g1404, g3723, g3817, g93, g4501, g287, g2724, g4704;
wire g22, g2878, g5220, g617, g637, g316, g1277, g6513, g336, g2882, g933;
wire g1906, g305, g8, g3368, g2799, g887, g5327, g4912, g4157, g2541, g2153;
wire g550, g255, g1945, g5240, g1478, g3080, g3863, g1959, g3480, g6653, g6719;
wire g2864, g4894, g5681, g3857, g3976, g499, g5413, g1002, g776, g28, g1236;
wire g4646, g2476, g1657, g2375, g63, g6012, g358, g896, g967, g3423, g283;
wire g3161, g2384, g3361, g6675, g4616, g4561, g2024, g3451, g2795, g613, g4527;
wire g1844, g5937, g4546, g3103, g2523, g3303, g2643, g6109, g1489, g5390, g194;
wire g2551, g5156, g3072, g1242, g47, g3443, g4277, g1955, g6049, g3034, g2273;
wire g6715, g4771, g6098, g3147, g3347, g2269, g191, g2712, g626, g2729, g5357;
wire g4991, g6019, g4709, g6419, g6052, g2927, g4340, g5929, g4907, g3317, g4035;
wire g2946, g918, g4082, g6486, g2036, g577, g1620, g2831, g667, g930, g3937;
wire g5782, g817, g1249, g837, g3668, g599, g5475, g739, g5949, g6682, g6105;
wire g904, g2873, g1854, g5084, g5603, g4222, g2495, g2437, g2102, g2208, g2579;
wire g4064, g4899, g2719, g4785, g5583, g781, g6173, g6373, g2917, g686, g1252;
wire g671, g2265, g6283, g6369, g5276, g6459, g901, g4194, g5527, g4489, g1974;
wire g1270, g4966, g6415, g6227, g3929, g5503, g4242, g5925, g1124, g4955, g5224;
wire g2012, g6203, g5120, g5320, g2389, g4438, g2429, g2787, g1287, g2675, g66;
wire g4836, g1199, g1399, g5547, g3782, g6428, g2138, g3661, g2338, g4229, g6247;
wire g2791, g3949, g1291, g5945, g5244, g2759, g6741, g785, g1259, g3484, g209;
wire g6609, g5517, g2449, g2575, g65, g2715, g936, g2098, g4462, g604, g6589;
wire g1886, g6466, g6365, g6711, g429, g1870, g4249, g6455, g3004, g1825, g6133;
wire g1008, g4392, g5002, g3546, g5236, g1768, g4854, g3925, g6509, g732, g2504;
wire g1322, g4520, g4219, g2185, g37, g4031, g2070, g4812, g6093, g968, g4176;
wire g4005, g4405, g872, g6181, g6381, g4765, g5563, g1395, g1913, g2331, g6263;
wire g50, g3945, g347, g5731, g4473, g1266, g5489, g714, g2748, g5471, g4540;
wire g6723, g6605, g2445, g2173, g4287, g2491, g4849, g2169, g2283, g6585, g121;
wire g2407, g2868, g2767, g1783, g3310, g1312, g5212, g4245, g645, g4291, g79;
wire g182, g1129, g2227, g6058, g4207, g2246, g1830, g3590, g392, g1592, g6505;
wire g6411, g1221, g5921, g106, g146, g218, g6474, g1932, g1624, g5062, g5462;
wire g2689, g6573, g1677, g2028, g2671, g1576, g4408, g34, g1848, g3089, g3731;
wire g86, g5485, g2741, g802, g2638, g4122, g4322, g5941, g2108, g6000, g25;
wire g1644, g595, g2217, g1319, g2066, g1152, g5252, g2165, g2571, g5176, g391;
wire g5005, g2711, g6023, g1211, g2827, g6423, g875, g4859, g424, g1274, g1426;
wire g85, g2803, g6451, g1821, g2509, g5073, g1280, g4815, g6346, g6633, g5124;
wire g1083, g6303, g5069, g2994, g650, g1636, g3921, g2093, g6732, g1306, g5377;
wire g1061, g3462, g2181, g956, g1756, g5849, g4112, g2685, g2197, g6116, g2421;
wire g1046, g482, g4401, g6434, g1514, g329, g6565, g2950, g4129, g1345, g6533;
wire g3298, g3085, g4727, g6697, g1536, g3941, g370, g5694, g1858, g446, g4932;
wire g3219, g1811, g3431, g6601, g3376, g2441, g1874, g4349, g6581, g6597, g5008;
wire g3610, g2890, g1978, g1612, g112, g2856, g6479, g1982, g6668, g5228, g4119;
wire g6390, g1542, g4258, g4818, g5033, g4717, g1554, g3849, g6704, g3199, g5845;
wire g4975, g790, g5913, g1902, g6163, g4125, g4821, g4939, g1056, g3207, g4483;
wire g3259, g5142, g5248, g2126, g3694, g5481, g1964, g5097, g3215, g4027, g111;
wire g4427, g7, g2779, g4200, g4446, g1720, g1367, g5112, g19, g4145, g2161;
wire g376, g2361, g4191, g582, g2051, g1193, g5401, g3408, g2327, g907, g947;
wire g1834, g3594, g2999, g5727, g2303, g6661, g3065, g699, g723, g5703, g546;
wire g2472, g5953, g3096, g6439, g1740, g3550, g3845, g2116, g5677, g3195, g3913;
wire g4537, g1687, g2681, g2533, g324, g2697, g5747, g4417, g6561, g1141, g1570;
wire g2413, g1710, g6527, g6404, g3255, g1691, g2936, g5644, g5152, g5352, g4213;
wire g6120, g2775, g2922, g1111, g5893, g1311, g3267, g6617, g2060, g4512, g5599;
wire g3401, g4366, g3676, g94, g3129, g3329, g5170, g4456, g5821, g6299, g1239;
wire g3727, g2079, g4698, g3703, g1559, g943, g411, g6140, g3953, g3068, g2704;
wire g6035, g6082, g49, g1300, g4057, g5200, g4843, g5046, g2250, g319, g4549;
wire g2453, g5841, g5763, g3747, g5637, g2912, g2357, g4232, g164, g4253, g5016;
wire g3119, g1351, g1648, g4519, g5115, g3352, g6657, g4552, g3893, g3211, g5654;
wire g929, g3274, g5595, g3614, g2894, g3125, g3325, g3821, g4141, g4570, g5272;
wire g2735, g728, g6295, g5417, g2661, g1988, g5128, g1548, g3106, g4659, g4358;
wire g1792, g2084, g3061, g3187, g4311, g2583, g3003, g1094, g3841, g4284, g3763;
wire g3191, g4239, g3391, g4180, g691, g534, g5366, g385, g2004, g2527, g5456;
wire g4420, g5148, g4507, g5348, g3223, g4931, g2970, g5698, g3416, g5260, g1521;
wire g3522, g3115, g3251, g1, g4628, g1996, g3447, g4515, g4204, g4300, g1724;
wire g1379, g3654, g12, g1878, g5619, g71, g59, I28349, g19408, I21294, g13297;
wire g19635, g32394, I19778, g9900, g11889, g13103, g17470, g23499, g6895, g9797, g31804;
wire g6837, I15824, g20066, g33804, g20231, I19786, g24066, g11888, g9510, I22692, g12884;
wire g22494, g9245, g8925, g34248, g10289, g11181, I20116, g7888, g9291, g28559, g21056;
wire I33246, g10288, g8224, g21611, g16718, g21722, I12530, g16521, I22400, g23611, g10571;
wire g17467, g17494, g10308, g27015, g23988, g23924, g12217, g14571, g32318, g32446, g14308;
wire I24041, I14935, g34778, g20511, g26672, g11931, g20763, g23432, I18165, I18523, g21271;
wire I31776, g23271, g22155, I22539, I32231, g34786, g9259, I15190, g17782, g8277, g9819;
wire I16969, g32540, g25027, g19711, g22170, g13190, g7297, g17419, g20660, g16861, g21461;
wire g10816, g28713, g15755, g23461, I24237, g34945, g8789, g31833, I18006, I20035, I17207;
wire g30999, g25249, g9488, g19537, g17155, I16855, g15563, g23031, g30090, g30998, g25248;
wire g23650, g7138, g16099, g34998, g23887, g25552, g20916, g27084, g30182, g7963, g10374;
wire I32763, g19606, g19492, g22167, g22194, g7109, g7791, g34672, g16777, g20550, g23529;
wire g6854, g18930, g13024, g32902, g6941, g12110, g32957, g9951, g32377, g12922, g23528;
wire g12321, g28678, g32739, g21393, g23843, g26026, g25081, g20085, g23393, g19750, g30331;
wire g24076, g24085, g17589, g20596, g34932, g23764, g25786, I25869, g32738, g32562, g32645;
wire g14669, g20054, I26337, g24054, I20130, g17588, g17524, I18600, g23869, g32699, g10392;
wire I28576, I28585, I15987, g14668, g25356, g24431, g29725, I15250, g28294, g8945, g10489;
wire g11987, g13625, I25161, g17477, g23868, g32698, g31812, g11250, g25380, I32550, g7957;
wire g13250, g20269, g34505, g7049, g20773, g25090, g6958, g20268, g14424, g34717, g12417;
wire g25182, g12936, g20655, g8340, g13943, g21225, g24156, g23259, g24655, I12109, I18063;
wire g7715, g29744, g8478, g20180, g17616, g20670, I29447, g10830, I32243, g22305, g24180;
wire g32632, g31795, g9594, g6829, g7498, g23258, g26811, I16590, g10544, g15573, I27492;
wire g9806, g14544, I14653, I33044, I16741, g25513, g32661, g20993, g32547, g32895, g8876;
wire g24839, g23244, g24993, g22177, g16162, g11855, g20667, g17466, g9887, g6974, g24667;
wire g9934, g21069, g25505, g34433, g34387, g10042, g24131, g32481, g14705, I13321, g18975;
wire g19553, g19862, g30097, g8915, g16629, I16150, g21657, g16472, I20781, g21068, g14255;
wire I21477, g14189, g32551, g32572, g23375, I24781, I33146, g7162, g25212, g7268, I11740;
wire g7362, g12909, g9433, g26850, g12543, g17642, g20502, g10678, I22725, I13740, g23879;
wire g20557, g23970, g34343, g20210, I22114, g12908, g20618, g11867, g11894, I11685, g8310;
wire g23878, g21337, g20443, g10383, g23337, g19757, g9496, g14383, g17733, I16526, g8663;
wire g10030, g23886, I18614, g32490, g10093, g18884, g27242, I14576, g11714, g22166, g11450;
wire I17114, I27192, g23792, g23967, g23994, g32784, g9891, I18320, g28037, g8002, g9337;
wire g9913, g32956, I21285, g11819, g11910, g14065, g7086, g13707, g31829, g32889, g11202;
wire g8236, g33920, I21254, g24039, g25620, g21425, g29221, I17744, g23459, I16917, g20038;
wire g23425, g31828, g32888, I15070, g25097, g32824, g10219, g13055, g9807, I30901, g19673;
wire g24038, g14219, g19397, g21458, g6849, I15590, g28155, I13762, g13070, g23458, g32671;
wire I21036, g34229, g10218, I18034, g16172, g20601, g21010, g11986, g7470, I12483, g17476;
wire g17485, I16077, I14745, g11741, g22907, g23545, g23444, g25369, g32931, g33682, g6900;
wire g19634, g19872, g34716, I20542, I25598, g8928, g29812, I28241, g12841, g22594, I16688;
wire g9815, g8064, I18408, I20913, g23086, I32815, g30310, g8899, g11735, g29371, I11908;
wire g9692, g13877, I32601, g8785, g24169, g24791, g9497, I16102, g26681, g20168, g9154;
wire g25133, g34925, I26309, g9354, g27014, I27564, g24168, g23322, g32546, g9960, g22519;
wire g22176, g14201, g26802, g28119, g12835, g7635, g14277, g20666, g13018, I16231, g32024;
wire g25228, I19802, g19574, g7766, g19452, g6819, g16540, I19857, g22154, g7087, I33297;
wire g25011, g32860, I18891, g7487, I33103, g8237, g18953, I14761, g19912, g17519, g21561;
wire I12183, g21656, g6923, g26765, I25680, g22935, g17092, g34944, g10037, I32791, g32497;
wire g21295, g23353, g29507, I32884, g8844, g11402, g17518, g26549, g17154, g22883, g20556;
wire g23823, g17637, g20580, g26548, g10419, g11866, g11917, g32700, I26687, g32659, g21336;
wire g32625, g10352, g23336, I32479, g19592, g34429, g10155, g10418, g12041, g32658, g19780;
wire g16739, g12430, I16660, g34428, I21074, g23966, g22215, g28036, g27237, g32943, g20110;
wire g11706, g24084, g16738, g9761, g13706, g16645, g12465, I11992, g24110, g20922, g27983;
wire g20321, g23017, g32644, g33648, I21238, g34690, g6870, g9828, g20179, g34549, g8948;
wire g20531, g12983, g24179, g16290, g32969, g13280, g6825, g33755, g17501, g7369, g27142;
wire g8955, g20178, g10194, g19396, g17577, g13624, I14241, I21941, g24178, g14167, g32968;
wire g19731, g29920, g34504, g29358, g7868, I15102, I26195, I11835, I20891, g9746, g20373;
wire g32855, g23289, g24685, g24373, I33024, g8150, g10401, g22906, g20654, I16596, g34317;
wire g8350, g18908, g32870, g7535, g32527, I13007, g8038, g10119, I24474, g16632, g21308;
wire g8438, g23571, g28693, g23308, g31794, g6972, g31845, g8009, I31497, g7261, g24417;
wire g33845, g10118, I19775, g9932, g28166, g28009, g16661, I17507, g25549, g13876, g13885;
wire g32503, g23495, I31659, g14749, g32867, g32894, I31625, g14616, g34245, I32953, g8836;
wire g30299, g6887, g23816, g25548, g34323, g34299, I32654, g22139, g8918, g24964, g7246;
wire I11746, g26856, g13763, g14276, g31521, I32800, g32581, g32714, g32450, g10053, g23985;
wire g22138, g15739, I26705, g34775, I20750, g20587, g32707, g32819, g9576, g31832, I20982;
wire g23954, g24587, g8229, g9716, I22788, I26679, g12863, g8993, g15562, g32818, g10036;
wire g32496, g19787, g16127, g8822, g10177, g20909, g20543, I13684, g31861, g9848, g21669;
wire g19357, g17415, g6845, g7502, I15550, g32590, g9699, g9747, g24117, g24000, I33197;
wire g23260, g19743, I14584, g33926, g25245, g34697, g26831, g20569, I20840, g34995, g23842;
wire g32741, g13314, I23348, g25299, g32384, I19831, g33388, I18252, I16502, g20568, g23489;
wire g25533, g13085, g19769, g24568, g20242, g25298, g11721, g7689, g29927, I17121, g34512;
wire g21424, g23559, g13596, g23525, g23488, g28675, g23016, I32909, g7216, g11431, g12952;
wire g23558, g13431, g32801, g14630, g32735, g24123, g32877, g7028, I30686, g8895, g10166;
wire g17576, g17585, g20772, g9644, g22200, g23893, I15773, g11269, I15942, g14166, g8620;
wire g19881, g8462, g25232, g29491, g7247, g20639, I17173, g16931, I16468, g23544, g23865;
wire I12046, g32695, I31581, g11268, g20230, g12790, g17609, g29755, g7564, g9152, g20638;
wire I18509, g9818, g13655, g34316, g17200, g32526, g20265, g29981, g6815, I12787, g12873;
wire I22028, I29211, g8788, I18872, I23333, g30989, g33766, g19662, g21610, g14454, g23610;
wire g10570, g34989, g8249, g20391, g32457, g21189, g24992, I33070, g20510, g23189, g11930;
wire g12422, g26736, g9186, g17745, g34988, g22973, g34924, g6960, g9386, I15667, I32639;
wire g21270, g32866, g32917, g23270, g19482, g21678, g17813, g12834, g20579, g34432, g7308;
wire g11965, g8085, g9599, g10074, g19710, g18983, g24579, g34271, g19552, g21460, g21686;
wire g9274, g20578, g26843, g23460, g23939, g21383, g19779, I19843, g9614, I33067, g17674;
wire g12021, g14238, g20586, g23030, g32706, g23938, g32597, I18574, g25316, g8854, g21267;
wire g24586, I32391, g23267, g9821, I13236, I18205, g34145, I16168, g26869, g32689, g15824;
wire g20442, g10382, I18912, I22240, g32923, g33451, g19786, I14833, g16659, g12614, g22761;
wire g9280, g10519, g34736, g10176, I16479, g27320, g16987, g32688, g32624, I23312, g13279;
wire I16217, I21115, g16658, I22604, g10518, g10154, g12905, g20615, g33246, g9083, g23875;
wire g25080, g24116, g14518, g23219, I18051, g30330, g13278, g26709, I29969, g8219, g27565;
wire I17491, I16486, g20041, g9636, g22214, g7827, g12122, g20275, g24041, g19998, g8431;
wire g11468, g16644, g13039, g8812, g15426, g22207, g6828, g19672, g34132, g17400, I12890;
wire g29045, g34960, g11038, g16969, g6830, g17013, I18350, g8005, g20237, g21160, g7196;
wire g11815, g8405, g9187, g16968, I27552, I15677, g31859, I32116, g20035, g31825, g32876;
wire g32885, g34161, g16197, g24035, g11677, g21455, I12003, g8286, g8765, g17328, g31858;
wire g13975, g32854, g7780, I12779, g16527, g25198, g30259, g25529, g14215, g32511, g23915;
wire g32763, I15937, I17395, I28434, g30087, g11143, g19961, g26810, I29894, I14033, g34471;
wire g9200, g25528, I21934, g31844, I31597, g8733, g19505, g23277, g7018, g8974, I11726;
wire I32237, I17633, g32660, g7418, I13726, g9003, g6953, g7994, g29997, g11884, g21467;
wire I16676, g25869, g10349, g23494, g26337, I32806, g8796, I32684, g32456, g34244, I33300;
wire g20130, g22683, g13410, I12826, g21037, g24130, g32480, g10083, g10348, g32916, g14348;
wire g12891, g8324, g26792, g20523, I16417, I21013, g32550, g9637, g23984, g18952, g24165;
wire g30068, g34810, g31227, g17683, g23419, g34068, g21352, g13015, g8540, g23352, g25259;
wire g25225, g21155, g34879, g21418, g22882, g28608, g23418, g32721, g20006, I26466, I15556;
wire g32596, g9223, g12109, g19433, g23170, g7197, g22407, g34878, g19387, I16762, g6848;
wire g7397, I27449, g15969, I20846, g19620, g12108, g10139, I15223, I17612, I24396, g6855;
wire g17414, g27492, g8287, I17324, g9416, g13223, g24437, g25244, g19343, g34994, I17098;
wire g32773, g32942, g9251, g20703, g29220, I11635, g23589, g10415, g18422, g32655, g8399;
wire g11110, g29911, g19369, g33377, g34425, g12381, g23524, g27091, g28184, g32670, g33120;
wire I12026, I21100, g8898, g20600, I16117, g34919, g19368, I32222, g20781, g16877, g23477;
wire g32734, g33645, g22759, I17140, g26817, g7631, g34918, g17584, I26693, g10664, I20929;
wire g32839, g32930, g20372, g30079, g19412, g7257, g22758, g24372, g16695, g25171, g20175;
wire g7301, I16747, g8291, g11373, g23864, g25886, g23022, g32667, g32694, g32838, I31550;
wire g33698, g24175, g29147, g32965, g12840, g6818, g17759, g6867, g16526, g23749, I15800;
wire g15714, g9880, g23313, g25994, g8344, g9537, g29950, g24063, g17758, g26656, g20516;
wire g10554, g18905, g24137, g32487, g24516, g7751, g23285, g26680, g32619, g8259, g21305;
wire g21053, g32502, g14609, g15979, g10200, g23305, g32557, g13334, g29151, g29172, I24787;
wire g9978, g30322, g10608, g29996, I12811, g10115, I16639, g21466, g32618, I18662, g8088;
wire g6975, g9417, g34159, g11762, g7041, g9935, I13606, g11964, g21036, g7441, g20209;
wire g33661, g33895, g9982, g21177, g21560, g16077, g9234, I15587, g32469, I27368, I18482;
wire g20208, g14745, g13216, g17141, I11750, I18248, g19379, g26631, g12862, g17652, g34656;
wire g8215, g30295, g22332, g9542, I16391, g26364, g32468, g6821, I18003, g19050, g34680;
wire g8951, g16689, g34144, g34823, g20542, g16923, g20453, g16280, g6984, g32038, g24021;
wire g28241, g29318, g16688, g16624, g22406, g8114, g10184, g12040, I16579, g16300, g19386;
wire g10805, I22785, g20913, I18778, g34336, g32815, g14184, g19603, g19742, g13117, g17135;
wire g12904, g20614, g32601, I15569, g9554, g20436, g23874, g8870, g32677, g33127, g25322;
wire I31694, I32834, g32975, g21693, g20607, g13569, g8650, I12896, g20320, I18647, g20073;
wire I28832, I33131, g30017, g20274, g9213, g24073, g20530, g21665, g25158, I21744, g20593;
wire I17754, g23665, g25783, I17355, g32937, g19429, I23345, g33385, I21849, g29044, g10761;
wire g7411, g25561, g18891, g20565, I31619, I15814, g24122, I23399, g8136, g19730, g19428;
wire g12183, g9902, I18233, g33354, I33210, g32791, g23476, g23485, I25555, g31824, g32884;
wire g33888, g8594, g19765, g6756, g24034, g7074, g11772, g10400, g20641, g26816, g21454;
wire I33279, g23555, I32607, g7474, g17221, g19690, g30309, g7992, g9490, I14563, g16511;
wire g9166, g20153, g23570, I32274, g23914, g32479, g32666, I13483, g11293, g24153, I31469;
wire g6904, g32363, I12112, g12872, g13638, g34308, g9056, g23907, g32478, g32015, g19504;
wire g9456, g33931, I32464, g8228, g9529, g7863, g20136, g20635, I27742, g13416, g25017;
wire I25567, I25594, I18897, g24136, g32486, I13326, g23239, g33426, g11841, g9155, I14395;
wire g6841, I17420, g23567, g32556, I32797, I14899, g8033, g23238, g11510, g13510, g17812;
wire g34816, I20647, g32580, g9698, g28441, g26260, I14633, g9964, I13252, g20164, g34985;
wire I20999, g23941, g18091, g19128, g23382, g24164, g25289, g21176, g21185, g23519, I27730;
wire g12047, g16307, g13835, g34954, g13014, g25023, g24891, I33143, g19626, g25288, g25224;
wire I20233, g16721, I12793, g23518, g23154, g26488, g26424, g20575, g31860, g13007, g25308;
wire g8195, g8137, g32922, g8891, g19533, g24474, g20711, I16193, g16431, I27549, g27051;
wire g32531, I13847, I31791, g20327, g23935, g24711, g34669, g26830, g27592, g12051, g20537;
wire g24109, g32740, g15885, g8807, g11615, g9619, g17507, I24331, g34668, g13116, g16773;
wire I18148, g24108, I28162, g32186, g34392, g32676, g32685, g33659, g28399, g30195, g7400;
wire g8859, g32953, g19737, g11720, g20283, g6811, g34195, g20606, g33250, g16655, g10882;
wire I18104, g10414, I13634, g31658, I13872, g13041, g32654, g9843, g33658, g16180, g30016;
wire g9989, I24448, g11430, g22541, g34559, g12350, g10407, g32800, g32936, g19697, I31486;
wire g23215, g12820, I17699, g23501, g6874, I29965, I32109, I21033, g20381, g8342, g11237;
wire g9834, g9971, I21234, g24982, g26679, g34830, g34893, g9686, g22359, g8255, g17473;
wire g20091, I22366, g24091, g7183, g8481, I12128, g17789, g29956, g29385, g34544, g15480;
wire I26664, g22358, g32762, g9598, g24174, g8097, g25260, g32964, g29980, g7779, g34713;
wire g8497, g13142, g21349, g8154, I28591, g17325, g8354, g18948, g7023, g31855, g10206;
wire g14441, g14584, g9321, g7423, g9670, I22547, g25195, g16487, g23906, g26093, g30610;
wire g18904, g32587, g15085, I32982, g23284, g19445, g10725, g21304, g25525, g34042, g25424;
wire I20433, g23304, g25016, g6978, I33179, g7161, g19499, g17121, g7361, g22682, g10114;
wire g20192, g9253, I16821, I17661, g27929, g25558, g23566, g32909, g10082, g32543, g34270;
wire I27232, g19498, g34188, g7051, g10107, g22173, g34124, g9909, g12929, g25830, g27583;
wire g20663, g27928, g25893, g8783, g7451, g32908, g6982, g7327, g24522, g33894, g11165;
wire g8112, g8218, g34939, g9740, g8267, g25544, g32569, g34383, g29190, I32840, g17291;
wire g14744, g16286, g21139, g21653, g26837, g7633, g34938, g23653, g9552, g15655, I31800;
wire g10399, g32568, g32747, I18310, I20369, g18062, g21138, g24483, g19432, I19837, g30065;
wire I11820, g23138, I26799, g20553, g31819, g8676, I15727, I32192, g10398, I18379, g14398;
wire g10141, g29211, g10652, g10804, g6800, I13152, g9687, g31818, g32814, g20326, g23333;
wire g13222, g19753, g16601, g17760, g16677, I22889, g20536, g20040, g13437, I20412, g32751;
wire g32807, g32772, g28463, g32974, g8830, g24040, g7753, g20702, g30218, g25188, g32639;
wire g20904, I17956, g23963, g19650, g28033, g8592, g7072, g14332, I11691, I28540, g32638;
wire g7472, g19529, g12640, I15600, g22927, g9860, g10406, I24228, g20564, g10361, I25576;
wire g7443, g8703, g14406, g19528, g19696, g34160, g25267, g19330, I17181, I17671, I29363;
wire g23585, g32841, g11236, I21291, g7116, g22649, g10500, g27881, g19365, g20673, g32510;
wire g9691, g31801, I15821, I12056, g24183, I32904, g14833, g19869, g21609, g19960, g23609;
wire g24397, g29339, g12881, g7565, g22903, g13175, g34915, I16593, I25115, g32579, g8068;
wire I13020, I32621, g23312, I31569, I28301, g25219, I27271, g21608, g24062, g17649, g20509;
wire g23608, g34201, g9607, g24509, g32578, g32835, g33695, g34277, g25218, g9962, g11790;
wire g14004, g17648, g20508, g9158, g27662, g17491, g22981, g20634, I21029, g21052, g28163;
wire g8677, g25837, g7533, g19709, g32586, I22211, g9506, g17604, g34595, g7697, g10613;
wire g23745, I18504, I22024, g32442, I31814, g19471, g30037, g12890, g16580, g23813, g7596;
wire I31751, I31807, g16223, g10273, g33457, I32062, I12199, g10106, g9311, I11743, g22845;
wire I12887, g34984, g32615, I15834, g13209, g8848, g20213, I15208, g33917, g21184, g34419;
wire g9615, g21674, g10812, g32720, g30155, g8398, g28325, g12779, g22898, g9174, g34418;
wire g17794, g26836, g17845, g9374, g20574, g20452, I15542, g32430, g10033, g10371, g32746;
wire g32493, g22719, g24452, I26100, g7936, g9985, g24047, g12778, I18245, I12764, g23732;
wire g8241, I20793, g20912, g19602, g32465, g7117, I18323, g19657, g22718, g16740, I12132;
wire g19068, g15169, g28121, g9284, g19375, g10795, I25692, g9239, g33923, g9180, g16186;
wire g16676, g16685, I20690, I29936, I17658, g9380, g12945, g31624, g32806, g20072, g32684;
wire g33688, g29707, g9832, I15073, g19878, g24051, g24072, g34589, g17718, g17521, g16654;
wire g20592, g27998, I16575, g15479, g9853, I15593, g8644, g6989, g9020, g24756, I32452;
wire I12709, g21400, g20780, g7922, g8119, g13530, g23400, g12998, g34836, g13593, g28173;
wire g18929, g32517, g23013, I28572, g12233, I31586, g23214, g11122, I14902, I14301, g12182;
wire g29978, g12672, g7581, g21329, g22926, g25155, g9559, g13565, g6971, g8818, I25005;
wire g14421, I19704, g25266, g25170, g9931, g23539, g17573, g7597, g11034, g23005, g13034;
wire g17247, I32051, g30022, g34118, I16606, g15580, g12932, g23538, g34864, I16492, g17389;
wire g17926, g16964, g24152, g19458, g30313, g34749, g17612, g24396, g8211, g29067, g9905;
wire g10541, g16423, g27961, g8186, g34313, I13552, g10473, g17324, g32523, I24128, g31854;
wire g14541, g16216, I29909, I33041, g12897, g13409, g16587, g17777, g25167, g25194, I13779;
wire I26584, g9630, g29150, g34276, g34285, g7995, g30305, g11136, g30053, g8026, g25524;
wire I27970, g18827, g34053, g7479, g9300, g10359, I32820, g8426, g32475, g14359, g8170;
wire g7840, g22997, g32727, g10358, g33660, g32863, g29196, I32846, g14535, g24405, g8125;
wire g30036, g14358, g25119, I22819, g8821, g16000, g15740, I25683, I29242, g32437, g14828;
wire g23235, g33456, g10121, g11164, g25118, g26693, g8280, g23683, g15373, g9973, g33916;
wire I22111, g7356, I17819, g16747, g20583, g32703, I12994, I15474, g24020, g19532, g22360;
wire g9040, g28648, g18881, I13672, g13474, I25882, g20046, g9969, g19783, I17111, g16123;
wire g24046, g17871, g16814, g21414, g32600, g7704, I16663, g23515, g28604, g23882, g23414;
wire g32781, I23099, g31596, g8106, g14173, I23324, g20113, g21407, g31243, I17590, g19353;
wire g24113, I32929, g32952, g19144, g12811, g27971, g8187, g32821, g8387, g25036, I31523;
wire g7163, g29597, g25101, g20105, g24357, g25560, g10029, g8756, g22220, g13303, g24105;
wire I17094, I18031, g29689, g14029, g29923, g25642, g32790, g9648, g32137, g10028, g9875;
wire g32516, g31655, I29579, g28262, I24445, g20640, I17801, g20769, g17472, I26406, g12368;
wire I16040, I20499, I12086, g33670, I31727, g32873, g8046, g25064, g16510, g19364, g20768;
wire g28633, g8514, I19238, g34570, g34712, g21725, g11796, g16579, g33335, g8403, g23759;
wire g13174, I21766, I17695, g26941, g34914, g31839, g33839, I32827, g8345, g8841, I14671;
wire g7157, I12159, g22147, g26519, g16578, g15569, g8763, I16564, g23435, g31667, g31838;
wire g23082, g32834, g9839, g30074, g26518, g17591, g12896, g17776, g27011, I27561, g15568;
wire g15747, g25009, I13723, I26004, I18868, I23360, g18945, g30567, I30962, g17147, g22858;
wire g34594, I13149, g17754, I16847, g26935, g25008, g32542, g8107, I32803, I25399, g31487;
wire g32021, g32453, I29720, g11192, g22151, I11620, I21162, I12144, I12823, I18709, g20662;
wire g21399, g23849, g22996, g23940, g25892, I20753, I15663, g23399, g32726, g32913, g24027;
wire I18259, g9618, g11663, g16615, g22844, g13522, g34941, g13663, g21398, g23848, g25555;
wire g32614, g7626, I12336, g23398, I32881, g8858, g33443, g16720, g9282, g34675, I20650;
wire g23652, g32607, g8016, g10981, g8757, g32905, g14563, g8416, g27112, g20710, g16746;
wire I20529, I21911, g17844, g20552, g32530, g9693, g13483, I33264, I15862, g17367, g32593;
wire g18932, g6985, I33137, g20204, g19687, I21246, g24003, g23263, I12631, g8522, g20779;
wire g22319, g12378, g34935, g23332, g32565, g32464, g25239, g19954, g11949, I24393, g19374;
wire g20778, g34883, g10794, g9555, g18897, I15536, g10395, g22227, g24778, g9804, g10262;
wire g24081, g21406, g16684, g11948, I21776, I15702, g14262, g12944, I18810, g23406, g9792;
wire g32641, g6832, g32797, g23962, g31815, g23361, g28032, I32482, g11702, g7778, g15579;
wire g31601, g8654, I16452, I18879, g9621, g10191, g23500, g24356, g13621, g21049, I11896;
wire g25185, g17059, g20380, g26083, g14191, g30729, I15564, g25092, g24999, g26284, I18337;
wire g34501, g27730, g10521, g12857, I19348, g21048, g25154, g20090, g17058, g32635, g8880;
wire g31937, g8595, g24090, g19489, g20233, g33937, g12793, I11716, g20182, g20651, g20672;
wire I17876, g23004, I27495, g7475, g21221, g24182, g19559, g23221, I14644, g11183, g29942;
wire g22957, g31791, g7627, g19558, g6905, g16523, g8612, g23613, g9518, g15615, I17763;
wire I31607, g13062, g7526, g7998, g11509, g22146, g26653, g20513, g17301, g20449, g28162;
wire g10389, g32891, I15872, g13933, g23947, g31479, g31666, I27954, g18097, g21273, g17120;
wire g19544, g23273, g19865, g17739, g10612, g11872, g23605, g9776, g10099, g15746, g16475;
wire g20448, g34304, I12954, g10388, I32651, g32575, g32474, g19713, g7439, g29930, g22698;
wire g29993, g16727, g17738, g17645, g20505, g21463, g23812, g32711, g8130, g14701, I17456;
wire I23318, g8542, g24505, g8330, g24404, g10272, g9965, g29965, I33034, g14251, I17916;
wire g20026, g32537, I18078, g20212, g23234, g24026, g9264, g15806, I21058, g25438, g6973;
wire I17314, I32449, g19679, I18086, g27245, g34653, g9360, g9933, g32606, g10032, I29236;
wire g32492, g19678, I15205, g14032, g10140, g29210, g9050, g17427, I13802, g13574, I25514;
wire I13857, g17366, g7952, g25083, g25348, g9450, I14450, g16600, g19686, g25284, g21514;
wire I11793, g11912, g26576, I26682, g28147, I27558, g32750, I12016, I18125, g10061, g13311;
wire g28754, g32381, g7616, I19484, g23507, g34852, g20433, g25566, g18896, g24149, g20387;
wire g28370, I28866, I22180, g16821, g21421, g27737, I12893, g7004, g9379, g23421, g13051;
wire g20097, g32796, g7527, I33164, g24097, g26608, g11592, g20104, g7647, g34664, I27713;
wire I13548, g10360, g23012, g24104, g17226, g25139, g17715, g6875, g9777, g17481, I25541;
wire g32840, I28597, g28367, I31474, g24971, g27880, g25138, g34576, g16873, g23541, g31800;
wire g12995, g7503, g7970, g13350, g23473, g33800, g8056, I13317, g11820, g33936, g8456;
wire g12880, I22131, I24078, g23789, I17839, g32192, I33109, I15846, I16357, I25359, I19799;
wire g30312, I12189, I19813, g24368, g21724, g23788, g8155, g34312, g26973, g34200, g7224;
wire g32522, g23359, g32663, g8355, g8851, I13057, g14451, I23366, I18364, I22619, I17131;
wire I22502, g22980, g21434, I22557, g21358, g6839, g23434, g24850, g30052, I19674, g8964;
wire I29913, g27831, I11626, g11413, g34921, g13413, g34052, g23946, g24133, g29169, g18096;
wire g18944, g20229, g32483, g19617, g19470, g22181, g11691, g19915, g12831, g26732, I16803;
wire I12030, I17557, g9541, g32553, g32862, g7617, g16726, I26649, g34813, g10776, g19277;
wire g32949, g9332, g14591, g14785, I21226, I22286, g7516, g21682, I18224, g9680, g9153;
wire g10147, g20716, g27989, g29217, g34973, g25554, I15929, I18571, g21291, g32536, g14147;
wire g30184, I31796, g10355, g32948, g23291, g16607, g19494, g11929, I11737, g34674, g8279;
wire g16320, g20582, g32702, g9744, g10370, g31000, g32757, g32904, g6988, I14866, g16530;
wire g26400, g11928, g25115, g13583, g32621, g8872, g22520, I22601, g10151, g28120, I32228;
wire I11697, g10172, g20627, I12837, g7892, g34934, g9558, g20379, g8057, g32564, I13995;
wire g24379, g8457, g8989, g19352, g22546, g23760, g20050, g23029, g6804, g24112, g10367;
wire g10394, I25028, g24050, g9901, g34692, I22143, I21784, g23506, g23028, I18752, I28480;
wire g31814, g32673, g32847, g20386, I21297, g8971, g22860, g24386, g20603, g9511, g27736;
wire g7738, g31807, g8686, g13302, g20096, g24603, g33772, g7991, I23354, g24096, g29922;
wire g34400, g7244, g12887, g10420, I17143, g22497, g25184, g32509, g31639, g10319, g17088;
wire g32933, g30329, g9492, I21181, g16136, g7340, g20681, g9600, I23671, g32508, g9574;
wire g31638, g9864, g32634, g32851, g32872, g33638, g35001, g30328, g7907, g11640, g11769;
wire g34539, g9714, g12843, g17497, g22987, g34328, g10059, g23927, I18842, g24429, g19524;
wire I29891, g7517, g22658, g29953, g10540, g10058, g31841, g24428, I32096, g33391, g19477;
wire g12869, g16164, g23649, g26683, g7876, g25692, g15614, g22339, g20765, g8938, I19235;
wire I20495, g29800, g10203, g12868, g21903, g14203, g20549, g23648, g13881, I16090, g22338;
wire g23491, I20816, g23903, I33252, I32681, g10044, g34241, g27709, g21604, I22580, I16651;
wire g20548, g8519, g8740, g31578, g25013, g31835, g32574, I20985, g24548, I31564, g17296;
wire g25214, g27708, I12418, g17644, g20504, g30100, g23563, g10377, g32912, g8606, I18865;
wire I20954, g19748, g10120, g22197, g14377, I11753, g22855, g19276, g9889, g13027, g7110;
wire I14660, g33442, g22870, g22527, I21860, g34683, g28127, g25538, g29216, I32690, g11249;
wire I28838, I13031, g14738, g13249, g14562, g14645, I30861, g20129, g16606, g17197, g18880;
wire g23767, g23794, g21395, g24129, g32592, g20057, g32756, g23395, g24057, g20128, I12167;
wire g14290, g17870, g17411, g17527, g23899, g7002, g13003, g24128, g11204, I14550, g7824;
wire g30991, g6996, g25241, g11779, I18270, g16750, g22867, g34991, g7236, g9285, g20626;
wire g27774, I27401, I11843, g23898, g9500, g20323, I21250, g29117, g24626, g33430, g23191;
wire g20533, g10427, g12955, g32820, I18460, g8341, g10366, g24533, g25100, g12879, g22714;
wire g11786, g14366, g17503, I14054, g9184, g23521, g28181, g25771, g20775, g18831, I15647;
wire I23339, g32846, g9339, I19759, g19733, I24558, g12878, g26758, I27749, I20830, g12337;
wire g32731, g31806, g22202, g33806, g9024, I12749, g11826, g17714, g12886, g22979, g20737;
wire g22496, g10403, I21969, g23440, g13999, g7222, g27967, g27994, g33142, g19630, g9809;
wire g20232, I14773, g29814, g17819, g17707, I33047, g30206, g7928, g26744, g12967, g23861;
wire g23573, g32691, g18989, g8879, g8607, g11233, I18875, g21247, g23247, g11182, I11708;
wire g7064, g17818, g9672, I13708, g20697, g14226, g9077, g17496, I19345, g22986, g8659;
wire g25882, g23926, g8358, g18988, I32775, g9477, g8506, I30766, g9523, g24995, g34759;
wire g7785, g16522, g23612, g10572, I25534, I17964, g23388, I15932, g17590, g19476, g12919;
wire I12808, g6799, g26804, g20512, g34435, g23777, g23534, I26451, g13932, g32929, g8587;
wire I14839, g23272, g11513, g19454, g7563, g17741, g12918, I18160, I15448, g17384, g32583;
wire g32928, g19570, g19712, g6997, g22150, g11897, I22000, g10490, g9551, g9742, g9104;
wire g23462, g9099, g34345, g9499, g11404, g15750, g34940, g13505, I15717, g16326, g18887;
wire g20445, I31820, I12064, g23032, g10376, g10385, g25206, g12598, g14376, g14385, g34848;
wire g19074, g17735, g14297, g20499, g7394, g10980, g11026, I26785, g12086, g32787, g13026;
wire g31863, I14619, g10354, I23315, I33152, g19567, g14095, g29014, g22526, I17569, g9754;
wire g21061, g28126, g18528, g20498, g6802, g8284, g23061, g8239, g28250, g10181, g25114;
wire g7557, g8180, I17747, g12322, g27977, g32743, g32827, g25082, g8591, g30332, g24056;
wire g9613, g12901, g20611, g17526, g12977, g20080, g7471, g9044, g20924, g19519, g24080;
wire g19675, g9444, g9269, g22866, I17814, g32640, g20432, g32769, g23360, g29116, g19518;
wire g8507, g9983, g12656, I15620, I17772, g25849, g9862, I27555, g23447, g32768, g32803;
wire g25399, g12295, I23384, g10190, g29041, g13620, g12823, I17639, I27570, I15811, I21067;
wire I18822, g16509, I32056, g11811, I12712, g20145, g34833, g34049, I13010, g31821, g32881;
wire I32988, g24031, I33020, g16508, I24455, g26605, g20650, g23629, g21451, g16872, I12907;
wire g22923, I17416, g23472, g15483, g9534, g9729, g9961, g7438, g25263, g29983, g20529;
wire g22300, g26812, I21019, g27017, I27567, g15862, g8515, g34221, g8630, g21246, I27238;
wire g23246, g20528, g20696, g25135, g20330, g9927, g32662, g8300, g32027, I32461, g19577;
wire g17688, g9014, g20764, g10497, I25591, g32890, I33282, I27941, g9414, g7212, g19439;
wire g9660, g9946, g20132, g24365, g20869, g13412, g23776, g34947, I12382, g24132, g32482;
wire g24869, g24960, g19438, I12519, g17157, I12176, g9903, g13133, g32710, I12092, g14700;
wire g21355, g32552, g31834, g23355, g34812, g10658, g21370, g23859, g28819, g16311, g32779;
wire I17442, g18878, g24161, g29130, I32696, I32843, g7993, g20709, g11011, g22854, g34951;
wire g34972, g23858, g13011, I12935, g32778, g18886, I31803, g9036, I18313, g25221, I22275;
wire g8440, g20708, g22763, g9679, g23172, g13716, I17615, g20087, g32786, g33726, I32960;
wire g8123, g19566, g14338, g24087, I18276, I18285, g28590, g23844, g32647, g23394, I32868;
wire g9831, g32945, g33436, g22660, g15509, I19012, g17763, g8666, g10060, I18900, g27976;
wire g27985, I32161, g32826, g25273, g29863, g24043, g10197, I21300, g22456, g12976, g15634;
wire I23688, I23300, g14197, g32090, g9805, g9916, g19653, g33346, I18101, I32225, g10527;
wire I12577, g10411, g23420, g9749, I18177, I18560, g32651, g18918, g32672, I19789, g24069;
wire g22550, I33027, g26788, g26724, g20657, g20774, I26427, g8655, g23446, I16057, I28908;
wire g19636, g23227, g30012, g19415, g24068, g24375, g21059, I33249, g7462, g23059, g31797;
wire g6838, g13096, g33641, g32932, g33797, I31482, g19852, g22721, g10503, I16626, g21058;
wire g6809, g32513, I20864, g23058, g32449, g14503, g16691, I24022, g19963, g12842, g34473;
wire I12083, g17085, I31779, g24171, g32897, g32961, g23203, g8839, g34789, g7788, g11429;
wire g17721, g29372, g10581, I16775, g13857, g32505, g20994, g9095, g32404, I14800, g33136;
wire g9037, g14714, g33635, g24994, g14315, g30325, g34788, g11793, g11428, g26682, g9653;
wire g17431, g13793, g22341, g32717, g34325, I15765, I18009, g21281, g18977, I31786, I32970;
wire g22156, g27830, g21902, g34920, g8172, g8278, g34434, g23902, g23301, g34358, g28917;
wire g23377, I32878, g22180, g24425, g19554, g10111, g12830, g12893, I11816, g16583, g7392;
wire g20919, g15756, I25146, g34946, I25562, g19609, g8235, g8343, I18476, g34121, I14964;
wire g19200, g21562, g9752, g12865, g20010, g8282, g20918, g23645, g8566, I18555, g24010;
wire g9917, I32967, I32994, g10741, I21480, g7854, g13504, g25541, g20545, g20079, g20444;
wire g21290, g32723, I31672, g10384, g8134, g23290, I33182, I13374, g8334, g24079, g21698;
wire g14384, g22667, g34682, g29209, g20599, g6926, I16512, g23698, I12415, g11317, g20078;
wire I12333, g32433, g19745, g24078, g6754, g12705, g20598, g32620, I28579, g20086, g19799;
wire g25325, I32458, g11129, I25366, g8804, g10150, g24086, g16743, g21427, g15731, g9364;
wire g10877, g23427, g25535, g32811, I12963, g14150, g21366, g32646, g8792, g7219, g19798;
wire I28014, g11128, g7640, I18238, g10019, g28157, I15626, g22210, g20322, g32971, g7431;
wire I32079, g7252, g16640, g29913, g34760, g7812, g16769, g20159, g34134, g25121, g20901;
wire g13626, g20532, g17487, I27576, I15533, g24159, g13323, g24125, g6983, I18382, g21661;
wire g17502, g16768, I19927, g20158, g8113, g12938, I16498, g23403, g23547, g23895, I13424;
wire g24158, g33750, I18092, g7405, g13298, g19732, I22264, I30980, I24008, g29905, g20561;
wire g20656, g9553, I18518, I18154, g23226, g7765, g20680, g26648, g20144, g10402, g23715;
wire g23481, g32850, g31796, g19761, I12608, g12875, I21734, g6961, g8567, I21930, g34927;
wire g7733, I22422, I15697, I17873, g31840, I32158, g12218, g32896, g12837, g23127, g6927;
wire I21838, g25134, g10001, g22975, g13856, I23694, I29248, g9888, g10077, g13995, I33149;
wire g8593, g29153, g24966, g7073, I12799, g20631, g17815, g10597, g23490, g25506, g9429;
wire I13705, I29204, g32716, g7473, g16249, g18976, g14597, g19539, g6946, g24017, g11512;
wire g34648, g24364, g17677, g34491, I22542, g16482, I17834, g31522, g32582, g7980, g21297;
wire g18954, g23376, g23385, I25095, g19538, g6903, g7069, g9281, I12805, g26990, g34755;
wire g23889, I13124, I18728, I21210, g23354, I14579, g22169, I26700, g34770, g12470, g7540;
wire g8160, g22884, g34981, g23888, g23824, I15831, g32627, g28307, g32959, g32925, g21181;
wire g22168, g10102, g10157, g31862, g32958, I15316, I19719, g8450, g24023, g26718, I32364;
wire g17791, g20571, g9684, g11316, g9745, g12075, I17436, g28431, g9639, I18906, g9338;
wire g24571, g10231, I18083, g9963, I26296, g33326, g17410, I12761, g11498, g34767, g14231;
wire g26832, g34845, g32603, g6831, I22464, g23931, g32742, I29233, g9309, I23306, g30990;
wire I18304, g19771, g25240, g32944, I29182, g29474, g34990, g11989, I25190, g16826, g17479;
wire g21426, g8179, g12037, g20495, g23426, g25903, g27984, I13875, g33702, g9808, g19683;
wire g23190, I16709, g11988, I21815, g17478, g28156, I12013, g17015, g32681, I32309, I12214;
wire g16182, g16651, I22153, g23520, g27155, g9759, g18830, I16471, g17486, g7898, g25563;
wire g32802, g32857, g22223, g13271, g34718, g24985, g34521, g32730, g23546, I24215, g32793;
wire I18653, g20374, g23211, I30644, g19882, g19414, g26701, g7245, g17580, g11753, I29961;
wire I12538, g26777, g20643, I18138, g9049, g23088, g31847, g32765, g19407, g9449, g16449;
wire g11031, g22922, g23860, I15650, g32690, g9575, g32549, I15736, I14684, I18333, g22179;
wire I29717, g25262, I11617, g11736, g20669, I17136, g16897, I26503, g34573, g7344, g25899;
wire g13736, g32548, I18852, I32687, g34247, I32976, I32985, g22178, g9498, g6873, g20668;
wire g34926, g32504, g31851, I15843, I32752, g9833, g10287, g7259, g21659, I33050, g14314;
wire g16717, g17531, g12836, g20195, I26581, g8997, g23987, g10085, g8541, g23250, g24489;
wire I23363, g14307, I27235, g17178, g6869, g34777, g12477, g20525, I15869, g18939, g8132;
wire g28443, g34272, g24525, g24424, I11623, g13132, g17685, g17676, g13869, g20558, g8680;
wire g22936, I13623, I21486, g17953, I22327, g23339, g8353, g18938, g23943, g18093, I13037;
wire I29149, g14431, g31213, g11868, g12864, g13868, g6917, g8744, g23338, g18065, g24893;
wire g12749, g19435, g9162, g9019, g17417, I18609, g7886, g20544, g23969, g32626, g28039;
wire I32195, I13352, g11709, g30997, g10156, g20713, g21060, g34997, I12991, g23060, g23968;
wire g18875, g32533, g8558, g28038, I32525, g13259, g33912, g19744, g16620, g7314, g10180;
wire I14006, I17108, I14475, g11471, g19345, g25099, g13087, g32775, g25388, g25324, I14727;
wire g13258, g12900, g19399, g20610, g7870, g21411, g17762, g20705, g34766, g23870, I16010;
wire g23411, g23527, g28187, I14222, I21922, g25534, g15932, g25098, g10335, I23321, g7650;
wire g27101, g25272, g29862, g24042, g33072, g20189, g19398, g20679, I29368, g17423, g16971;
wire g11043, g12036, g9086, g32737, I18813, g17216, g20270, g9728, g19652, I30986, I17750;
wire g22543, g17587, g9730, I31504, g24124, g8092, g14694, g29948, g8492, g9185, g23503;
wire g23894, g19263, g32697, g27064, I18674, g25032, g20383, g32856, I28913, g11810, g25140;
wire g9070, g8714, g7594, g31820, g10487, g32880, g13068, g25997, g7972, g24030, g20267;
wire g24093, g10502, g26776, g23714, I27758, g23450, I29228, g32512, g7806, I15878, g20065;
wire g31846, g7943, g24065, g11878, g19361, I20609, I12758, g23819, g12874, g26754, g34472;
wire g25766, g28479, I32678, g23202, g14443, g23257, g26859, g27009, g26825, g21055, g23496;
wire g7322, g16228, g20219, g23055, g6990, g17242, g34246, g10278, g33413, g29847, I29582;
wire g23111, g12009, g21070, g6888, g22974, g32831, g33691, g32445, I32938, I32093, I13276;
wire g16716, g9678, g10039, g10306, g32499, g23986, g30591, g6956, g18984, g8623, I11809;
wire g34591, I18214, g12892, g34785, g16582, g17772, g34776, g11425, g10038, g32498, g23384;
wire g17639, I12141, g34147, g9682, g9766, g15811, g16310, g7096, g10815, g13458, g24160;
wire I15918, g9305, g7496, g33929, g16627, g17638, g22841, g34950, g12914, g13010, g32611;
wire g7845, I33232, g25451, g32722, g25220, g32924, g33928, g19947, g7195, g12907, g20617;
wire g17416, g7395, g7891, g8651, g16958, g9748, g13545, g23877, g19273, g20915, g7913;
wire g27074, g28321, I32837, g30996, g25246, g34151, I12135, g10143, g29213, g34996, g23019;
wire I33261, g8285, g12074, I25695, g9226, g20277, g16603, g16742, g23196, g34844, I22564;
wire g16096, g23018, g32753, g12238, g32461, I21242, g10169, g24075, g17579, g19371, g20595;
wire g23526, g6808, g20494, g14169, g8139, I16289, I32455, g7266, g29912, g29311, g10410;
wire g20623, g27675, I12049, g9373, g17014, g27092, g9091, g20037, g31827, g32736, I32617;
wire g13322, g32887, I32470, g24623, g33827, g9491, I14905, g24037, g34420, g16429, I11665;
wire g20782, g21457, g13901, g23402, I13166, g32529, g23457, g25370, g8795, g10363, I24400;
wire g10217, I14593, g30318, g14363, g14217, g9283, I14346, g16428, g9369, g32528, g32696;
wire g9007, I21230, g32843, g6957, g24419, g32393, g9407, I15295, I11892, g34059, g8672;
wire g9920, I15144, I13892, g31803, g32764, g24155, g24418, I32467, g20266, g8477, g34540;
wire g11823, g13680, g17615, g12883, g13144, g22493, g7097, g23001, g34058, g24170, g32869;
wire I18882, g32960, I18414, g7497, I14797, g19421, g17720, I33056, I25689, g9582, g11336;
wire g7960, g32868, g8205, I32782, g10223, g21689, g23256, I12106, I12605, g17430, g17746;
wire g20853, g34044, g21280, g23923, I14409, g29152, g29846, I32352, I29002, g21300, g20167;
wire g20194, g20589, g32709, g11966, g23300, I12463, g17465, g8742, g13966, g10084, g24167;
wire g9415, g19541, g30301, g10110, g11631, g19473, g18101, g11017, g20588, g20524, g32708;
wire I32170, I12033, g13017, I28174, I29245, g32471, g19789, g24524, g24836, g16129, g25227;
wire g14321, g34739, g10531, g17684, g27438, g14179, g25025, g7267, g24477, g10178, g26632;
wire g24119, g27349, I31650, g23066, I28390, g9721, g23231, g34699, g19434, g16626, g8273;
wire g10685, I16489, g16323, g24118, g10373, g14186, g14676, g24022, g34698, g7293, g12906;
wire g16533, g20616, I18114, g23876, I18758, g13023, g18874, I31528, g25044, I19661, g29929;
wire g16775, I18107, g10417, I25511, g32602, g32810, I13637, I20882, g32657, g32774, g33778;
wire g7828, g32955, g21511, g29928, I26670, g20704, g23511, g34427, I32119, g32879, g8572;
wire g20053, g32970, g10334, g19682, I14537, g24053, g25120, I17780, g17523, g20900, g8712;
wire g7592, I16544, I18849, g18008, g32878, g31945, g21660, g24466, I16713, g9689, g10762;
wire g25562, g18892, g20036, g31826, g32886, I33161, I18398, g20101, g24036, I12541, g20560;
wire g16856, g21456, I26667, g11985, g17475, g24101, I23684, g32792, g23456, g13976, g24177;
wire g24560, I15954, g32967, g10216, g14423, g8534, I16610, g9671, g20642, g23480, g27415;
wire I20584, g23916, g9030, g19760, I32305, I14381, g16512, I16679, g23550, g26784, g9247;
wire I33258, I32809, g18907, g7624, g32459, g20064, g7953, g30572, g24064, g28579, g9564;
wire I18135, g23307, g32919, g23085, g32458, I24759, g14543, g33932, g9826, g10117, g10000;
wire g26824, I16460, g20874, g21054, g32918, g23243, g20630, g11842, g21431, g9741, g8903;
wire g23431, I13906, g32545, g9910, g17600, I19671, g34490, g20166, g20009, I22583, g27576;
wire g27585, g20665, g25547, g32599, I20744, I31810, g9638, g21269, g24166, g24665, g7716;
wire g7149, g34784, g7349, g30297, g27554, g20008, g34956, g17952, g32598, g13016, I22046;
wire g23942, I20399, g23341, g18092, g21268, I14192, I18048, I28062, g25226, g22137, g21156;
wire g17821, g8178, g6801, I21006, g28615, I16875, g25481, I15893, I31878, g19649, I32874;
wire g21180, I14663, g21670, I18221, g16722, g16924, g20555, g32817, I28851, I28872, I32693;
wire g8135, I21222, g19491, g34181, g34671, g20570, g20712, g11865, I22302, g13865, g20914;
wire g21335, g18883, g32532, g32901, g14639, g10230, g23335, I32665, g19755, g6755, g12921;
wire g23839, I17787, g17873, g23930, g23993, g32783, g19770, I29199, g30931, g8805, I14862;
wire g8916, I16160, g21694, g23838, g9861, g10416, I15705, g9048, I17302, g32561, g32656;
wire g23965, I31459, g20239, I32476, g11705, I22640, g24074, I22769, g26860, I14326, g34426;
wire g11042, g16031, g20567, g20594, g32680, g10391, I16455, g32823, g20238, g25297, g13255;
wire g9827, g13189, g22542, g13679, g28142, g31811, g23487, g14510, g31646, g9333, I14702;
wire g19794, g11678, g12184, g16529, g29081, g12805, g13188, g19395, g23502, I27927, g20382;
wire I16201, I23351, I31545, I23372, g26700, g7258, I33079, g11686, g16528, g7577, g7867;
wire g13460, g15831, I26479, I12927, g26987, g11383, g10014, g23443, I15030, I18795, g21279;
wire g24176, g24185, g23279, g32966, g19633, g7717, g30088, g24092, I32074, g29945, g6868;
wire g11030, g20154, g22905, g32631, g19719, g21278, g11294, g24154, I32594, g8037, g23278;
wire g13267, g29999, g32364, g6767, g17614, g22593, g9780, g16960, g20637, g26943, g8102;
wire g13065, g19718, g21286, g8302, g14442, g29998, g17607, g21468, g17320, g21306, g31850;
wire g8579, g23306, I29225, I31817, g7975, g33850, g17530, g10116, g9662, g9018, g11875;
wire g8719, g27013, g7026, I32675, g9467, g19440, g16709, g17122, g34126, g34659, I12770;
wire I12563, g12013, g23815, g34987, I25677, I15837, I33158, g7170, g19861, g10275, g19573;
wire g8917, g16708, g22153, g21677, g33228, g10430, g14275, g25546, g32571, I31561, I17249;
wire g25211, I32935, g22409, g19389, g17641, g20501, g26870, g30296, g20577, g34339, g9816;
wire g34943, I20951, g25024, g33716, I31823, g19612, g34296, g7280, g29897, g7939, g22136;
wire g29961, g8442, g22408, g22635, I12767, g14237, g8786, g23937, g10035, g32495, g29505;
wire g19777, g17409, I12899, g7544, g8164, g9381, I15617, I13805, I18788, g8364, g32816;
wire I15915, g24438, g11470, g17136, g10142, g17408, g34060, g29212, g7636, g9685, I26676;
wire g9197, I18829, g32687, g9397, I18434, g33959, g9021, I12719, g16602, g21410, g34197;
wire I27718, I16401, g16774, g23410, g8770, I29337, g34855, I26654, I22380, g16955, g32752;
wire g8296, g25250, g27100, g32954, g8725, g24083, g33378, g21666, g23479, I26936, g32643;
wire g6940, I15494, g13075, g23363, I18344, g7187, g7387, g20622, g11467, g13595, I17999;
wire g20566, g7461, I15623, g23478, g13494, g23015, g8553, I26334, I19707, g25296, g10130;
wire g16171, g33944, g19061, g26818, g16886, I27573, g32669, I15782, g23486, g26055, g13037;
wire g10362, g29149, g7027, I19818, g19766, g21556, I12861, g10165, g13782, g17575, g28137;
wire g11984, g16967, I22331, g32668, g32842, g17711, g7046, I32284, g20653, g27991, I33288;
wire g31802, g9631, g17327, g25060, g32489, g8389, I13329, I27388, g31857, g7446, g18200;
wire g29811, g23223, g7514, g19360, g11418, g34714, g8990, g12882, g9257, g22492, g25197;
wire g29343, g7003, I13539, g22303, I27777, g9817, g32559, g34315, g10475, I17932, g24138;
wire g32525, g32488, g11170, g34910, I29444, g8171, g10727, g7345, g7841, I12534, g20636;
wire I19384, g8787, g32558, g34202, g23084, g24636, g6826, g10222, g7191, g30055, g17606;
wire g20852, g32830, g23922, g23321, g32893, I18028, g21179, I24920, g26801, I24434, g29368;
wire g9751, g34070, g8281, g32544, g19629, g32865, g19451, g21178, g34590, g19472, g24963;
wire g20664, g34986, g32713, g7536, g9585, g8297, g10347, g21685, I16733, I12997, g28726;
wire g34384, g23953, g30067, g11401, g22840, g21654, I29977, g7858, g32610, g20576, g20585;
wire g23654, I12061, g32705, g34094, g13477, g8745, g28436, g8138, g8639, g24585, I22149;
wire g19071, g23800, I23711, g20554, g23417, g32679, g16322, g8791, g10351, g23936, g10372;
wire I23327, g25202, g19776, g19785, g34150, I32963, g16159, g22192, g20609, g28274, g15171;
wire g34877, g10175, I17723, g12082, g17390, g28593, g32678, g13022, g7522, g23334, g25055;
wire g19147, g30019, g7115, g12107, g8808, g19754, g7315, g16158, g20608, g25111, g9669;
wire g19355, I12360, g25070, g32460, g32686, I22343, g24115, g32939, I18903, g30018, g32383;
wire g19950, g14063, g19370, I19917, I14046, I17148, g16656, g9772, I26638, g20921, g12345;
wire I16476, g14790, g20052, g23964, I23303, g32938, g28034, g33533, g29310, g16680, g24052;
wire I17104, g12940, g17522, g21423, g12399, g9743, I16555, g23423, g8201, g9890, g13305;
wire g6827, g14873, g23216, g11900, g19996, g29379, g29925, g13809, I23381, I15036, g8449;
wire g12804, g9011, g19367, g19394, I12451, g6846, g9856, g8575, g13036, g32875, g30917;
wire I14827, g11560, g13101, g14209, g7880, g13177, g34917, g8715, g20674, g7595, g23543;
wire g6803, g16966, g7537, g24184, I18845, I32921, g16631, g14208, I18262, g29944, g22904;
wire g23000, I26578, g23908, g17326, g32837, g31856, I13206, g8833, g30077, g9992, g20732;
wire g23569, g25196, g10542, I31610, I23390, g13064, g24732, g14453, g7017, I30992, g7243;
wire g19446, g34597, I12776, I13759, I18191, g23568, I33255, I33189, g8584, g8539, g23242;
wire I32973, I29571, g34689, I33270, g34923, g9863, I12355, g16289, g9480, I17228, g6994;
wire g21123, g18100, g34688, g9713, g10607, g12833, g22847, g16309, I12950, g23814, g10320;
wire g32617, g28575, g32470, g10073, I18832, I31686, g7328, g32915, g10274, g29765, g10530;
wire g7542, I12858, g28711, g13009, g16308, g9569, g13665, g27004, g30102, g8362, I13744;
wire g31831, g32201, g24013, I33030, I12151, g10122, g6816, I12172, g17183, g17673, g17847;
wire I26430, g13008, g15656, I21483, g20329, I33267, g8052, I18861, g21293, g20207, g23230;
wire g15680, g20539, g25001, g17062, g20005, g13485, g20328, g32595, g32467, g32494, g19902;
wire g24005, g17509, g14034, g19957, g16816, g20538, g9688, g28606, g6847, g13555, g18882;
wire g32623, g18991, I28897, g19739, I25391, g9976, g17508, g29317, g10153, g23841, I22096;
wire g23992, g32782, g23391, g19146, g19738, g33080, g21510, g23510, g10409, g16752, I21757;
wire I33218, I25579, g16954, g29129, g22213, g19699, g8504, g34511, g10136, g16643, g10408;
wire g9000, g32822, g13074, I24191, g29128, g14635, I12227, g13239, g19698, g9326, I15238;
wire g12951, g25157, g23578, g8070, g13594, I16438, g23014, I25586, g8470, g20100, g7512;
wire g34660, I30983, g9760, g20771, g22311, g24100, g26054, g7490, I15382, I14647, g25231;
wire g7166, g20235, g19427, I26130, g11941, g19366, I17857, g32853, g24683, g33736, g11519;
wire I14999, g16195, g34480, g16489, g34916, g13675, I20861, g32589, g7456, g15224, g7148;
wire g6817, g7649, g22592, g22756, g16525, g15571, g26942, g9924, g10474, g32588, g32524;
wire g9220, g31843, g32836, g33696, g30076, g30085, g7851, I33075, g9779, g26655, g13637;
wire g20515, g34307, g23041, I20388, g32477, I18360, g21275, g24515, I31494, g24991, I12120;
wire g10109, g30054, g21430, g27163, g34596, g8406, g17756, I27738, g23430, g23746, g23493;
wire g7964, g7260, g8635, g24407, g34243, g29697, g9977, g19481, g10108, I14932, g29995;
wire I33037, g34431, g12012, g32118, g15816, g8766, g18940, g8087, I31782, g32864, g23237;
wire I19734, g7063, g10606, g21340, g32749, g32616, g23340, g23983, I22128, g34773, g9051;
wire g23684, g25480, g34942, g32748, I15577, g8748, g11215, g19127, g9451, g28326, I32991;
wire I14505, I33155, g13215, g26131, g34156, g13729, g25550, g20441, g20584, g32704, I21047;
wire g10381, g28040, g33708, I33170, g19490, g25287, g34670, I29939, g9999, I17128, g23517;
wire g33258, g32809, g32900, g25307, g32466, g7118, g7619, g16124, I19487, g19376, g19385;
wire I17626, g17413, g9103, g32808, I26952, g24759, I18071, g19980, g25243, g34839, g17691;
wire g20114, g16686, g34930, g11349, g34993, g12946, g15842, g32560, g20435, g8373, I15906;
wire g24114, g8091, I33167, g6772, g29498, g24082, I15284, g16030, g7393, g13906, g10390;
wire g21362, g24107, g32642, g9732, g23362, g34131, g29056, g22928, g9753, I26516, g23523;
wire g31810, g8283, g25773, I27481, g18833, g31657, g7971, g13304, I20447, I28582, I18825;
wire I18370, g24744, I31477, g29080, g7686, g33375, g8407, g17929, g9072, g25156, I29218;
wire g8920, g8059, g32733, I33119, g14192, I18858, g9472, g19931, g25180, g6856, I12572;
wire g15830, g17583, g8718, I18151, g34210, g32874, I28925, g9443, g21727, I22512, g20652;
wire g28508, g32630, g7121, g23863, g32693, I31616, g21222, I23396, g7670, g23222, I18367;
wire g26187, g29342, g9316, g25930, g7625, g32665, I31748, I13473, g19520, g6992, g12760;
wire g9434, g13138, g17787, g7232, g10553, g25838, I27784, I15636, I33276, I33285, g18947;
wire I27385, g30039, g30306, g25131, I33053, g15705, g26937, g17302, g32892, g23347, g24135;
wire g32476, g32485, g33459, I31466, g7909, g30038, g23253, I12103, g11852, g17743, g9681;
wire I22499, g10040, I22316, g32555, I18446, g14536, g19860, g33458, g7519, g24361, g11963;
wire g25557, g32570, g32712, g25210, g32914, I25351, g9914, I20355, g33918, g23236, g20500;
wire g10621, g34677, g29365, g14252, I22989, g13664, g20049, g23952, g23351, g32907, I31642;
wire g33079, g24049, I14896, g29960, g21175, g22881, g23821, g10564, g15938, g16075, g9413;
wire g19659, g14564, g24048, I11682, g11576, I33064, I25790, I17989, g20004, g13484, g32567;
wire g32594, g19658, g23264, g25286, g16623, g10183, I15609, g7586, g23516, g25039, I28548;
wire g10397, g6976, g14183, g14673, g11609, g9820, g16782, g12903, g20613, I21787, I22461;
wire g31817, g13312, I18301, g32941, g32382, g11608, g19644, g10509, I18120, g32519, I22031;
wire I27546, g32185, g18421, g14509, I15921, g32675, g8388, I23357, g20273, g20106, g12563;
wire g20605, g21422, I26409, g30217, g8216, g10851, I12089, g10872, g9601, g23422, g32518;
wire I16328, g24106, g24605, I14050, g29043, I16538, g13745, g32637, g31656, I20318, g17249;
wire I28002, g32935, g24463, I21769, I17650, I28128, g20033, g31823, I32613, g32883, g17248;
wire I30641, I31555, I14742, g19411, g19527, g17710, g24033, I17198, g12845, g27990, g16853;
wire I12497, g23542, g9581, g23021, g23453, g10213, I32947, g12899, g21726, g16589, g25169;
wire g29955, g9060, I32106, g23913, g15915, g9460, g24795, g29970, g7659, g12898, g22647;
wire g17778, g16588, g25168, g23614, g25410, g18829, I12987, I15732, g8741, g10047, I32812;
wire g19503, g29878, g15277, g21607, g22999, g23607, g21905, g14205, g26654, g20514, I25530;
wire g32501, g32729, g18828, g31631, g10311, g23320, g23905, g9739, g32577, g33631, I14730;
wire g18946, g29171, g21274, g14912, g30321, g23274, g20507, g23530, g22998, g27832, I32234;
wire g34922, I24281, g26936, g15595, g32728, g21346, g25015, g6977, I20957, g19714, I13240;
wire g7275, g22182, g29967, g29994, g34531, g9995, I12644, I11903, g23565, g10072, g32438;
wire I14690, g8883, g7615, g12440, g27573, I20562, g25556, g24163, I33176, g7174, g19979;
wire g16748, g7374, g12861, g17651, g17672, g34676, g8217, I16515, I17471, g9390, g21292;
wire g11214, g32906, g7985, g16285, g8466, I19762, g22449, g34654, g20541, I12855, g16305;
wire g10350, g13329, g16053, g9501, g6999, g16809, g21409, g22897, g7239, I12411, g23409;
wire g8165, g32622, g8571, g8365, I26381, g24789, g32566, g19741, I30537, g29079, g7380;
wire g21408, g10152, g7591, g23408, g8055, g10396, g20325, g24359, g19067, g20920, g20535;
wire I13990, g20434, g9704, g31816, g8133, g24920, g24535, I18376, g24358, I18297, I12503;
wire g17505, g17404, g10413, g8774, g32653, g19801, I32473, g17717, I17879, g34423, g15588;
wire I22886, g32138, I17970, I20895, g24121, I18888, g8396, g9250, g34587, I13718, g12997;
wire g10405, g32636, I23998, I32788, g32415, g14405, g19695, g8538, I12819, g29977, I12910;
wire g16874, g32852, g11235, I32535, I25327, g8509, g35002, g19526, g16630, g16693, g26814;
wire g34543, I22425, g24173, g32963, g22148, g7515, g12871, g29353, I12070, I22458, g23537;
wire g9568, g31842, g32664, g30569, I16345, g8418, I19772, g34569, g22646, I22918, g17433;
wire I25606, g8290, I17425, g18903, g30568, g23283, g19866, g11991, I17919, g13414, I22444;
wire g23492, g25423, g23303, I31622, g32576, g24134, g8093, g32484, g34242, g24029, g33424;
wire I11701, g10113, g17811, g17646, I11777, g20506, I28199, I25750, g20028, I12067, I32173;
wire g32554, I18089, g24506, I20385, g7750, g24028, I24784, g34123, g16712, g26841, g32609;
wire g21381, I27735, I29239, g31830, g23982, g10357, g26510, g14357, g34772, I12735, g8181;
wire g28779, g32608, g8381, g19689, g7040, g25117, I16135, g25000, g8685, g7440, g8700;
wire g28081, g32921, g33713, g8397, g19688, g9626, g8021, g16594, g26835, g13584, g18990;
wire g32745, I29185, g22896, I18700, g23840, g15733, g32799, g18898, g23390, g32813, g22228;
wire g6820, g33705, g25242, g7666, I17159, g20649, I17125, I22561, I23149, g31189, g34992;
wire I17901, g34391, g32798, I22353, g28380, g20240, I23387, g32973, I30904, g34510, g22716;
wire g23192, g16675, g20648, g10881, I17783, g20903, g32805, g13082, g32674, g24648, g7528;
wire g12859, g13107, g34579, g7648, g26615, g12950, g20604, g9683, g23522, g18832, I13360;
wire g24604, g30578, g33460, g33686, g19885, g26720, g7655, g11744, g20770, I26508, g9778;
wire I14271, g20563, g27996, g32732, g24770, g8631, g25230, g32934, g24981, I24089, g11849;
wire I16613, g17582, g12996, g10027, g23483, I18060, I23369, g14662, g8301, g19763, g25265;
wire I32240, g29976, g12844, g7410, g11398, g23862, g12367, g32692, g32761, I32648, g18926;
wire I18855, I11629, g11652, g9661, g13141, g29374, g20767, g26340, g21326, g18099, I18411;
wire g30116, I14650, g33875, I24497, g10710, g20899, I12300, g10003, g23948, I32770, g18098;
wire g10204, I29438, g21904, g14204, g16577, g20633, g23904, I16371, g31837, g14779, g21252;
wire I22289, g32329, g29669, g34275, g19480, g23252, g17603, g20191, g34430, g17742, g32539;
wire g10081, g17096, I18894, g6995, g7618, g8441, g22857, I22571, I11785, g7235, g7343;
wire I14365, g30237, I16795, g25007, g32538, g24718, I32794, g14786, g29195, g9484, g30983;
wire g9439, g17681, g7566, g6840, g8673, g16349, g34983, g18997, g10356, g33455, g21183;
wire g21673, g7693, g11833, g17429, g7134, g21397, g23847, g13049, g10380, g30142, g18061;
wire g16284, g19431, g34142, g25116, g17428, I22816, g7548, g11048, g8669, g10090, g20573;
wire g10233, g20247, g29893, I24060, g16622, g23509, g10182, g28620, I21959, g20389, g8058;
wire I14708, I28458, I29139, g8531, g19773, g24389, g8458, g24045, g12902, g20612, g23508;
wire I16163, I20870, g32771, g8743, g20388, g20324, g8890, I23378, g29713, g24099, g24388;
wire g20701, g20777, g20534, g22317, g31623, g32683, I17976, g25465, g19670, g24534, g8505;
wire g20272, g34130, g24098, g14331, g12738, I19863, g9616, g17504, I16541, g8011, g25340;
wire g25035, I17374, g8411, g8734, g19734, g13106, g27698, g29042, g13605, g10897, I33214;
wire I20867, I27314, g6954, g19930, g6810, g9527, I14069, g11812, g7202, I16724, g10404;
wire I12314, g13463, g31822, g32515, I31539, g32882, I14602, I15033, g19694, g7908, I32388;
wire g24032, g22626, I21802, I16829, g25517, g11033, g11371, I16535, g18911, g23452, g10026;
wire g32407, g9546, g13033, g21205, g11234, g10212, I14970, g29939, g17128, g7518, I17668;
wire I20819, I22525, I22488, I17842, I20910, g16963, g23912, I17392, g34222, g9970, g24061;
wire I29585, g29093, g34437, g20766, I26929, g8080, I18526, g31853, g19502, g8480, g19210;
wire g17533, g25193, g8713, g21051, g7593, I17488, g15348, g19618, g19443, I14967, g12895;
wire I12773, g16585, g13514, g25523, g31836, g32441, g32584, I32997, g24360, g29219, g15566;
wire g20447, g14149, g10387, g16609, g19469, I28336, g10620, g17737, g22856, g29218, g22995;
wire g32759, g16200, I33235, g23350, g25006, g32725, g24162, I32766, g7933, g16608, g19468;
wire g9617, g23820, g34952, g34351, g13012, g32758, g7521, I32871, g25222, g7050, g20629;
wire g23152, I12930, I13699, g9516, I21002, g20451, g21396, g31616, I14079, g30063, I22124;
wire g9771, I29973, g26834, g20911, I16028, g10369, g32744, I31515, g24911, g19677, I18280;
wire g12490, g17512, I17679, g21413, g9299, I15788, g23413, g27956, g32849, g9547, g10368;
wire g32940, g7379, g8400, g11724, I17188, g31809, I12487, g11325, g20071, g32848, g9892;
wire g24071, g11829, g12889, g11920, I11632, g20591, g25781, g10412, g20776, g20785, g31808;
wire g32652, g32804, g14412, g7289, I12618, g12888, g26614, g10133, g20147, I17938, g34209;
wire g7835, g24147, g10229, I18066, g12181, g26607, g17499, g22989, g23929, g17316, g11344;
wire g34208, I14158, g19410, g24825, g22722, g17498, g22988, g8183, g23020, I15682, g23928;
wire g8608, I18885, g30021, I32071, g19479, g19666, g6782, g25264, g16692, g25790, I29013;
wire g25137, g9340, I13715, g17056, I29214, g11291, I32591, g24172, g23046, g32962, g9478;
wire I14823, g19478, g24996, g17611, g17722, g9907, g13173, g34913, g10582, I16755, I29207;
wire g14582, g33874, g9959, g7674, g8977, g24367, g24394, I16770, g32500, g34436, g9517;
wire g9690, g17432, g23787, I27677, g29170, g32833, g18957, g21282, g16214, g17271, I32950;
wire g23282, I26710, g7541, g10627, I25105, g34320, g27089, g10379, g23302, I25743, g31665;
wire g25209, g19580, g30593, g33665, g6998, g22199, g34530, g10112, g34593, g7132, g12546;
wire I22470, g10050, g27088, g18562, g34346, g10378, g25208, g30565, g7153, g7680, g8451;
wire g22198, g22529, g34122, g15799, I21831, g13506, g12088, g13028, g20446, g10386, g29194;
wire g9915, g12860, g22528, g6850, g14386, g23769, I11980, g22330, I13889, g25542, g7802;
wire g20059, g32613, g8146, g10096, g20025, g8346, g24059, g33454, g14096, g24025, g9214;
wire g17529, g20540, g12497, g30292, I16898, g23768, I12884, I22467, g20058, g24540, g33712;
wire I26356, I18307, g32947, g19531, g24058, g22869, g17528, g7558, g32605, g8696, g34409;
wire I21722, g22868, I16521, g17764, I12666, g10429, g11927, g23881, g10857, g32812, g25073;
wire g32463, g16100, I32446, g19676, g19685, g31239, g25274, g24044, g16771, g34408, I22419;
wire g19373, g26575, g10428, g32951, g32972, g16235, g32033, I32059, g8508, g19654, I31361;
wire g9402, g9824, g8944, g8240, g18661, g20902, g18895, g19800, I18341, g19417, g21662;
wire g24377, g7092, I31500, g24120, g23027, g32795, g25034, I23342, g17709, g33382, I12580;
wire g8443, g19334, g20146, g20738, I18180, g25641, g20562, g9590, g21249, I15981, g24146;
wire g6986, g23249, I14687, g11770, I21199, I30998, g20699, g16515, g10504, g11981, g9657;
wire g12968, g17471, g25153, I26448, g8316, g17087, g23482, I25552, g32514, I18734, g24699;
wire g21248, g14504, g19762, g23248, g19964, I22589, g20698, g27527, g25409, g34575, I25779;
wire g32507, g9556, I18839, g23003, g8565, g21204, g33637, g29177, g30327, g33935, g34711;
wire g12870, I11860, g25136, g34327, I18667, I18694, g32421, I23330, I23393, g10129, I29441;
wire g11845, g9064, I18131, g8681, g10002, I25786, g10057, g9899, I32645, g7262, g24366;
wire g20632, I15633, I32699, I33273, g30606, g8697, I33106, I14668, I25356, g19543, g30303;
wire g8914, I19796, g17602, g12867, g12894, I17401, g16584, g17774, g23647, g18889, g17955;
wire g18980, g32541, g7623, g10323, g23945, g16206, I25380, g18095, g23356, g32473, I31463;
wire g19908, g22171, g13191, g26840, g20661, I12654, g21380, g10533, g20547, g23999, g32789;
wire g18888, g23380, g33729, I18443, g19569, I14424, I14016, I17118, g16725, I22748, g13521;
wire g22994, g34982, g32788, g32724, g19747, g23233, g21182, g6789, g11832, g23182, g20715;
wire g23651, g32829, g28080, g32920, I18469, g32535, g25327, g32434, I14830, I21258, g24481;
wire I14893, g25109, g12818, g20551, g20572, g9194, g32828, g18931, g6987, g32946, g10232;
wire I17276, g7285, g11861, g22919, g16744, I17704, g12978, g14232, g9731, g23331, I13968;
wire I32547, g19751, I24839, g9489, g19772, g25283, g34840, g20127, I22177, g23449, g26483;
wire g28753, g9557, g13926, g24127, g13045, g10261, I17808, g9071, g26862, g11388, g23897;
wire g13099, g11324, g23448, g23961, g32682, g24490, I14705, g19638, I17101, g34192, I21810;
wire I16629, g16652, g17010, g23505, I27543, g26326, g8922, g20385, I14679, g13251, I23375;
wire g13272, g19416, g20103, g7424, g24376, g24385, g34522, g7809, I18143, g24103, g23026;
wire g18088, g24980, I16246, I30971, I12117, g24095, g26702, g17599, I12000, g25174, g28696;
wire g31653, g6991, g33653, I14939, g7231, g20671, I17733, g27018, g31138, g32760, g17086;
wire g24181, g7523, g19579, g22159, g29941, g13140, g7643, I21792, I12568, g12018, I22009;
wire g34553, g10499, I22665, I13581, I18168, I24278, I14267, g32506, g8784, I31724, g33636;
wire g29185, I32956, g30326, g21723, g29092, I32297, g34949, g10498, I32103, g34326, g13061;
wire I31829, I18479, g31852, g6959, I31535, g30040, I13202, g19586, I12123, g17125, g17532;
wire g27402, g34536, I17166, g28161, g7634, g15758, g21387, I22485, I29221, g23433, I28419;
wire I13979, I32824, g24426, g8479, g20190, g22144, I24038, g23620, g28709, g10080, I17008;
wire I32671, g8840, g9212, g12866, I21918, I17892, g21343, I26925, g8390, g32927, g15345;
wire g14432, g17680, g17144, g26634, g26851, g11447, g7926, I15162, g20546, g20089, g23971;
wire I26378, g19720, g20211, I25369, g24089, I19851, g27597, g21369, I33291, g12077, g32649;
wire g25553, g20088, I27391, g8356, I20937, g9229, I13094, g14753, I33173, g24088, g19493;
wire g24024, g14342, g34673, g34847, g31609, g29215, g10031, g32648, g32491, g32903, g25326;
wire g14031, g9822, g10199, I11801, I14455, g16605, g11472, I27579, I29371, g12923, g31608;
wire g18527, g20497, g32604, g34062, I28588, g32755, I30959, g10198, g12300, g11911, g16812;
wire g21412, g32770, g34933, g14198, g32563, I32089, I33134, g13246, g20700, g20659, g34851;
wire g20625, g10393, g24126, g24625, g14330, g24987, g8954, g7543, g31799, g23896, g25564;
wire g8363, g18894, g31813, g21228, g33799, g10365, g22224, g33813, g8032, g19517, g23228;
wire I18373, g29906, g29348, g16795, g10960, I17675, g23011, g31798, g32767, g32794, I14623;
wire g11147, g11754, I17154, I23680, g25183, g32899, g7534, g31805, g17224, g16514, g12885;
wire g22495, g17308, g23582, g32633, g32898, I32659, g15048, g9620, g9462, I23336, I19756;
wire g19362, g7927, g34574, g32719, I12041, g20060, g34047, g18979, g19523, g24060, g8912;
wire I16120, g33934, g10708, g20197, g6928, I12746, g21379, g34311, I12493, g22976, g22985;
wire g32718, g32521, g10087, g23925, g8357, g18978, g7946, g7660, g29653, I22729, g26820;
wire g21050, g20527, I13597, g11367, g28918, g32832, I20321, g23378, g13394, I31491, g33761;
wire g24527, g7903, g30072, g17687, I31604, g28079, g10043, I13280, g7513, g26731, g34592;
wire I11688, I16698, g29333, g16473, I31770, g32861, g9842, g23944, g32573, g18094, g31013;
wire I14589, g25213, g19437, g20503, g9298, g28598, I18909, g9392, g32926, I32855, g7178;
wire g7436, I14836, g8626, g21681, g29963, g16724, g22842, g23681, I18117, g32612, g16325;
wire g18877, I23309, g25452, g15371, g25047, g32099, g10375, I21288, g34820, g16920, g20714;
wire g20450, g23429, g32701, g12076, g7335, g7831, I14119, g32777, g32534, g12721, g34152;
wire g20707, g21428, I22622, g20910, g34846, g23793, g12054, g17392, g19600, g10337, g24819;
wire g19781, g17489, I24334, g20496, g7805, g7916, g25051, g25072, g24818, g32462, I14749;
wire g24979, g21690, g22830, g19952, g24055, g7749, g19351, I12523, g23549, g27773, g20070;
wire g20978, g24111, g28656, g9708, g24070, g24978, g34691, g29312, g20590, g22544, g22865;
wire g23548, g8778, g29115, g7947, I20216, g24986, I14305, g9252, I26880, g23504, g13902;
wire g13301, g31771, g19264, g18917, g19790, g20384, g12180, g9958, g29921, g13120, I18293;
wire g24384, g25820, I26512, I17653, g20067, g32766, g6955, g29745, g24067, g24094, g11562;
wire g17713, I18265, g34929, g27930, I12437, g27993, g8075, g32871, g30020, g30928, g22189;
wire g8475, g26105, g9829, g12839, g6814, g12930, g7873, g26743, g26827, g34583, g7632;
wire g34928, g7095, I17636, g21057, g23002, g10079, g11290, g24150, g23057, I28594, g9911;
wire g7495, g14545, g7437, g17610, I27253, I30995, g12838, g23128, I20569, I17852, g10078;
wire g21245, g24019, g17189, g23245, I13287, g26769, g8526, g19208, g20695, I20747, I31701;
wire g21299, g30113, g9733, g10086, g23323, g23299, g9974, I32067, g17188, I11721, g17124;
wire g17678, g34787, g26803, g12487, g20526, I22576, I28185, I18835, I13054, g24526, g19542;
wire g30302, g7752, I16181, g18102, g8439, g9073, g32629, g34302, I26989, I32150, g30105;
wire g6836, g7917, I14630, g27279, g32472, g10159, g34827, g10532, g32628, g17093, g6918;
wire g32911, g14125, g15344, g10158, g11403, g11547, g13895, g20917, I33140, I28883, g23232;
wire g24866, g19905, I12790, I17609, g34769, I11655, g18876, g18885, g10353, g25046, g6993;
wire g10295, g8919, g21697, g29013, I29981, g34768, g12039, g13715, I22745, g29214, g27038;
wire g9206, g32591, I15572, g23995, g32776, g32785, I30989, g19565, g24077, g20706, I11734;
wire g23880, g12038, g20597, I21042, g32754, I14570, g33435, g25282, I21189, g14336, g27187;
wire g7296, g23512, g8616, g28752, g20923, g27975, g32859, g32825, g32950, g28954, g26710;
wire g18660, g20624, g22455, g12975, g7532, I13694, I16024, g32858, g33744, g7553, g8404;
wire g15506, g31849, g8647, g14631, g10364, g19409, I14567, g12143, g20102, g16767, g20157;
wire g25640, g12937, g28669, g26081, g8764, g22201, g24102, g23445, g31848, g18916, g24157;
wire g32844, g9898, g33848, g28260, g17617, g18550, g25768, g25803, g31141, I26960, g22075;
wire g18314, g33652, g18287, g27410, g16633, g30248, g34482, g23498, g28489, g26356, g18307;
wire g29771, g30003, g34710, g16191, g22623, g21989, g30204, g13671, g26826, g27666, I31246;
wire g18721, g22037, g25881, g26380, g33263, g18596, g32420, g28488, g27363, g23056, g27217;
wire g29683, g18243, g33332, I17692, g21988, g26090, g21924, g28558, g18431, g26233, I31071;
wire g26182, g26651, g12015, g34081, g27486, g31962, g24763, g33406, g18269, g33361, g15903;
wire g18773, I31147, g18341, g29515, g29882, g18268, g29991, g21753, g31500, g18156, g18655;
wire g33500, g24660, g33833, g32203, g18180, g26513, g17418, I27409, g34999, g18670, g34380;
wire g25482, g32044, I24684, g16612, g21736, g11546, g21887, g30233, g18734, I31151, g16324;
wire I31172, g18335, g16701, g22589, g32281, g34182, g28255, g16534, g28679, g11024, g16098;
wire I13937, g18993, g24550, g32301, g14643, g24314, g22588, g21843, g32120, g24287, g28124;
wire g15794, g18667, g18694, g12179, g24307, g29584, g27178, g21764, g11497, g18131, g29206;
wire g13497, g28686, g32146, g28939, g24721, g22119, g21869, g27186, g31273, g34513, g21960;
wire g27676, g27685, g15633, g33106, g18487, g27373, g29759, g22118, g32290, g11126, g12186;
wire g28267, g17401, g21868, g18619, g18502, g22022, g34961, g12953, g18557, g33812, g18210;
wire g29758, g17119, g33463, I31227, g18618, g18443, g24773, g21709, g18279, g30026, g33371;
wire g30212, g16766, g26387, g27334, g34212, g28219, g21708, g18278, I16111, g26148, g23708;
wire g16871, g29345, g22053, g23471, g26097, g18469, g24670, g33795, g28218, g29940, g26104;
wire g18286, g22900, g27762, g15861, g8690, g27964, g18468, g25331, g18306, g12762, g22036;
wire g25449, g13060, g31514, g32403, g27216, g33514, g22101, g24930, g29652, g29804, g17809;
wire I31281, g28160, g15612, g25448, g18815, g30149, g25961, I27381, g33507, I31301, g20131;
wire g15701, g10705, g18601, g13411, g18187, g18677, g14610, g28455, g33421, g21810, g17177;
wire g21774, g29332, g23657, g28617, g34097, g21955, g23774, g22064, I24600, I31146, g25026;
wire g34104, g27117, g21879, g34811, g21970, g18143, g24502, g28201, g19536, g19948, g29962;
wire g21878, I16695, g32127, g31541, g24618, g26229, g33473, g18169, g21886, g27568, g18791;
wire g31789, g28467, g28494, g33789, g21792, g16591, g22009, g22665, g18168, g18410, g21967;
wire g21994, g31788, g33724, g32376, g19564, g33359, g25149, g17693, g22008, g32103, g24286;
wire g18479, g18666, g33829, g18363, g32095, g18217, g33434, g24306, g33358, g25148, g11496;
wire g15871, g18478, g30133, g33828, g28352, g11111, g14875, g34133, g21919, g30229, g25104;
wire g11978, g26310, g23919, g32181, g33121, g18486, g27230, g27293, g29613, g28266, g19062;
wire g33344, g14218, g21918, g30228, g26379, g18556, g25971, g24187, g34228, g30011, g27265;
wire I31226, g16844, g18580, g26050, g27416, g26378, g13384, g29605, g18223, g23599, g27992;
wire g22074, g27391, g24143, g25368, g27510, g34582, g32190, g26096, g29951, g18110, g34310;
wire g25850, g15911, g28588, g28524, I31127, g18321, g24884, g30925, g21817, g11019, g18179;
wire g13019, g18531, g30112, g28477, g33760, g24410, g32089, g25229, g30050, g29795, g34112;
wire g11018, g18178, g18740, g26857, g34050, g21977, g22092, g23532, g23901, g34378, g16025;
wire g33506, I24530, g32088, g24666, g22518, g21783, I31297, g24217, g18186, g15785, g18676;
wire g18685, g34386, g18373, g29514, g24015, g30096, g22637, g17176, g34742, g28616, g34096;
wire g18654, g16203, g28313, g27116, I27509, g21823, g27615, g18800, g15859, I31181, g18417;
wire g24556, g28285, g34681, I27508, g15858, g27041, g32126, g18334, g27275, g19756, g33927;
wire g28254, g27430, g34857, g10822, g24223, g27493, g16957, g25959, g30730, g25925, g28466;
wire g25112, g21966, g18762, g25050, g20084, g32339, g31240, g19350, g34765, g27340, g27035;
wire g18423, g29789, g32338, g33491, g33903, g24922, g26129, g18216, g24321, g16699, g27684;
wire g28642, g18587, g25096, g29788, g26128, g14589, g29535, I31211, g27517, g10588, g18909;
wire g32197, g18543, g26323, g24186, g14588, g24676, I16721, g18117, g16427, g25802, g22083;
wire g32411, g23023, g19691, g24654, g28630, g29344, g18569, g30002, g27130, g30057, g22622;
wire g18568, g18747, g25765, g27362, g31990, g33899, g18242, g10616, g27523, g30245, I31126;
wire g26232, g33898, g21816, g18123, g18814, g33719, g24762, g10704, g34533, g18751, g18807;
wire g21976, g21985, g15902, g18772, g28555, g33718, g34298, g28454, g33521, g18974, g26261;
wire g32315, g24423, g21752, g27727, I31296, g18639, g28570, g28712, g21954, g27222, g29760;
wire g33832, g18230, g29029, g17139, g18293, g17653, g15738, g18638, g27437, g33440, g32055;
wire g17138, g18265, g25129, g15699, g30232, g32111, g18416, g25057, g32070, g33861, g28239;
wire g25128, g17636, g11916, g33247, g28567, I31197, g27347, g18992, g18391, g24908, g28238;
wire g21842, g18510, g30261, g23392, g24569, g25323, g31324, g33099, g13287, g27600, g10733;
wire g18579, g31777, g33701, g24747, g32067, g21559, g31272, I16618, g15632, g28185, g10874;
wire g18578, g25775, g23424, g27351, g27372, g19768, g14874, g16671, g21558, g27821, g32150;
wire g28154, g18586, g29649, g33462, g21830, g26611, g20751, g10665, g28637, g18442, g32019;
wire g24772, g29648, g27264, g22115, g27137, g21865, g31140, g32196, g13942, g24639, g32018;
wire g26271, g29604, g30316, g21713, g34499, g24230, g13156, g18116, g24293, g18615, g22052;
wire g10476, g24638, g29770, g16190, g29563, I31202, g34498, g18720, g26753, I31257, g25880;
wire g14555, g24416, g16520, g21705, g30056, g18275, g26145, I31111, g18430, g18746, g27209;
wire g32402, g18493, g33871, g30080, g28215, g26650, g34080, g16211, g27208, g18465, g29767;
wire g29794, g21188, g33360, g18237, g29845, g23188, I16143, g28439, g18340, g29899, g29990;
wire g21939, g25831, g15784, g18806, g18684, g26393, g14567, g24835, g29633, I31067, g24014;
wire g15103, g34753, g21938, g18142, g34342, g30145, g30031, g27614, g32256, g18517, g27436;
wire g30199, g29718, g29521, g16700, g31220, g33472, g16126, g28284, g10675, g25989, g27073;
wire g30198, g32300, g14185, g25056, g28304, g33911, g34198, g26161, g34529, g21875, g25988;
wire I31196, g25924, g27346, g34528, g17692, g18130, g34696, g18193, g22013, g32157, g34393;
wire g26259, I24508, g18362, g23218, g29861, g29573, g33071, g21837, g34764, g22329, g10883;
wire g18165, g23837, g18523, g26087, g27034, g13306, g31776, g34365, g26258, g19651, g33785;
wire g29926, g34869, g28139, g22005, g31147, g28653, g13038, g27292, g29612, g24465, g12641;
wire g22538, g27153, g33355, g29324, g34868, g7396, g25031, g30161, g18475, g33859, g26244;
wire g29534, g33370, g24983, g27409, g16855, g18727, g28415, g24684, g28333, g33858, g34709;
wire g18222, g10501, g16870, g27136, g27408, g27635, g21915, g30225, g31151, g18437, g24142;
wire I31001, g31996, g34225, I31077, g26602, g30258, g11937, g15860, g34087, g23201, g33844;
wire g33367, I31256, g18703, g22100, g18347, g19717, g14438, g30043, g18253, g25132, g30244;
wire g26171, g15700, I24051, g18600, g20193, g18781, g28585, g24193, g28484, g33420, g30069;
wire g29766, g18236, g21782, g17771, g20165, g34069, g21984, I31102, g26994, g27474, g28554;
wire I31157, g18351, g18372, g24523, g32314, g29871, g33446, g27711, g16707, g21419, g32287;
wire g34774, g18175, g18821, g34955, g27327, g34375, g16202, g28312, g28200, g32307, g14566;
wire g32085, I31066, g29360, g21822, g22515, I31231, g22991, g27537, g28115, g31540, g25087;
wire g32054, g24475, g7685, g18264, g18790, g18137, I27513, g18516, g34337, g24727, g34171;
wire g16590, g24222, g16986, g27303, g11223, g25043, g32269, g21853, g28799, g26079, g34967;
wire g28813, g29629, g32341, g31281, g15870, g26078, g32156, g25069, g24703, g31301, g18209;
wire g29628, g33902, g21836, g31120, g32180, g23836, g26086, g28674, g13321, g25068, g25955;
wire g30919, g18208, g16801, g16735, g23401, g25879, g24600, g25970, g31146, g30010, g30918;
wire g32335, g11178, g11740, g18542, I18803, g18453, g29591, g29785, g31290, g22114, g26159;
wire g26125, g21864, g34079, g22082, g27390, g18726, g26977, g30599, g22107, g30078, g21749;
wire g26158, g17725, g26783, I31287, g18614, g28692, g28761, g34078, g18436, g25967, g30598;
wire g14585, g29859, I31307, I31076, g30086, g21748, g15707, g15819, g18607, g34086, g18320;
wire g24790, g21276, g21285, g26295, g29858, g21704, g18274, g22849, g33366, g27522, g26823;
wire g15818, g18530, g25459, g18593, g18346, g19716, g21809, g23254, g28214, g15111, g22848;
wire g18122, g23900, g34322, g14608, g15978, g18565, g26336, g30125, g18464, g21808, g29844;
wire g34532, g15590, g29367, g28539, g10921, g27483, g30158, g33403, g24422, I31341, g32278;
wire g27553, g18641, g18797, g25079, I31156, g18292, g16706, g31226, g32286, g34561, g16597;
wire g18153, g27326, g25078, g31481, g32039, g33715, g32306, g34295, g33481, g22135, g27536;
wire g18409, g27040, g25086, g21733, g10674, g18136, g18408, g18635, g24726, g27252, g24913;
wire g21874, g25817, g32187, g26289, g24436, g25159, g10732, g22049, g25125, g27564, g25901;
wire g26023, I31131, g34966, g31490, g10934, g24607, g25977, g26288, g33490, g19681, g24320;
wire g28235, g26571, g23166, g23009, g22048, g26308, g29203, g18164, g28683, g32143, g31784;
wire g34364, g33784, g31376, g31297, g27183, g33376, g27673, g22004, g23008, g33889, g11123;
wire g24464, I24027, g16885, g32169, g18575, g18474, g29902, g30289, g29377, g13807, g18711;
wire g32168, g32410, g28991, g13974, g18327, g24797, g30023, g21712, I24482, g18109, g27508;
wire g16763, g27634, g34309, g21914, g24292, g30224, g18537, I24710, g34224, g30308, g22106;
wire I24552, g29645, I24003, g17613, g34571, g18108, g14207, g21907, I31286, I13862, g15077;
wire g24409, g25966, I31306, g13265, g18283, g15706, g18606, g18492, g18303, g24408, g24635;
wire g34495, g22033, g27213, g18750, g31520, I31187, g33520, g18982, g18381, g34687, g21941;
wire g26842, I27429, g27452, g21382, g29632, g31211, g26195, g34752, g23675, g18174, g27311;
wire g18796, g28725, g32084, g32110, g16596, g28114, g25571, g33860, g32321, g16243, g29661;
wire g29547, g29895, g28107, g10683, g32179, g21935, g18390, g31497, g33497, g20109, g24327;
wire g21883, g32178, g15876, g24537, g11116, g20108, g34842, g18192, g22012, g26544, I27504;
wire I18620, g25816, g33700, g33126, g31987, g29551, g29572, g26713, I31217, g34489, g24283;
wire g18522, g27350, g18663, g24606, g25976, g24303, g16670, g27820, g34525, g28141, g34488;
wire g28652, g13493, g25374, g31943, I24505, g21729, g26610, g33339, g33943, g31296, g34558;
wire g16734, g23577, g18483, g24750, g32334, g21728, g33338, g28263, g16930, g23439, g11035;
wire g18553, g13035, g26270, g31969, g29784, g26124, g22920, g16667, g20174, g29376, g27413;
wire g34865, g16965, g18949, g31968, g18326, g24796, g11142, g27691, g17724, g29354, I27533;
wire g18536, g23349, g22121, g29888, g33855, g14206, g21906, g18702, g21348, g18757, g31527;
wire g23083, g23348, g15076, g33870, g33411, g33527, g26294, I31321, g16619, g30042, g18252;
wire g18621, g25559, g30255, g25488, g28833, g16618, g34679, g18564, g30188, g24192, g30124;
wire g16279, g34678, g27020, g31503, I18716, I31186, g33503, g24663, g33867, g17682, g34686;
wire g13523, g18183, g18673, g25865, g26218, g18397, g30030, g30267, g34093, g33450, g22760;
wire g22134, g27113, g32242, g18509, g22029, g31707, g34065, g33819, g33707, g18933, g33910;
wire g24553, g26160, g28273, g7696, g18508, g22028, g27302, g18634, g21333, g23415, g27357;
wire g25042, g31496, g33818, g24949, g33496, g19461, g27105, g24326, g30219, g17134, g21852;
wire g15839, g34875, g28812, g33111, g34219, g31070, g19145, g24536, g29860, g17506, g25124;
wire g15694, g15838, g21963, g24702, g34218, g24757, g31986, g19736, g24904, g28234, g32293;
wire I31216, g25939, g26277, g18213, g32265, g25030, g25938, g25093, g31067, g24564, g29625;
wire g29987, g19393, g16884, g18574, g23484, g18452, g18205, g31150, g23554, I31117, g18311;
wire g33801, g24673, g33735, g33877, I24582, g30915, g29943, g34470, g16666, g25875, g31019;
wire I18765, g29644, g29338, g30277, g13063, g31018, g32014, g29969, g30075, g26155, g14221;
wire g21921, g26822, I31242, g16486, g18592, g23921, g18756, g34075, g31526, g24634, g30595;
wire g33526, g24872, g29968, g21745, g18780, g12027, g14613, g27249, g21799, g29855, g17770;
wire g21813, g23799, g27482, g15815, g28541, g10947, g18350, I24603, g33402, g29870, g29527;
wire g27710, g21798, g34782, I27529, g18820, g26853, g28789, g21973, g32116, g27204, g33866;
wire g22899, g21805, g22990, I27528, g18152, g25915, g32041, g18396, g22633, g17767, g18731;
wire g30266, g28535, g15937, g25201, g22191, g16179, g29867, g29894, g19069, g21732, g16531;
wire g13542, g21934, g18413, g24912, g26119, g24311, g16178, g18691, g15884, g33689, g32340;
wire g29581, g32035, g31280, g17191, g17719, g21761, g29315, g27999, g26864, g26022, g13436;
wire g18405, g31300, g30167, g30194, g30589, I24690, I24549, g26749, g27090, g29202, g25782;
wire g32142, g13320, g26313, g28291, g29979, g34588, g22861, g27651, g34524, g33102, I31007;
wire g26276, g26285, g34401, g34477, g22045, g18583, g29590, g34119, g26254, g31066, g31231;
wire g29986, g22099, g27932, g27331, g30118, g24820, g26808, g16762, g20152, g22534, g29384;
wire g22098, g32193, I31116, g24846, g26101, g33876, g33885, g26177, g18113, g18787, g32165;
wire g24731, I31041, g18282, g34748, g27505, g27404, g31763, g18302, g33511, g15084, g18357;
wire g19545, g29877, g15110, g18105, g10724, g22032, g30254, g18743, g27212, g10829, I31237;
wire g21771, g10828, g18640, g18769, g22061, g30101, g30177, g29526, g17140, g26630, g34560;
wire g18768, g18803, g31480, I31142, g33480, g24929, g22871, g26166, g27723, g15654, g31314;
wire g28240, g27149, g30064, g17766, g27433, g27387, g15936, g25285, g29866, g27148, g21882;
wire g21991, g26485, g23991, g27097, g33721, g19656, g27104, g16751, g16807, g27646, g25900;
wire g34874, g23407, g33243, g28563, g25466, g19680, g33431, g16639, g26712, I17741, g18662;
wire g32175, g30166, g30009, g24302, g16638, g33269, g34665, g22472, g18890, g13492, g27369;
wire g24743, g30008, g18249, g33942, g33341, g18482, g14506, g29688, I31006, g29624, g14028;
wire g18248, g16841, g18710, g34476, g34485, g18552, g24640, g24769, g19631, g18204, I31222;
wire g27412, g34555, g18779, g22071, g24803, g33734, g30914, g21759, g15117, g23725, g18778;
wire g25874, g27229, g31993, g21758, g26176, g26092, g18786, g27228, g24881, I31347, g22859;
wire g26154, g30239, g17785, g25166, g31131, g18647, g34074, g30594, g18356, g29876, g29885;
wire g21744, g30238, g34567, I31600, g28440, g18826, g18380, g19571, g33487, g22172, g29854;
wire g21849, g21940, I31236, g15814, g31502, g28573, g25485, g33502, g29511, g31210, I31351;
wire g18233, g28247, g21848, g15807, g18182, g27310, g18651, g18672, g34382, g30185, g34519;
wire g17151, g21804, g34185, g27627, g25570, g27959, g28612, g34092, g30154, g28324, g24482;
wire g31278, g34518, g32274, g27050, g27958, g25907, g24710, g27378, I31137, g18331, I27364;
wire g24552, g33469, g28251, g30935, g28272, g31286, g32122, g18513, g21332, g18449, I26972;
wire g27386, g19752, g33468, g15841, g25567, g27096, g18448, g29550, g32034, g25238, g16806;
wire g29314, g22059, g21962, g18505, g21361, g22025, g18404, g24786, g33815, g32292, g10898;
wire g18717, g22058, g31187, g32153, g24647, g33677, g31975, g13252, g18212, g29596, g24945;
wire g10719, g16517, g21833, g30215, g32409, g14719, g34215, g30577, g34577, g25518, g27428;
wire g13564, g22044, g26304, g31143, I24709, I31021, g24998, g12730, g27765, g24651, g24672;
wire g14832, g29773, g27690, g16193, g27549, g31169, g11397, g18723, g25883, g28360, g22120;
wire g33884, g15116, g18149, g27548, g31168, g32164, g18433, g33410, g18387, g24331, g30083;
wire g13509, g27504, g18620, g18148, g21947, g30284, g34083, g34348, I31593, g33479, g34284;
wire g21605, I31346, g33363, g13508, g18104, g18811, g18646, I31122, g14612, g31478, g8234;
wire g31015, g18343, g24897, g29839, g30566, g33478, g24961, g21812, g17146, g34566, g28451;
wire g16222, g31486, g32327, g29667, g29838, g27129, g33486, g32109, g21951, g26852, g21972;
wire g27057, g19610, g18369, g24717, g27128, g28246, I31292, g32108, g30139, g18368, g34139;
wire g16703, g22632, g31223, g21795, g32283, g27323, g30138, g27299, g29619, g32303, g34138;
wire g11047, g18412, I31136, g11205, g13047, g27298, g29618, g19383, g34415, g18133, g23514;
wire g26484, g33110, g13912, g34333, g24723, g31321, g18229, g33922, g14061, g33531, g18228;
wire g24387, g26312, g34963, g26200, g32174, g21163, g21012, g28151, g18716, g31186, g33186;
wire g24646, g33676, g33373, g16516, g27697, g18582, g27995, g31654, g30576, g22127, g34585;
wire g34484, g18310, g29601, g31936, g33417, I31327, g21789, g26799, g29975, g34554, g18627;
wire g15863, g18379, g30200, g21788, g33334, g18112, g16422, g23724, g25852, g18378, g22103;
wire g34115, g21829, g29937, g14220, g21920, g23920, g22095, g16208, g25963, g28318, g18386;
wire g30921, g28227, g21828, g15703, g17784, g23828, g18603, g21946, g18742, g27445, g33423;
wire g29884, g23121, g24229, g34745, g27316, g24228, g18681, I31091, g24011, g32326, g29666;
wire g17181, g16614, g17671, g29363, g23682, g18802, g18429, g32040, g24716, I24680, g33909;
wire g34184, g18730, g15821, g27988, g18793, g18428, g24582, g33908, g28281, g16593, g12924;
wire g27432, g13020, g18765, g28301, g24310, g16122, g18690, g28739, g18549, g11046, g25921;
wire g13046, g26207, g24627, g29580, g21760, g20112, g31242, g22089, g27461, g33242, g18548;
wire g15873, g28645, I31192, g27342, g24378, g16641, g27145, g22088, g18504, g22024, g31123;
wire g32183, g19266, g33814, g28290, g32397, g13282, g27650, g29110, g25973, g18317, g33807;
wire g31974, g29321, g33639, g26241, g34214, g29531, g31230, g18129, g30207, g16635, g27696;
wire g34329, g27330, g27393, g28427, g24681, g29178, g29740, g30005, g22126, g18128, g21927;
wire g26100, g19588, g33416, g29685, I31326, g18245, g27132, g34538, g18626, g15913, g24730;
wire g31992, g18323, g33841, g18299, g18533, g28547, g33510, g24765, g18298, g27161, g30241;
wire I31252, g31579, g18775, g24549, g28226, g21755, g29334, g16474, g23755, g27259, g19749;
wire g32047, g33835, g9968, g21770, g32205, g21981, g22060, g10902, g18737, g27087, g28572;
wire g12259, g24504, g32311, g25207, g29762, g18232, g34771, g29964, g16537, g11027, g30235;
wire I18713, g25328, g11890, g24317, g15797, g18697, g27043, g32051, g16283, g29587, I31062;
wire g18261, g21767, g21794, g21845, g12043, g16303, g10290, g24002, g21990, g11003, g18512;
wire g23990, I27524, g33720, g19560, g29909, g27602, g31275, g34515, g34414, g28889, g31746;
wire g27375, g26206, g31493, g32350, g21719, g33493, g24323, g24299, g13778, g13081, g29569;
wire g21718, g33465, g31237, g10632, g24298, g33237, g32152, g18445, g24775, g29568, g29747;
wire g32396, g33340, g21832, g18499, g18316, g33684, g16840, g31142, g22055, g18498, g32413;
wire g19693, g22111, I31047, g21861, g34584, g22070, g13998, g31517, g26345, g28426, g33517;
wire g29751, g29807, I31311, g29772, g22590, g16192, g26849, g29974, g15711, g18611, g27459;
wire g21926, g18722, g26399, g25414, g25991, g23389, g29639, g15109, g26848, I16646, g26398;
wire g22384, g18432, I24705, g29638, I31051, g21701, I31072, g18271, g30082, g34114, g15108;
wire g21777, g34758, g26652, g31130, g22067, g22094, g34082, g30107, g21251, I24679, g33362;
wire g11449, g27545, g16483, g18753, g18461, g31523, g32020, g18342, g33523, g29841, g19914;
wire g29992, g27599, g34744, g18145, g29510, g32046, g18199, g22019, g27598, g18650, g18736;
wire g27086, g31475, g29579, g17150, I24030, g33475, g16536, g18198, g22018, g18529, g21997;
wire g32113, g34398, I31152, g33727, g24499, g29578, g33863, g19594, g29835, g34141, g16702;
wire g24316, g31222, g32282, g27817, g15796, g18696, g18330, g32302, g18393, g24498, g29586;
wire g16621, g12817, g21766, g26833, g26049, g30263, g32105, g28658, g18764, g20056, g18365;
wire g27158, g21871, g25107, g22457, g15840, g18132, g26048, g28339, g30135, g24722, g34135;
wire I18782, g7948, g29615, g16673, g18161, g34962, g19637, g26613, g18709, g22001, g22077;
wire g25848, g14190, g27336, g30049, g18259, g29746, g34500, g18225, g33351, g33372, g18708;
wire g28197, g25804, g18471, g33821, g26273, g30048, g22689, g18258, g16634, g20887, g23451;
wire g24199, g24650, g23220, g24887, g30004, I31046, g22624, g21911, g30221, g31790, g33264;
wire g31516, g24198, g33790, g33516, g29806, g29684, g18244, g26234, g22102, g24843, g33873;
wire g24330, g22157, g24393, I24075, I31282, g25962, g16213, g24764, g29517, I31302, I31357;
wire g21776, g21785, I27519, g18602, g18810, g15757, g18657, g22066, g18774, g7918, g18375;
wire g31209, g33422, g34106, g32248, g21754, I27518, g10625, g27309, g23754, g28714, g16047;
wire g25833, g14126, g16205, g27288, g28315, g33834, g31208, g32204, g21859, g21825, g21950;
wire g26514, g22876, g18337, g28202, g30033, g28257, g21858, g29362, g18171, g30234, g34371;
wire g24709, g31542, g31021, g29523, g23151, g28111, g14296, g21996, g24225, g15673, g18792;
wire g15847, g23996, g24708, g14644, g33913, g16592, g21844, g21394, g32356, g29475, g18459;
wire g18425, g33905, g33073, g12687, g25106, g26541, g34514, g15851, g15872, g18458, g19139;
wire g27374, g33530, g21420, g34507, g31122, g32182, g20069, g33122, g8530, I31027, I24524;
wire g33464, I16129, g20602, g28150, g16846, g18545, g25951, g26325, g24602, g25972, g18444;
wire g25033, g25371, g20375, g24657, g24774, g16731, g26829, g27669, g17480, g19333, g29347;
wire g18599, g22307, g22076, g22085, g26358, I27349, g23025, g27260, g32331, g31292, g26828;
wire g27668, g23540, g18598, g22054, g28695, g31153, g27392, g29600, g26121, g20171, g34541;
wire g17307, g15574, g33409, I24616, g29952, g27559, g29351, g27525, g27488, g18817, g15912;
wire g14581, g18322, g33408, I31081, g24967, g10707, g18159, g27558, g25507, g22942, g18125;
wire g18532, g26291, g30920, I24704, g19585, g14202, g16929, g18158, g14257, g21957, g18783;
wire g23957, g29516, g14496, g22670, g21739, I31356, g25163, g18561, g18656, g30121, g25012;
wire g18353, g18295, g21738, g10590, g17156, g17655, g18680, g18144, g18823, g34344, g21699;
wire g28706, g28597, I31182, g18336, g24545, g33474, g28256, g15820, g28689, g32149, g27042;
wire g33711, g30173, g34291, g31327, g27255, g28280, g22131, g29834, g33327, g34173, I24064;
wire g29208, g25788, g32148, g28624, g28300, g27270, g32097, I31331, g27678, g18631, g32104;
wire g7520, g18364, g32343, g31283, g27460, g27686, g25946, g31492, g24817, g30029, g33492;
wire g19674, g24322, g12939, g27030, g20977, g13299, g24532, g32369, g27267, g27294, g29614;
wire g30028, g28231, g24977, g34506, g16803, g31750, g29607, g18289, I31026, g29320, g33381;
wire I31212, g29073, g12065, g18309, g29530, g24656, g29593, g33091, g18288, g18224, g21715;
wire g22039, g29346, g25173, g24295, g18571, g18308, g24680, g27219, g32412, g24144, g33796;
wire g19692, I24555, g29565, g26604, g17469, g13737, g22038, g23551, g23572, g10917, g12219;
wire g27218, g30927, g18495, g33840, g29641, g29797, g16662, g13697, g28660, g18816, g32011;
wire g27160, g10706, g15113, g19207, g18687, g28456, I31097, g17601, g22143, g21784, g22937;
wire g26845, g14256, g21956, g18752, g27455, g26395, g30604, g33522, g18374, g29635, g21889;
wire g23103, g27617, g15105, g21980, g10624, g28550, g18643, g7469, g32310, g16204, g28314;
wire g21888, g21824, g26633, g34563, I17542, g27201, g27277, I24675, g33483, g26719, g24289;
wire g18669, g32112, g25927, g32050, g24309, g33862, g18260, g28243, g24288, g27595, g24224;
wire g18668, g27467, g27494, g31949, g18392, g29891, g24308, g21931, g18195, g22015, g18489;
wire g34395, g31948, g32096, g28269, g29575, g15881, g18559, g25491, g18525, g18488, g18424;
wire g28341, g29711, g33904, g24495, g28268, g31252, g29327, g26861, g33252, g13080, g18558;
wire g28655, g30191, g16233, g29537, g34191, g16672, g27822, I27539, g26389, g18893, g25981;
wire g24687, I31011, g27266, g26612, I27538, g26388, g18544, g26324, g32428, g29606, g21024;
wire g18713, g13461, g22084, g31183, g26251, g22110, g24643, g26272, g33847, g21860, g16513;
wire g28694, g29750, g29982, g29381, g18610, g34861, g30247, g18705, g13887, g25990, g23497;
wire g33509, g24669, g31933, g30926, g30045, g18255, g18189, g27588, g15779, g18679, g31508;
wire g34389, g17321, I31112, g34045, g30612, g33508, g24668, g21700, g30099, g33872, g18270;
wire g29796, g17179, g24392, g22685, g18188, g18124, g21987, g18678, g34388, g16026, g28557;
wire g34324, g15081, g13393, g16212, g24195, g28210, g32317, g27119, g30098, g34701, g10721;
wire g20559, g30251, g34534, g23658, g30272, g34098, g19206, g15786, g18460, g18686, g24559;
wire g18383, g29840, g24488, I31096, g24016, g27118, g22417, g11960, g32129, g21943, g25832;
wire g21296, g24558, g18267, g18294, g27616, g26871, g17654, g32128, I17575, g27313, g29192;
wire g30032, g21969, g26360, g25573, g30140, g27276, g27285, g29522, g32323, g24865, g29663;
wire g34140, g22762, g15651, g21968, g10655, g15672, g27305, g25926, g24713, g25045, g18219;
wire g27254, g30061, g33311, g21855, g34061, g14180, g23855, g22216, g18218, g21870, I17606;
wire g28601, g28677, g27036, g29553, g26629, g27177, g27560, g34871, g24189, g31756, g24679;
wire g11244, g29949, g32232, g20188, g18160, g29326, g10838, g28143, g31780, g25462, g24188;
wire g22117, g29536, g22000, g21867, g18455, g24686, g24939, g29757, I31317, g33350, g32261;
wire g18617, g18470, g20093, g33820, g29621, I24576, I24585, g10619, g21714, g23581, g24294;
wire g31152, g25061, I31002, g18201, g33846, I31057, g21707, g21819, g29564, g18277, g14210;
wire g21910, g26147, g30220, g28666, g33731, g28217, g22123, g21818, g17747, g21979, g16896;
wire g27665, g30246, g25871, g20875, g18595, g28478, g18467, g18494, g19500, g24219, g26858;
wire g21978, g11967, g18623, g20218, g30071, g17123, g24218, g21986, g34071, g18782, g27485;
wire g28556, g29509, g32316, g33405, g21741, g26844, g18419, g27454, g26394, g18352, g29634;
wire g29851, g29872, g28223, g15104, g34754, g18155, g21067, g18418, g18822, g30825, g19613;
wire g32056, g18266, g11010, g34859, g18170, I31232, g10677, g22992, g34370, I24674, g21801;
wire g28110, g21735, g21877, g23801, g34858, g30151, g30172, g24915, I31261, g27594, g28531;
wire g17391, g22835, g28178, g18167, g18194, g18589, g22014, g34367, g31787, g34394, g25071;
wire g33113, g33787, g32342, g29574, g31282, g22007, g15850, g29205, g18588, g18524, g28676;
wire g32145, g14791, g32031, g24467, g27519, g33357, g27185, g25147, g32199, g18401, g28654;
wire g33105, g14168, g18477, g26203, g33743, g16802, g18119, g27518, g27154, g34319, g32198;
wire g22116, g16730, g24984, g18118, g21866, g21917, g30227, g31769, g23917, g33640, g26281;
wire g32330, g29592, g30059, g22720, I31316, g30025, g25151, g16765, g15716, g18749, g22041;
wire g26301, g13656, g18616, g18313, g33803, g24822, g26120, g30058, g16690, g11144, g18748;
wire g8643, g25367, I31056, g21706, g18276, g18285, g29350, g26146, g30203, g18704, g34203;
wire g18305, g33881, g30044, g18254, g18809, g21923, g22340, g32161, g22035, g28587, g26290;
wire g18466, g23280, g27215, g27501, g15112, I31271, g30281, g18808, g25420, g24194, g24589;
wire g34281, g29731, g22142, g27439, g34301, g18177, g18560, g30120, g28543, g24588, g32087;
wire g34120, I31342, g32258, g28117, g18642, g25059, g33890, g19788, I31031, g16128, g34146;
wire g34738, g33249, g34562, g28569, g21066, g25058, g16245, g32043, g33482, g32244, g31710;
wire g33248, g10676, I27514, g18733, g27083, g27348, g33710, g22130, g27284, g24864, g22193;
wire g28242, g21876, g21885, g26547, g10654, g11023, g15857, g23885, g27304, g24749, g32069;
wire g12284, g14654, g24313, g22165, g18630, g21854, g15793, g18693, g23854, g31778, g24748;
wire g26226, g32068, g33081, g17193, g21763, g18166, g24285, g25902, g18665, I31132, g31786;
wire g25957, g24704, g25377, g33786, g24305, g16737, g26572, g22006, g28639, g24900, g33647;
wire g32337, g27139, g28293, g33356, g22863, g27653, g28638, g32171, I31161, g18476, g18485;
wire g29787, g26127, g27138, g28265, g34661, g18555, g18454, g25290, g14216, g21916, g30226;
wire g18570, g18712, g33233, g31182, g31672, g27333, g24642, g34226, g14587, g29743, I31087;
wire g34715, g34481, g23314, g32425, g26103, g34572, g10543, g26095, g27963, g23076, g29640;
wire g25366, g29769, g18239, g21721, g33331, g27664, g18567, g18594, g31513, g32010, g33513;
wire g29803, g18238, g26181, g26671, g28586, g24630, g31961, g33897, g17781, g31505, g28442;
wire g33505, g18382, g24009, g33404, g29881, g21773, g18519, g11016, g21942, g13525, g18176;
wire g18185, g22063, g18675, g34385, g33717, g24008, g32086, g30095, g31212, g28116, g18518;
wire g18154, g27312, g24892, g26190, g24485, g24476, I31337, g16611, g27115, g11893, g13830;
wire g22873, g25551, g18637, g25572, I31171, g30181, g30671, g18935, g32322, g24555, g29662;
wire g9217, g21734, g32159, g24712, g29890, g24914, g21839, g21930, g25127, g21993, g32158;
wire g22209, g15856, g15995, g33723, g28237, g21838, g22834, g15880, g31149, g21965, g26088;
wire g26024, g22208, g29710, g28035, g29552, g33433, g23131, g32295, g10841, g29204, g31148;
wire g30190, g13042, g16199, g18215, g25103, g27184, g16736, g18501, g18729, g22021, g27674;
wire g25980, g18577, g33104, g25095, g33811, g33646, g19767, g32336, g34520, g23619, g33343;
wire g21557, g18728, g18439, g30089, g24941, g26126, g30211, g11939, g23618, g25181, g34089;
wire g16843, g18438, g34211, g26250, g13383, g24675, g29647, g30024, g33369, I24048, g17726;
wire g16764, g34088, g13030, g22073, g18349, g14586, g13294, I31086, g29380, g33368, g34860;
wire g16869, g27692, g28130, g28193, g26339, g25931, g18906, g18348, g24637, g19521, g22122;
wire g12692, g12761, g18284, g16868, g34497, g28165, g28523, g18304, g29182, g29651, g33412;
wire I31322, g16161, g15611, g15722, g18622, g22034, g15080, g18566, g30126, g14615, g27214;
wire g34700, g31229, g10720, g21815, g30250, g27329, g32309, g27207, g33896, g31228, g27539;
wire g29331, g32224, g34658, g23187, g26855, g21975, g27328, g25089, g32308, g20215, g29513;
wire g18139, g27538, g18653, g24501, g24729, g25088, g17292, g11160, g17153, I24033, g18138;
wire I26531, g21937, I17552, g34338, g24728, g16244, I31336, g14035, g15650, g34969, g10684;
wire g28703, g18636, g18415, g31310, g18333, g30060, g21791, g28253, g21884, g11915, g34968;
wire g23884, g30197, g31959, g33379, g19462, g25126, g25987, I31017, g13277, g28236, g34870;
wire g34527, g24284, g18664, g27235, g24304, g26819, g27683, g24622, g33742, g26257, g31944;
wire g11037, g18576, g18585, g14193, g18484, g22109, g32260, g28264, g34503, g34867, g25969;
wire g18554, g29620, g33681, g22108, g18609, g27414, g32195, g24139, g25968, g18312, g33802;
wire g33429, g33857, g29646, g30315, g34581, g18608, g27407, g18115, I27534, g33730, g32016;
wire g33428, g34707, g30202, g25870, g30257, g25411, g26094, g31765, g24415, g7763, g24333;
wire g29369, g14222, g21922, g22982, g30111, g18745, g33690, g30070, g34111, g18799, g22091;
wire g23531, g13853, g18813, g30590, g21740, g16599, g26019, g25503, g18798, g28542, g31504;
wire g28453, g27206, g33504, g24664, g29850, g19911, g34741, g16598, g15810, g13524, g17091;
wire g18184, g21953, g18805, g18674, g23373, g30094, g27759, g25581, g25450, g32042, g21800;
wire g24484, g29896, g27114, g32255, g31129, g32189, g21936, g18732, g27435, g18934, g30735;
wire g24554, g27107, g32270, g16125, g16532, g25818, g28530, g31128, g32188, g25979, g28346;
wire g7251, g24312, g18692, g18761, g33245, g24608, g25978, g13313, g15967, g30196, g31323;
wire g29582, g31299, g17192, g34196, g21762, g21964, g25986, g32030, g24921, I31016, g31298;
wire g34526, g18400, g10873, g26077, g24745, g29627, g18214, g28292, g29959, g22862, g28153;
wire g18329, g25067, g25094, g18207, g26689, g29378, g13808, g18539, g11036, g26280, g18328;
wire g27263, g21909, g31232, g25150, g22040, g25801, g26300, g34866, g28136, g18538, g15079;
wire g27332, g29603, g24674, g29742, g21908, g15078, g33697, g30001, g31995, g33856, g26102;
wire g12135, g31261, g26157, g27406, g34077, g27962, g27361, g33880, I31042, g18241, g34706;
wire g21747, g32160, g30256, g25526, g28164, g26231, g33512, g14913, g27500, g29857, g15817;
wire g14614, g24761, g19540, g21814, g18771, g16023, g16224, g11166, g18235, g21751, g21807;
wire g21772, g26854, g15783, g21974, g22062, g18683, g25866, g24400, g27221, g33831, g28327;
wire g29549, g34102, g26511, g34157, g23639, I31267, g10565, g28537, g31499, g33499, g14565;
wire g29548, g23293, g24329, g30066, g22851, g28108, g30231, g15823, g34066, g10034, g25077;
wire g33498, g23265, g24328, g28283, g18515, g23416, g18414, g31989, g14641, g28303, g27106;
wire g21841, g21992, g34876, g18407, g25923, g31988, g33722, g33924, g32419, g15966, g28982;
wire g31271, g12812, g34763, g15631, g27033, g27371, g32418, g26287, g27234, g25102, g21835;
wire g32170, g13567, g22047, g26307, g26085, g29626, g33461, g16669, g33342, g29323, g23007;
wire g31145, g18441, g18584, g24771, g18206, g29533, g12795, g16668, g16842, g17574, g33887;
wire g18759, g22051, g22072, g18725, g32167, g32194, g25876, g33529, I31201, g27507, I31277;
wire g18114, g28192, g18758, g31528, g26341, g18435, g33528, g34287, g19661, g33843, g21720;
wire g33330, g26156, g18107, g27421, g34085, g28663, g32401, g34076, g30596, g26180, g26670;
wire g21746, g33365, g32119, g30243, g31132, g18744, g34054, g31960, g33869, g14537, g18345;
wire g19715, I31037, g29856, g17780, g21465, g18399, g29880, g33868, g26839, g27541, g30269;
wire g22846, g21983, g28553, g25456, g18398, g29512, g32313, I31352, g21806, g26838, g18141;
wire g30268, g18652, g18804, g34341, g25916, g16610, g16705, g17152, g31225, g32276, g27724;
wire g34655, I31266, g27359, g30180, g27325, g30670, g31471, g32305, g32053, g33471, g34180;
wire g33087, g18263, g32254, g27535, g26487, g27434, g27358, g25076, g25085, g18332, g19784;
wire g28252, g12920, g18135, g34335, g25054, g24725, g30930, g32036, g27121, g29316, g19354;
wire g33244, g32177, g18406, g13349, I31167, I18785, g26279, g18361, g24758, g23130, g34667;
wire g34694, g17405, g11083, g34965, g30131, g31069, g19671, g29989, g18500, g22020, g27682;
wire g23165, g28183, g28673, g33810, g27291, g29611, g33657, g26286, g29988, g29924, g34487;
wire g13566, g22046, g26306, g24849, g33879, g24940, g24399, g34502, g30210, g34557, g23006;
wire g23475, g33878, I31022, g18221, g22113, g21863, g26815, g24141, g34279, g11139, g33886;
wire g27134, g30278, g27029, g18613, g31792, g32166, g32009, g25993, g31967, g31994, g22105;
wire I31276, g27028, g29199, g32008, g25965, g29650, g29736, g16160, g29887, g21703, g18273;
wire g24332, g18106, g20135, g18605, g13415, g21347, g13333, g33425, g28213, g15679, g18812;
wire g10948, g18463, g33919, g24406, g29528, I31036, g24962, g29843, g21781, g29330, g16617;
wire g25502, g15678, I31101, I31177, g18951, g30187, g18371, g8721, g28205, g18234, g34187;
wire g17769, g21952, g28311, g23372, g29869, g21821, g17768, I26530, g18795, g30937, g29868;
wire g27649, g34143, g16595, g21790, g24004, g33086, g27648, g24221, g27491, g26486, g18514;
wire g29709, g34169, g21873, g18507, g22027, g23873, g15875, g30168, g29708, g33817, g11115;
wire g33322, g34410, g27981, g25815, g31125, g32176, I31166, g26223, g31977, g33532, g33901;
wire g34479, g34666, g25187, g18163, g15837, g32154, g34363, g25975, g34217, g22710, g30015;
wire g21834, g22003, g34478, g28152, g26084, g28846, g24812, g19855, g33353, g25143, g34486;
wire g18541, g27395, g33680, g18473, g27262, g26179, g12794, I17529, g34556, g18789, g21453;
wire g22081, g29602, g29810, g29774, g34580, g26178, g16194, g27633, g21913, g29375, g30223;
wire g13805, g18788, g18724, g25884, g18359, g34223, g18325, g26186, g23436, g18535, g18434;
wire g18358, g31966, g30084, g27521, g29337, g17786, g30110, g25479, g34084, g15075, g31017;
wire g34110, g25217, g33364, g18121, g22090, g30179, g24507, g18344, g19581, g34179, g27440;
wire g21464, g28020, g28583, g30178, g9479, g24421, g34178, g34740, g16616, g10756, g18682;
wire I31176, g30186, g27247, I31092, g18291, g24012, g17182, g21797, g34186, g34685, g25580;
wire g18173, g27389, g34953, g27045, g31309, I24699, g32083, g32348, g23292, g25223, g16704;
wire g27612, g31224, g32284, g28113, g26423, g27099, g15822, g27388, g27324, g24541, g32304;
wire g30936, g28282, g12099, g27534, g27098, g28302, g25084, g27251, g27272, g25110, g16808;
wire g19384, g18760, g18134, g25922, g34334, g24788, g31495, g24724, g29599, g33495, g22717;
wire g16177, g24325, g25179, g26543, I27503, g18506, g22026, g27462, g33816, g29598, g16642;
wire g25178, g15589, g32139, g27032, g34964, g33687, g31976, g31985, g19735, g27140, g30216;
wire g27997, g28768, g15836, g31752, g34216, g31374, g29322, g33374, g16733, I18671, g29532;
wire g29901, g32333, g15119, g20682, g13771, g25417, g23474, g24682, g22149, g29783, g21711;
wire g26123, g15118, g34909, g24291, g30000, g29656, g34117, g15749, g18649, g22097, g27360;
wire g33842, g18240, g22104, g17149, g33392, g18648, g18491, g31489, g26230, g25964, g33489;
wire g21606, g27162, g34568, g34747, g23606, g29336, g15704, g30242, g18604, g21303, g16485;
wire g18755, g31525, g31488, g31016, g33525, g33488, g28249, g15809, g18770, g22369, g18563;
wire g18981, g21750, g28248, g29966, g28710, g15808, g21982, g27451, g26391, I26948, g23381;
wire g27220, g33830, g29631, g32312, g32200, g33893, g28204, g27628, g34751, g29364, g10827;
wire g25909, g32115, g25543, g12220, g27246, g33865, g21796, g30230, g25908, g18767, g18794;
wire g34230, g18395, g32052, g18262, g22133, g25569, g21840, g25568, g18633, g17133, g34841;
wire g18191, g18719, g22011, g15874, g24649, g29571, g11114, g31270, g16519, g16176, g16185;
wire g25123, g18718, g15693, g18521, g31188, g25814, g27370, g31124, g32184, g28998, g33124;
wire g33678, g24491, g24903, g28233, g16518, g28182, g25772, g28672, g24755, g27151, g34578;
wire g16637, g22310, g18440, g13345, g26275, g30007, I24546, g34586, g18573, g29687, g22112;
wire g18247, g29985, g10890, g21862, g22050, g23553, g18389, g29752, I31312, g29954, g21949;
wire g15712, g18612, g15914, g25992, g18388, g19660, g18324, g24794, g31219, g34116, g24395;
wire g25510, g18701, g26684, g21948, g22096, g32400, g18777, g18534, I14198, g32013, g30041;
wire I31052, g18251, g21702, g31218, g16729, g18272, g21757, g25579, g30275, I24700, g27227;
wire g33837, I24625, g32207, g26517, g34746, g34493, g25578, g15567, g27025, g24191, g24719;
wire g18462, g25014, g32328, g29668, g29842, g27540, g23564, g27058, g30035, g18140, g34340;
wire g27203, g19596, g26130, g29525, g21847, g34684, g10999, g13833, I18819, g26362, g27044;
wire g31470, g23397, g33470, g33915, g32241, g26165, g17793, g10998, g18766, g13048, g23062;
wire g27281, g24861, g24573, g34517, g28148, g14233, g21933, g27301, I14225, g27957, g7804;
wire g25041, g13221, g27120, g17690, g29865, g21851, g21872, g23872, g15883, g18360, g31467;
wire g31494, g28343, I24527, g19655, g33467, g33494, g24324, g27146, g27645, g26863, g18447;
wire g30193, g24777, g27699, g16653, g18162, g25983, g29610, g30165, g22129, g34523, g22002;
wire g22057, g17317, g22128, g33352, I31207, g16636, g18629, g25142, g18451, g26347, g18472;
wire g32414, g29188, g33418, g33822, g18220, g26253, g30006, g31266, g31170, g21452, g18628;
wire g27427, g34475, g17057, g24140, g22299, g29686, g24997, g18246, g21912, g29383, g30222;
wire g34863, g28133, g22298, g26236, g28229, g19487, g29938, g26351, g28228, g25130, g26821;
wire g27661, I31241, g27547, g18591, g31194, g31167, g18776, g18785, g15083, g21756, g18147;
wire g25165, g30253, g16484, g18754, g31524, g33524, g18355, g26264, g33836, g21780, g29875;
wire g32206, g26516, g13507, g27481, g30600, g18825, g18950, g18370, g31477, g33401, g33477;
wire g20162, g30236, g14148, g29837, g14097, g21820, g11163, I24067, g9906, g18151, g31118;
wire g18172, g28627, g32114, g28959, g30175, g32082, g33864, g27127, g21846, g28112, g32107;
wire g15653, g24629, g23396, g18367, g18394, g31313, g24451, g21731, g24220, g20628, g27490;
wire g13541, g30264, g34063, g13473, g30137, g19601, g24628, g32345, g34137, g31285, g34516;
wire g27376, g27385, g33704, g29617, g31305, I24695, I24018, g27103, g33305, g22831, g23691;
wire g26542, g34873, g26021, g18420, g15852, g27095, g18319, g33809, g33900, g33466, g16184;
wire g16805, g21405, g16674, g29201, g32141, g22316, g18318, g18446, g33808, g24785, g18227;
wire g7777, g27181, g30209, g22498, g33101, g19791, g24754, g29595, g29494, g30208, g16732;
wire g21929, g32263, g18540, g10896, g22056, g26274, g29623, g32332, I31206, g21928, g22080;
wire g25063, g24858, g29782, g18203, g26122, g16761, g29984, g34542, g22432, g12931, g29352;
wire g25873, g30614, I24597, I31082, g18281, g27520, g21787, g15115, I31107, g22342, g18301;
wire g30607, g32049, I24689, g26292, g33693, g18377, g19556, g30073, g22145, g18120, g26153;
wire g18739, g21302, g22031, g27546, g30274, g31166, g34073, g10925, g16207, g27211, g32048;
wire g16539, g21743, g21827, g11029, g17753, g18146, g18738, g13029, g15745, g18645, g30122;
wire g24420, g24319, g29853, g16538, g17145, g26635, g11028, g18699, g34565, g15813, g31485;
wire g29589, g33892, g18290, g17199, g24318, g33476, g33485, g21769, g30034, g22843, g24227;
wire g18698, I31141, g25453, g29588, g29524, g29836, g21768, g21803, g28245, g15805, g28626;
wire g30153, g28299, g27700, g22132, g29477, g32273, g32106, g18427, g14681, g19740, g20203;
wire g33907, g18366, I31332, g21881, g27658, g18632, g25905, g17365, g22161, g33074, g34136;
wire g33239, g25530, g27339, g29749, g29616, g7511, g26711, g31238, g32234, g25122, g18403;
wire g18547, g25565, g24301, g28232, g20739, g13491, g22087, g30164, g31941, g33941, g18226;
wire g21890, g13604, g31519, g18715, g27968, g28697, g31185, g18481, g33519, g29809, g33675;
wire g24645, g28261, g26606, g28880, g18551, g22043, g26303, g31518, g31154, g18572, g33518;
wire g29808, g21710, I31221, g24290, g29036, g27411, g34474, g24698, g21779, g26750, g12527;
wire g23779, g18127, g22069, g25408, g30109, g26381, g34109, g29642, g33883, g21778, g22068;
wire g26091, g18490, g30108, g32163, g32012, g34108, g24427, g21786, g27503, I24054, g30283;
wire I31106, g18784, g18376, g18385, g29733, g18297, g17810, g18103, g10626, g34492, g13633;
wire g25164, g21945, g28499, g18354, g29874, g27714, g21826, g21999, g26390, g31501, g18824;
wire g27315, g33501, g29630, g24403, g29693, g30982, g34750, g16759, g18181, g21998, g18671;
wire g34381, g23998, g33728, g27202, g19568, g30091, g32325, g29665, g16758, g34091, g24226;
wire g13832, g28722, g28924, g30174, g29008, g12979, g24551, g24572, g33349, g25108, g21932;
wire g32121, g18426, g33906, g13247, g29555, g21513, g18190, g22010, g23513, g34390, g10856;
wire g11045, g15882, g27384, g29570, g29712, I24694, g33304, g14261, g18520, g21961, g22079;
wire g27094, g30192, g31566, g13324, g29907, g32291, g16804, g21404, g28199, g22078, g23404;
wire g32173, g18546, g25982, I31012, g18211, g21717, g28198, g24297, g22086, g25091, g20095;
wire I24619, g29567, g29594, g12735, g31139, g28528, g28330, g26252, g11032, g34483, g18497;
wire g32029, g24671, g14831, g22125, g29382, g27526, g34862, g29519, g32028, g19578, g33415;
wire g22158, g14316, g33333, g18700, g17817, g18126, g18659, g18625, g18987, g29518, g18250;
wire g24931, g15114, g25192, g26847, g34948, g18658, g27457, g26397, g15082, g23387, g31963;
wire g29637, g22680, g34702, g15107, g23148, g34757, g17783, g25522, I31121, g24190, g18339;
wire g18943, g29883, g18296, g21811, g28225, g23104, g23811, g23646, g18644, g28471, g16221;
wire g18338, g30564, g9967, g28258, g21971, g34564, g15849, g31484, g24546, g33484, g16613;
wire I31291, g15848, g19275, g31554, g30673, g27256, g19746, g28244, g34183, g18197, g22017;
wire g15652, g15804, g34397, g25949, g27280, g31312, g29577, g30062, g27300, g10736, g10887;
wire g31115, g18411, g25536, g25040, g26213, g34509, g21850, g28602, g23412, g28657, g25904;
wire g33921, g19684, g34508, g10528, g34872, I18740, g24700, g28970, g24659, g14528, g26205;
wire g23229, g16234, g29349, g22309, g20658, g18503, g22023, g26311, g24658, I24015, g10869;
wire g22308, g28171, g33798, g21716, g30213, g24296, g18581, g18714, g26051, g18450, g31184;
wire g34213, g18315, g33805, g33674, g24644, g29622, g29566, g18707, g18819, g18910, g18202;
wire g30047, g18257, g26780, g30205, g32191, g18818, g18496, g34205, g31934, g18111, g21959;
wire g21925, g26350, g25872, g28919, g14708, I18762, g28458, g24197, g24855, g27660, g16163;
wire g22752, g15613, g18590, g21958, g21378, g23050, g28010, g23958, g24411, g30051, g26846;
wire g18741, g34072, g23386, g30592, g18384, g29636, g21742, g17752, g27480, g34756, g23742;
wire g28599, g21944, g33400, g29852, g17643, g15812, g13319, g27314, g24503, g27287, g32045;
wire I24685, g33329, g31207, g18150, g10657, g18801, g18735, g25574, g27085, g32324, g29664;
wire g33328, g21802, g22489, g21857, g23802, g16535, g20581, g10970, g23857, g13059, g13025;
wire g30152, g24581, g24714, g32098, g24450, g21730, g24315, g21793, g32272, g22525, g28159;
wire I31262, g10878, g18196, g22016, g28125, g15795, g18695, g28532, g34396, I18568, g24707;
wire g30731, g29576, g29585, g21765, g28158, I27523, g18526, g27269, g29554, g23690, g19372;
wire g26020, g33241, g34413, g17424, g11044, I31191, g27341, g10967, g29609, g27268, g32032;
wire g25780, g15507, g32140, g28144, g18402, g18457, g24590, g29608, g27180, g19516, g20094;
wire g27335, g33683, g13738, g25152, g22042, g26302, g26357, g29799, g30583, g16760, g27667;
wire I31247, g18706, g18597, g27965, g13290, g29798, g22124, g27131, g30046, g18256, g29973;
wire g18689, g31991, g33515, g33882, g18280, g29805, g33414, g22686, g22939, g18688, g18624;
wire g32162, g18300, g24196, g33407, g34113, g27502, I31251, g11427, g22030, I31272, g22938;
wire g27557, g22093, g23533, g11366, g27210, g21298, g29732, g28289, g21775, I16671, g13632;
wire g18157, g23775, g22065, g34105, g28224, g34743, I17585, g28571, g24402, g29761, I31032;
wire g18231, g21737, g32246, g27469, g22219, g25928, g8583, g27286, g33441, g31206, g10656;
wire g27039, g22218, g28495, g32071, I31061, g21856, g10823, g14295, g21995, g31759, g23856;
wire g14680, g33759, g33725, g24001, g21880, g29329, g25113, g18511, g29207, g25787, g32147;
wire g18763, g31758, g33114, g24706, g26249, g33758, g22160, g27601, g33082, g21512, g29328;
wire g27677, g25357, g29538, g11127, g24923, g25105, g10966, g31744, g24688, g26204, g24624;
wire g24300, I24579, g26779, g33345, g32151, g32172, I31162, g31940, g18456, g33849, g30027;
wire g33399, g21831, g26778, g34662, g16845, g11956, g18480, g32367, g34890, g28668, g34249;
wire g13095, g30482, g24231, g13888, g26945, g30552, g34003, g23989, g29235, g28525, g34204;
wire I28566, g14309, I30330, g24854, g30081, g32227, g33962, g19575, g27556, g25662, g28544;
wire g30356, g27580, g34647, g26932, I31859, g33049, g30380, g34826, g16926, I25736, I31858;
wire g33048, g7684, g25710, g28610, g26897, g34090, g26961, g28705, g28042, g30672, g34233;
wire g13211, g33004, g31221, g23198, I31844, g27179, g28188, g33613, g34331, g30513, g30449;
wire g33947, g34449, g25647, g24243, g33273, g28030, g33605, g25945, g28093, g30448, g34897;
wire g34448, g30505, g29114, g30404, g28065, g27800, g24269, g34404, g33951, g33972, g24341;
wire g33033, g24268, g25651, g25672, g33234, g34026, g32427, g13296, g23087, g29849, g13969;
wire g26343, g19522, g29848, g24335, g26971, g34723, g30433, g34149, g30387, g24965, g32226;
wire g29263, g34620, g34148, g25717, g27543, g30104, g33012, g19949, g30343, g34646, g24557;
wire g24210, g27569, g34971, g33541, g31473, g28075, g30369, g24443, g19904, g23171, g24279;
wire g26896, g34369, g28595, g14030, g30368, g24278, g25723, g28623, g34368, g33788, g31325;
wire g32385, g31920, g32980, g30412, g33535, g24468, g32354, g34850, g34412, g28419, g27974;
wire g33946, g25646, g28418, g20187, g26959, g26925, g34011, g26958, g29273, g31291, g17570;
wire g33291, g26386, g32426, g28194, g28589, g26944, g20169, g27579, g29234, g30379, g34627;
wire g27578, g17594, g28401, g31760, g34379, g33029, g32211, g30378, g21901, g20217, g33028;
wire g30386, g24363, g26793, g28118, g13526, g24478, g34603, g25716, g28749, g26690, g25582;
wire g28748, g28704, g24580, g31927, g30429, g28305, g28053, g32987, g32250, g34802, g25627;
wire g30428, g34730, g34793, I26643, g13077, I18492, g28101, g33240, g13597, g28560, g31903;
wire g30549, g25603, g25742, g31755, g33604, g30548, g10589, g29325, g13300, g31770, g30504;
wire g28064, g33563, g33981, g25681, g28733, g26299, g30317, g25730, g22304, g14119, g31767;
wire g33794, g34002, g33262, g31899, g34057, g28665, g30128, g33990, g24334, g25690, g26737;
wire g29291, g31898, g34626, g30533, g22653, g30298, g23687, g26880, g24216, g23374, g32202;
wire g22636, g26512, g32257, g13660, g32979, g29506, g34232, g32978, g28074, g33573, g31247;
wire g28594, g31926, g32986, g27253, g33389, g33045, g22664, g34856, g25626, g33612, g34261;
wire g34880, g8921, g30512, g33534, g27236, g32094, g31251, g22585, g33251, g24242, g33272;
wire g28092, I30124, g28518, g21893, g29240, g26080, I12583, g25737, g26924, g30445, g33032;
wire g34445, g30499, g33997, g25697, g25856, g30498, g25261, g33061, g24265, g26342, g31766;
wire g31871, g30611, g24841, g34611, g23255, g34722, g26887, g28729, g28577, g24510, g30432;
wire g28728, g29262, g27542, g27453, g23383, g24578, g30461, g30342, g34461, g26365, I18452;
wire g26960, g34031, g31472, g28083, g28348, g34199, g32280, g9984, g34887, g31911, g30529;
wire g33628, g27274, g31246, g25611, g19356, g25722, g28622, g28566, g30528, g9483, g30393;
wire g27122, g34843, g34330, g30365, g24275, g29247, g31591, g31785, g33591, g24430, g24746;
wire g32231, g25753, g31754, g28138, g24237, g33950, g29777, g24340, g25650, g25736, g29251;
wire g29272, g28636, g19449, g28852, g34259, g30471, g33996, g34708, g26657, g25696, g26955;
wire g34258, g24517, g26879, g26970, g25764, g28664, g26878, g16867, g25960, g34043, g26886;
wire g25868, g28576, g31319, g27575, g26967, g33318, g34602, g25709, g30375, g34657, g28609;
wire g33227, g9536, g33059, g33025, g25708, g34970, I29986, g23822, g33540, g27108, g33058;
wire g30337, g32243, g26919, g28052, g27283, g26918, g28745, g15968, I31854, g33044, g34792;
wire g32268, g23194, g33281, g31902, g30459, g30425, g33957, g24347, g34459, g25602, g12982;
wire g25657, g24253, g25774, g29246, g30458, g34458, g33562, g34010, g24236, g25878, g28732;
wire g33699, g32993, g30545, g30444, g29776, g24952, g24351, g33290, g26901, g34444, g24821;
wire g29754, g34599, g32131, g20063, g34598, g15910, g24264, g23276, g27663, g28400, g32210;
wire g21900, g16866, g28329, g30532, g32279, g34125, g22652, g13762, g34977, g25010, g31895;
wire g28328, g33547, g34158, g24209, g34783, g28538, g26966, g25545, g30561, g7673, g30353;
wire g24208, g25599, g34353, g29319, g25598, g33551, g33572, g30336, g29227, g13543, I31839;
wire I31838, g28100, g20905, g34631, g30364, g34017, g24274, g13242, g33956, g24346, g33297;
wire g25656, g31889, g33980, g24565, g21892, g25680, g16876, g29281, g31888, g20034, g29301;
wire g27509, g34289, g24641, g34023, g34288, g32217, g26954, I18449, g31931, g29290, g25631;
wire g30495, g32223, g29366, g27574, g34976, g26392, g27205, g33546, g30374, g16076, g34374;
wire I30728, g33024, g34643, g28435, g28082, g26893, g29226, g28744, g34260, g28345, g29481;
wire g30392, g30489, g33625, g32373, g33987, g31250, g25687, g30559, g30525, g30488, g30424;
wire g25752, g34016, g30558, g27152, g33296, g25643, g29490, g16839, g28332, g30544, g33969;
wire g25669, g28135, g29297, g33060, g33968, g26939, g25668, g33197, g28361, g32216, g27405;
wire g26938, g31870, I28147, g24840, g34610, g24390, g30189, g28049, g34255, g34189, g30270;
wire g28048, g20522, g26875, g32117, I23163, g31894, g31867, g30460, g30383, g34460, g30093;
wire g34030, g25713, g28613, g33581, g33714, g29520, g34267, g34294, g31315, g33315, g31910;
wire g13006, g25610, g31257, g25705, g28605, g33257, g32123, g33979, g33055, g16187, g25679;
wire g33070, g33978, g25678, g26915, g33590, g15965, g28371, I30745, g32230, g33986, g24252;
wire g25686, g33384, g33067, g12768, g29250, g32992, g32391, g30455, g34455, g11372, g31877;
wire g30470, g34617, g22648, I12611, g29296, g33019, g30201, g33018, I30761, g30467, g30494;
wire g34467, g34494, g29197, g34623, g34037, I30400, g27248, g30984, g27552, g31917, g30419;
wire g31866, g30352, g27779, g25617, g24213, g23184, g28724, g34352, g28359, g30418, g32275;
wire g31001, g28358, g34266, g33001, g34170, g24205, g33706, g33597, g32237, g31256, g33256;
wire g25595, g31923, g32983, g19879, g28344, g22832, g33280, g25623, g20051, g25037, g33624;
wire g34167, g34194, g26616, g19337, g28682, g29257, I23755, g30524, g27233, g16800, g29496;
wire g27182, g30401, g30477, g26305, g24350, g26809, g33066, g26900, g33231, g29741, g32130;
wire g34022, g28134, g31876, g31885, g32362, g34616, g25589, g29801, g29735, g25588, g34305;
wire g25836, g27026, g34254, g30466, g34809, g34900, g26733, g34466, g34808, g32222, g23771;
wire g26874, g34036, g30560, g34101, g31916, g34642, g25749, g25616, g28649, g33550, g32347;
wire g33314, g31287, g15800, g32253, g25748, g33287, g34064, g30733, g31307, g33076, g34733;
wire g26892, g25704, g22447, g33596, g33054, g32236, g8790, g32351, g32372, g34630, g34693;
wire g24282, g26914, g29706, g8461, g31269, g34166, g34009, g19336, g26907, g29256, g31773;
wire I30399, g31268, g32264, g34008, g29280, g33268, g30476, g30485, g29300, g31670, g8904;
wire I31863, g30555, g30454, g34454, g25733, g13091, g22591, g27133, g28719, g28191, g31930;
wire g32209, g33993, g25630, g28718, g25693, g29231, g33694, g32208, g33965, I12783, g25665;
wire g34239, g34238, g23345, g26883, I23162, g33619, g33557, g29763, g30382, g30519, g33618;
wire g28389, g30176, g28045, g30092, g31279, g24249, g33279, g25712, g28099, g30518, I22280;
wire g28388, g16430, g28701, g24248, g33278, g12925, g28777, g28534, g28098, g32346, g34637;
wire g24204, g33286, g31468, g31306, I31873, g33039, g29480, g27742, g22318, g25594, g33038;
wire g29287, g29307, g28140, g26349, g33601, g25941, g33187, g33975, g27429, g26906, g25675;
wire g29243, g26348, g30501, g28061, g34729, g32408, g30439, g34728, g34439, g29269, g25637;
wire g24233, g25935, g30438, g19525, g19488, g34438, g29268, I25613, g31884, g33791, g30349;
wire g34349, g8417, g30348, g22645, g34906, g29734, g30304, g33015, g34622, g25729, g26636;
wire g28629, g25577, g28220, g25728, g28628, g33556, g24212, g26963, g33580, g29487, g23795;
wire g28071, g29502, g27533, I29351, g28591, g25906, g28776, g30415, g30333, g34636, g22547;
wire g29279, g31922, g32982, g33321, g25622, g29278, g19267, g22226, g24433, g20148, g29286;
wire g27232, g7404, g29306, g28172, g33685, g7764, g33953, g24343, g26921, g25653, g32390;
wire g27261, g30484, g30554, g22490, g13820, g26813, g15727, g25636, g30609, g34609, g28420;
wire g30608, g28319, g30115, g29143, g34608, g17490, g26805, g31762, g23358, I30760, g31964;
wire g33964, g25664, g28059, g29791, g16021, g26934, g28058, g29168, g33587, g24896, g34799;
wire g25585, g25576, g29479, g34798, g31909, g28044, g33543, g19595, g29478, g19467, g25609;
wire g34805, g31908, g33000, g29486, g32252, g25608, g33569, g30732, g27271, I18495, g34732;
wire g26329, g33568, g25745, g29223, g26328, g28562, g14844, g34761, g28699, g27031, g33123;
wire I30755, g28698, g31751, g31772, g30400, g33974, g30214, g34013, g25805, g25674, g31293;
wire g33293, g30539, g34207, g22659, g22625, g25732, g34005, g28632, g33265, g30538, g29373;
wire I30262, g33992, g25761, g28661, g28403, g22644, I12782, g33579, g14044, g28715, I30718;
wire g33578, g31014, g27225, g33014, g23770, g26882, g28551, g31007, g27258, g34100, g33586;
wire g33007, g25539, g13662, g34235, g27244, g28490, g33116, g33615, g23262, g21899, g30515;
wire g30414, g28385, g33041, g28297, g21898, g34882, g28103, g24245, g33275, g28095, g30407;
wire g34407, g27970, g31465, g26759, g26725, g28671, g33983, g22707, g33035, g27886, g25683;
wire g29242, g26082, g11380, g30441, g34441, g24232, g34206, g26940, I25612, g34725, g24261;
wire g29230, g27458, g29293, g30114, g30435, g29265, g28546, g28089, g23251, g28211, g34107;
wire g19555, g28088, g30345, g30399, g34849, g34399, g25584, g28497, g33006, g30398, g26962;
wire g26361, g23997, g30141, g34804, g28700, g25759, g28659, g25725, g28625, g14888, g32357;
wire g27159, g27532, g25758, g34263, g34332, g33703, g28296, g31253, g27561, g33253, g25744;
wire g28644, g30406, g24432, g30361, g34406, g24271, g33600, g25940, g31781, g23162, g33236;
wire g30500, g29275, g28060, g33952, g24342, g25652, g26947, g8905, g29237, g28527, g33063;
wire g34004, g26951, g26972, g31873, g19501, g34613, g32249, g30605, g27289, g34273, g34605;
wire g18879, g28581, g27224, g30463, g27571, g28707, g34463, g23825, g30371, g28818, g34033;
wire g34234, g28055, g33542, g33021, g24259, g28070, g31913, g18994, g24471, g34795, g25613;
wire g24258, g33614, g17511, g32999, g33607, g31905, g31320, g30514, g32380, g31274, g25605;
wire g29222, g24244, g33274, g30507, g32998, g28094, g28067, g33593, g26789, g32233, g12954;
wire g23319, g30421, g33565, g34421, g26359, g28735, g23318, g30163, g33034, g26920, g34012;
wire g29253, g24879, g33292, g26946, g30541, g30473, g24337, g27489, g29236, g28526, g26344;
wire g27016, g30359, g34724, g28402, g30535, g30434, g19576, g30358, g34535, g29264, g29790;
wire g16928, g27544, g33164, g17268, g24919, g30344, g31891, g28077, g33891, g31474, g33575;
wire g24444, g30291, g25789, g32387, g25724, g28688, g33537, g22487, g28102, g33283, g27383;
wire g33606, g31303, g33303, g34029, g26927, g30506, g28066, g21895, g34028, g32368, g33982;
wire g25682, g29274, g24561, g24353, g26903, g35000, g11737, g9012, g26755, g28511, g32229;
wire g26770, g24336, g27837, g33390, g32228, g25760, g29292, g34649, g34240, g30491, g34903;
wire g23297, g34604, g26899, g30563, g26898, g28085, g28076, g28721, g28596, g28054, g33553;
wire g15803, g22217, g33949, g31326, g32386, g30395, g34794, g25649, I26644, g27037, g34262;
wire g33536, g33040, g33948, g25648, g28773, g31757, g31904, g34633, g25604, g25755, g33621;
wire g34719, g28180, g28670, g26926, g32429, g30521, g14511, g33564, g26099, g29283, g28734;
wire g28335, g29303, g24374, g30440, g34440, g25767, g28667, g33062, g22531, g27589, g16448;
wire g30389, g24260, g27524, g25633, g31872, g24842, g30388, g34612, g25719, g28619, g34099;
wire g30534, g19441, g25718, g28618, g34251, g28279, g26766, g30462, g23296, g34462, g28286;
wire g32245, g34032, g28306, g33574, g33047, I26741, g31912, g31311, g23197, g25612, g28815;
wire g29483, g16811, g25701, I30055, g24705, g33051, g24255, g33592, g30360, g24270, g26911;
wire I30741, g30447, g21894, g34447, g32995, g24460, g29904, g13657, g29252, g28884, g26785;
wire g24267, g30451, g30472, I30735, g34629, g17569, g34451, g34628, g34911, g26950, g22751;
wire g27008, g22639, g27555, g28580, g29508, g8476, g20160, g30355, g27570, g31929, g32989;
wire g30370, g25629, g27907, g16959, g31020, g31928, g14187, g32988, g28084, g33020, g33583;
wire g25628, g25911, g27239, g19605, g33046, g32271, g34172, g28179, g27567, g27238, g17510;
wire g30394, g30367, g24201, g24277, g25591, g33282, g28186, g28685, g31302, g28373, g25754;
wire g30420, g28417, g24782, g30446, g34446, g34318, g28334, g29756, g24352, g26902, g26957;
wire g34025, g31768, g26377, g30540, g13295, g15582, g24266, g32132, g9535, g31881, g28216;
wire g24853, g22684, g32259, g30377, g32225, g34957, g34377, g33027, I22912, g31890, g24401;
wire g30562, g31249, g19359, g34645, g19535, g31248, g28747, g34290, g33552, g13289, g33003;
wire g33204, g26895, g31779, I31843, g10800, g19344, g27566, g28814, g30427, g20276, g29583;
wire g32375, g14936, g30366, I30054, g24276, g28751, g28772, g34366, I31869, g34632, g25739;
wire g24254, I31868, g28230, g33945, g25738, g25645, g30547, g30403, g33999, g33380, g25699;
wire g34403, g29282, g28416, g16261, g32994, g33998, g29302, g25698, g29105, g30481, g7932;
wire g26956, g30551, I30734, g26889, g31932, g26888, g23721, g25632, g28578, g30127, g29768;
wire g34127, g31897, g30490, g33961, g25661, g27484, g30376, g30385, g26931, g30103, g34376;
wire g34297, g34103, g33026, g30354, g22516, g34980, g33212, g25715, g8679, g34095, g30824;
wire g28720, g28041, g17264, g28430, g32125, g28746, g32977, g19604, I30469, g29249, g26089;
wire g24907, I30468, g29482, g34931, g29248, g33149, g30426, g32353, g33387, g24239, g9055;
wire g28684, g32144, g33620, g34190, g24238, g30520, g28517, g30546, g33971, g29786, g25671;
wire g34024, g13938, g24518, g22530, g28362, g30497, g24935, I12903, g29233, g26969, I18421;
wire g32289, g22641, g34625, g26968, g17464, g31896, g34250, g32288, g28727, g16258, g33011;
wire g30339, g24215, g24577, g30338, g34644, g33582, g19534, g27241, g28347, g29717, g33310;
wire g26894, g33627, g31925, g32976, g32985, g24349, g16810, g25700, g28600, g25659, g25625;
wire g20083, g30527, g30411, g33050, g32374, g33958, g24348, g34411, g16970, g25658, g28372;
wire g23217, g33386, g26910, g33603, g25943, I30740, g13623, g25644, g30503, g28063, g34894;
wire g29148, g32392, g27515, g30450, g24653, g34450, g13155, g31793, g34819, g34257, g28209;
wire g30496, g8956, g34979, g34055, g33549, g28208, g26877, g34978, g33548, g27584, g25867;
wire g25894, g30384, g31317, g33317, g29229, g25714, g28614, g25707, g25819, g28607, g29228;
wire g25910, g28320, g31002, g28073, g33002, g33057, g34801, g34735, g32124, g29716, g24200;
wire g31245, g34019, g26917, g15792, g26866, g28565, g33626, g33323, g34695, g25590, g34018;
wire g30526, g32267, g32294, g33298, g25741, g28641, g31775, I30123, g8957, g24799, g30402;
wire g24813, I30751, g30457, g34402, g34457, g26923, g32219, g33232, g25735, g25877, g28635;
wire g32218, g27135, g33995, g34001, g33261, g25695, g31880, g30597, g34256, g29802, g34280;
wire g29730, g30300, g29793, g34624, g34300, g15125, g26876, g26885, g23751, g25917, g32277;
wire g24214, g31316, g33316, g22634, g24207, g22872, I29985, I22958, g34231, g29504, g25706;
wire g25597, g32037, g33989, g33056, g13570, g25689, g13914, g33611, g31924, g32984, g33988;
wire g25688, g28750, g25624, g26916, g30511, g20241, g32352, I30746, g24241, g33271, g27972;
wire g32155, g15017, g28091, g32266, g29245, g26721, g29299, g33031, g30456, g34456, g29298;
wire g24235, g13941, g31887, g28390, g30480, g30916, g29775, I26523, g25885, g30550, g30314;
wire g23615, g30287, g34314, g30307, g33393, g23720, I12902, g25763, g29232, g31764, g23275;
wire g34721, g31869, I30193, g30431, g33960, g25660, g29261, g31868, g26335, g19572, g22152;
wire g26930, g34269, g30341, g26694, g26965, g33709, g34268, g31259, g32285, g33259, g28536;
wire I30727, g31258, g24206, g13728, g28702, g30734, I22298, g30335, g34734, g25721, g28621;
wire g25596, I31853, g33043, g31244, g20082, g28564, g23193, I23756, g26278, g33069, g33602;
wire g25942, g31774, g7834, g30487, g31375, g33068, g33955, g24345, g25655, g31879, g30502;
wire g28062, g30557, g33970, g34619, I22880, g25670, g29271, g31878, I31864, g30443, g34618;
wire g24398, g30279, g34443, g25734, g28634, g28851, g31886, g29753, g25839, g34278, g30469;
wire g33967, g33994, g27506, g30286, g25694, g25667, g24263, g34286, g30468, g34468, g34039;
wire g34306, g29529, g22640, g34038, g31919, g32454, g25619, g15124, g26884, g28574, g31918;
wire g28047, g33010, g34601, g29764, g25618, g34975, g24500, g33545, g9013, g26363, g33599;
wire g32239, g28051, g27240, g28072, g33598, g32238, I29352, g28592, I31874, g34791, g22662;
wire g34884, g29259, g29225, g30410, g31322, g14062, g34168, g27563, g29258, g31901, g33159;
wire g30479, g33977, g30363, g25601, g12981, g24273, g25677, g31783, g23209, g30478, g34015;
wire g29244, g33561, g30486, g31295, g26922, g28731, g33295, g31144, g25937, g30556, g24234;
wire g13973, g29068, g25791, g28691, g29879, g26953, g28405, g33966, g25666, g33017, g26800;
wire g34321, g30531, g23346, g29792, g12832, g13761, g16022, g26334, g28046, g32349, g31289;
wire g30373, g33289, g22331, g26964, g34373, g33023, g31288, g23153, g33288, g31308, g33571;
wire g30417, g34800, g34417, g28357, g30334, g28105, g28743, g29078, g26909, I18385, g34762;
wire g25740, g26908, g28640, g30423, g33976, g33985, g24946, g25676, g25685, I30750, g33954;
wire g21891, g24344, g25654, g25936, g30543, I26522, g31260, g34000, g26751, g33260, g29295;
wire g31668, g14583, g25762, g28662, g26293, g33559, I30192, g33016, g25587, g33558, g23750;
wire g31893, g34807, g34974, g31865, g33544, g34639, g12911, g30293, g23796, g28778, g16239;
wire g34293, g34638, g34265, g30416, g27591, g34416, g29289, g25747, g28647, g33610, g29309;
wire g30391, g33042, g27147, g31255, g29288, g33255, g29224, g30510, g29308, g24240, g33270;
wire g28090, g30579, g27858, g25751, g28651, g29495, g33383, g25639, g34014, g33030, g31267;
wire g25638, g34007, g16883, g33267, g33294, g27394, g28331, g30442, g33065, g34442, g28513;
wire g31875, g29643, g34615, g33219, g24262, g28404, g34720, g34041, g28717, g30430, g30493;
wire g28212, g29260, g25835, g30465, g34465, g25586, g34237, g30340, g29489, g34035, g29488;
wire g34806, g23183, g28723, g33617, g31915, g25615, g30517, g28387, g31277, g25720, g24247;
wire g33277, g14182, g15935, g28097, g28104, g25746, g28646, g33595, g32235, g27562, g33623;
wire I30756, g33037, g30362, g34193, g24251, g24272, g31782, g27290, g28369, g30523, g33984;
wire g25684, g29255, g28368, g26703, g29270, g32991, g30475, g34006, g28850, g33266, g23574;
wire g13972, g34727, g26781, g30437, g26952, g29294, g29267, g19619, g8863, g19557, I22830;
wire g27403, g33589, g30347, g28716, g34347, g33588, g34253, g27226, g28582, g34600, g24447;
wire g14387, g34781, g27551, g27572, g33119, g28310, g34236, g30351, g30372, g25727, g33118;
wire g34372, g31864, g33022, g26422, g31749, g16052, g7450, g28050, g33616, g33313, g30516;
wire g34264, g28386, g34790, g31276, g25703, g28603, g24246, g33276, g28096, g32399, g33053;
wire g31254, g27980, g33254, g31900, g31466, g32398, I22267, g25600, g26913, g28681, g23405;
wire g29277, g30422, g33036, g28429, g33560, g24355, g28730, g26905, g25821, g28428, g30542;
wire g30453, g33064, g19363, g28690, g34021, g34453, g27426, g28549, g24151, g33733, g32361;
wire g34726, g28548, g31874, g30436, g19486, g34614, g29266, g34607, g30530, g28317, g33009;
wire g34274, g30346, g25834, g27024, I31849, g33008, g30464, g32221, g34464, g31892, I31848;
wire g28057, g34034, g33555, g34641, g34797, g25726, g33570, g31914, g34292, g28323, g33914;
wire g34153, g27126, g25614, g28533, g31907, g30409, g27250, g26891, g24203, g25607, g10802;
wire g15732, g28775, g30408, g29864, g34635, g25593, g33567, g33594, g32371, g29313, g24281;
wire g33238, g26327, g22225, g29748, g22708, g29276, g29285, g29305, g29254, g33176, g16882;
wire g30474, g25635, g31883, g30537, g19587, I30331, g34537, g13794, g34283, g30492, g34606;
wire g34303, g28316, g27581, g27450, I30717, g33577, g30381, g25575, g28056, g32359, g27257;
wire g29166, g25711, g28611, g24715, g32358, g34796, g29892, g27590, g29476, g29485, g31906;
wire g30390, g32344, g31284, g25606, g28342, g31304, g29914, g21897, g33622, g33566, g25750;
wire g26949, g28650, g30522, g27150, g34663, g29239, g26948, g24354, g27019, g26904, g29238;
wire g30483, g30553, g22901, g28132, g13997, g29176, g30536, g26673, g34040, g33963, g25663;
wire g34252, g34621, g28708, g26933, g28087, g33576, g33585, g24211, g28043, g33554, g32240;
wire g30397, I26742, g33609, g29501, g33312, g30509, g33608, g28069, g33115, g25702, g25757;
wire g28774, g30508, g31921, g28068, g32981, g28375, g33052, g34634, g25621, g31745, g21896;
wire g24250, g26912, g27231, g29284, g32395, g24339, g33973, g29304, g32262, g23716, g25673;
wire g32990, I18417, g24338, g11370, g30452, g34452, g13858, g33732, g30311, g24968, g25634;
wire g31761, g33692, g19475, g27456, g26396, g28545, g28078, g33013, g22669, g32247, I18543;
wire g28086, g32389, g30350, g34350, g33539, g32388, g33005, g27596, g11025, g28817, g33538;
wire g28322, g27243, g30396, g32251, g13540, g27431, g20202, g34731, g29484, g24202, g26929;
wire g24257, g30413, g24496, g31241, g26928, g17488, g25592, g25756, g28561, g28295, g28680;
wire g32997, g30405, g16173, g34405, g33235, g23317, I22852, g29813, g22679, g23129, g13699;
wire g34020, g25731, g28631, I28567, I24117, g32360, g16506, g15789, I30261, g34046, g31882;
wire g33991, g14078, g20196, g25691, g27487, g34282, g23298, g30357, g28309, g32220, g26881;
wire g16927, g25929, g28308, g27278, g29692, g24457, g14977, g25583, g33584, g34640, g19274;
wire g19593, g34803, g28816, g20077, g23261, g26890, g28687, g29539, g32355, g34881, g24256;
wire g32370, g28374, g24280, g25743, g28643, g27937, g32996, g34027, g29241, g13385, g11980;
wire g13889, g13980, g12169, I22761, I13443, I14185, g16719, I14518, g10224, g17595, g22984;
wire I12346, g12478, g21432, g28830, I14883, g19474, g11426, g11190, g9852, g23342, g27223;
wire I15089, g22853, g25003, I15088, g24916, g25779, g12084, g28270, g22836, g21330, g20076;
wire g21365, g23132, I22683, g28938, g9825, g7201, g15719, g27654, g22864, I20165, g14489;
wire g29082, g25233, g24942, I26459, g15832, g14830, I32431, g9972, I20222, g17748, g11969;
wire g20734, g28837, I25244, g11968, g13968, g15045, g12423, g27587, g20838, g13855, g19483;
wire g10610, g11411, I13110, g22642, g12587, g13870, g13527, g23810, g20619, g16628, I23119;
wire g10124, g12000, I23118, g22874, g10939, g13867, g14686, I12840, g29049, g16776, g13315;
wire g11707, I18530, g20039, I14609, I13334, g13257, g29004, g21459, g11979, g13496, g11590;
wire g12639, g22712, g23010, g7897, g24601, g13986, g12293, g24677, g12638, g24975, g10160;
wire g17712, g12416, g14160, g28853, g13067, g28167, I18635, g10617, g16319, I32187, I12252;
wire g14915, g22941, I17406, g12578, g27586, g12014, g14075, g15591, g28864, g10623, g17675;
wire g23656, g21353, I13751, g14782, I14400, g12116, g14984, g13866, I18537, g16281, g28900;
wire g14822, g14170, g15844, I22972, g21364, I13391, g13256, I13510, g11923, g12340, g12035;
wire g13923, I15300, g9830, g20186, g20676, g21289, I12205, g13102, g25429, g23309, g28874;
wire g29121, g21288, g7582, I13442, g13066, g24936, g31262, g10022, g14864, g8769, g7227;
wire I32186, g12523, g28892, g13854, g11511, I14991, g8967, g13511, g20216, g14254, g28914;
wire g29134, g28907, g12222, g29028, g22852, g14101, g25002, I29297, g14177, g11480, I26460;
wire I22946, I18536, I15287, I14206, g16956, I26093, I15307, g23195, g13307, I15243, g16181;
wire g12351, g24814, g22312, g28935, g24807, I15341, g14665, g24974, g31997, g14008, I14399;
wire I22760, g9258, g22921, g15715, g17312, g25995, g14892, g17608, I14398, g15572, I18634;
wire I15335, g34056, g14570, g11993, g13993, I23963, g9975, g21124, I14332, g13667, g13131;
wire g10567, g20007, I23585, g28349, g29719, g21294, g25498, g28906, g13210, g34650, g16625;
wire g17732, g10185, g11443, g12436, g11279, g14519, I29296, g14675, I25219, g27593, I26419;
wire I22755, g12073, g14154, g17761, I26418, g13469, g25432, g10935, g14637, I15306, g16296;
wire g25271, g7133, g12464, g7846, g12797, I22794, I22845, g7803, g31950, g12292, g9461;
wire g12153, g25199, I22899, g8829, g11975, I12204, g19513, g23617, g15024, I20205, g12136;
wire I22719, g9904, g13143, I13453, I22718, g33394, g11169, I29315, I15168, g13884, g11410;
wire g23623, g9391, I15363, g8124, g24362, g11479, g23782, g13666, g13479, g8069, I32517;
wire g13217, g10622, g10566, g13478, I13565, I13464, g13486, g25258, g23266, g13580, g10653;
wire g14139, g16741, I14789, g23167, g13084, g28973, g14636, I14788, g14333, I17462, g21401;
wire g27796, g20236, g12796, g9654, g15867, g25337, g28934, g14664, g16196, g11676, g34545;
wire I22871, g11953, g13676, g23616, g29355, g15581, g10585, g9595, g23748, I14291, g11936;
wire I15334, g12192, g10609, I13109, g22940, I12097, g25425, g12522, g23809, g17744, I17447;
wire g28207, g17399, g14921, g15741, I32516, g9629, I13750, g14813, g11543, I12850, g13909;
wire g23733, g15735, g15877, g9800, g14674, g11117, g29025, g13000, I22754, g29540, g23630;
wire g22833, g15695, g25532, g15018, I13390, g14732, g24905, I15242, g19857, g17500, I15123;
wire g14761, I22844, g21555, g16854, g11974, g31671, g27933, g19549, g8806, g11639, g9823;
wire g12933, I25907, g10207, I20204, g26752, g14005, g16660, I26439, g17605, g11992, I29314;
wire I26438, I12096, I23962, I17446, g28206, g25309, I13564, I12730, g7857, g28758, I29269;
wire g14771, g8913, g11442, I13183, g14683, g17514, g25495, g12592, I13509, I14247, I15041;
wire g10515, I13851, g25985, g14882, g34424, g14407, g19856, I23951, I15340, g26255, g12152;
wire g22325, g13983, g16694, g17788, g12413, g10584, g28406, I13452, g28962, I29279, g28500;
wire g10759, g15721, I29278, I14766, I15130, I15193, I29286, g14758, g11130, g14082, g11193;
wire g13130, g14107, g16278, g12020, g19611, g23139, g16306, I12261, g14940, I18627, g13475;
wire g14848, g27282, g21415, g16815, g13727, g15734, g14804, g25255, I13731, g12357, g31978;
wire I22824, I15253, g24621, I18681, g14962, g13600, I22931, g9645, g23576, g19764, g11952;
wire I15175, I32757, I14370, g26782, g13821, g14048, I15264, g22755, g28421, g26352, I12271;
wire g13264, g24933, g13137, g13516, g15039, g29060, g17755, g13873, I31974, g14947, g10605;
wire g12482, g25470, g13834, g16321, g10951, g28920, g24574, g14234, g31706, I18626, g28946;
wire g25467, g23761, g23692, g27380, g12356, g9591, g12999, g11320, g25984, g19886, I15122;
wire g13346, g19792, I14957, g26053, g13464, g13797, g11292, I32756, g11153, g29094, g12449;
wire I14290, g11409, I22894, I14427, g14829, I31983, g14434, g29018, I12878, g10946, g28927;
wire g14946, g9750, I11826, g14344, g24583, I13182, I17496, g28903, g14682, g12149, I14481;
wire g28755, g12148, g13109, g16772, g24787, g29001, g13108, g12343, g13283, I22801, g11492;
wire g12971, I12545, g9528, g12369, g28395, I14956, g11381, g28899, I18529, g28990, g17220;
wire I15174, g29157, g17246, g12412, I26049, g26382, g33930, g22754, g33838, g14927, g16586;
wire I22866, g21345, g27582, g9372, g28861, I20461, g25476, g8359, g24662, I24461, g10604;
wire g15751, g10755, g24890, g14755, g19495, g27925, I22923, g29660, g20248, g16275, g14981;
wire I14211, g9334, g12112, I17923, g33306, g11326, g20081, g14794, g14845, I14497, I24365;
wire I13850, g13040, g13948, g14899, g29085, g28997, g25382, I12289, g14898, I32204, I23950;
wire g15014, I12288, g24380, g12429, g14521, I25221, g12428, g28871, I17885, g9908, g22902;
wire I16780, g10573, g9567, g14861, g14573, g24932, g15720, g11933, I14855, g14045, g29335;
wire g13634, g13851, g27317, I12374, g25215, g7850, g12317, g29694, g14098, g17699, g25439;
wire g28911, g23972, g17290, I29253, g29131, I15213, I12842, g25349, g12245, g12323, I14714;
wire g22661, I13730, g27775, g16236, I14257, g28950, I15051, I14818, g9724, g22715, I23120;
wire g24620, g14871, I12544, g13756, I18680, g12232, g16264, g19875, I22930, g26052, g26745;
wire g17572, g11350, I22965, I32433, g24369, g12512, g21359, g13846, g10472, g11396, I12270;
wire I14735, g19455, g20133, g17297, g21344, g11405, g15781, g20011, g14776, g28203, g10754;
wire g29015, g13929, I12219, g25200, g14825, g14950, g11020, g12080, g13928, I12218, g14858;
wire g19782, g29556, g31747, g14151, g14996, g24925, g24958, g17520, g12461, I24364, g12342;
wire I22937, I26395, I14923, g12145, g11302, I15105, I23980, g24944, g13105, I16779, I12470;
wire g9092, I16778, g19589, I12277, I13499, I17884, g15021, I12075, g27365, g24802, g29186;
wire g29676, g7690, g15726, I13498, g24793, g26235, g14058, I26440, g28895, I14885, g11881;
wire I14854, g25400, g12225, g14902, g12471, I29303, g12087, g14120, g14739, g10738, I22922;
wire I25845, g14146, g32072, g19466, I15003, g12244, g13248, I14480, g28376, g13779, I22685;
wire g27955, g28980, I23987, g23719, I12401, g28888, g28824, I20488, I22800, I22936, g11356;
wire g8691, g13945, g19874, g17581, g17315, g28931, I23969, g14547, g14895, g11998, I22762;
wire g13672, g12459, g16663, g10551, g21388, g24880, g23324, g14572, I14734, I20189, g21272;
wire I13043, I14993, I20188, g13513, g14127, g21462, g11961, g12079, g28860, g13897, I20460;
wire I24383, g12078, I26071, I15212, g14956, I11879, g14889, g16757, I11878, g28987, g25435;
wire I23979, g24989, g12159, g12125, I21978, I22974, I23978, g24988, g24924, I15149, g21360;
wire I23986, g27295, g20271, g11149, I15148, g28969, I26367, I26394, g12144, g9543, g13097;
wire g10520, g13104, g12336, g14520, I14187, g7150, I25220, g20199, g11971, g28870, g34048;
wire I13079, I13444, I32432, g14546, g14089, g22688, g20198, g17706, g17597, I12074, I13078;
wire g14088, g14024, g17689, I18589, g24528, g17624, g28867, I18588, g7836, I20467, I14169;
wire I14884, g11412, g15702, g13850, g15904, g25049, g12289, g14659, g14625, g14987, g20161;
wire g22885, g12023, g28910, g13896, I23917, g25048, g12224, g14943, I13336, g27687, g14968;
wire g11959, g13627, I22684, I20167, g14855, I12729, g13050, g13958, I12728, g28877, g20068;
wire I26366, I14531, g13742, g11944, g7620, g8010, I14186, g17287, g12195, g17596, g25514;
wire g24792, g17243, g12525, g12016, g23281, g21301, g21377, g14055, g17773, I18485, g14978;
wire g15780, I17475, g14590, g24918, g17670, g22839, g23699, I29302, g25473, g14741, g27705;
wire g22838, g17734, g28923, g16282, g9442, g27679, I15129, g12042, I15002, I26095, g12255;
wire g11002, I15128, g13057, g14735, g12188, g12124, I13392, g11245, I15299, g12460, g12686;
wire I20166, g11323, g14695, g14018, I15298, g11533, g21403, g20783, g12294, g17618, g28885;
wire g22306, I22873, I11865, I14230, g17468, I21993, g15787, g14706, I14992, g21385, I14510;
wire g15743, g21354, g14688, g28287, g12915, I13383, g11445, g14157, g22666, g13499, I13065;
wire g14066, g13498, I15080, g17363, g28942, g17217, g21190, g14876, g14885, g14854, g10511;
wire g11432, I23601, g13432, I14275, g12155, g12822, g15027, I15342, g28930, I24439, g28965;
wire g30573, I24438, g15710, g9715, g28131, g31509, g10916, I12241, g33933, g12589, g12194;
wire g10550, g13529, I14517, g12588, g27401, g12524, g23659, g11330, g13528, g13330, g10307;
wire I15365, g14085, g17740, g13764, g8238, g14596, g12119, g14054, I22711, g7701, g21339;
wire g13960, g32057, g12118, g12022, g21338, I26070, I17474, g16723, g14773, g24544, g13709;
wire g25389, g12285, I15087, g14655, g11708, g13708, g12053, g16097, I26094, I24415, I15043;
wire g13043, g14930, g14993, I17381, g24678, g14838, g14965, g22908, g13069, g29702, g34162;
wire g15717, I13401, g11955, g13955, g11970, g28410, g19962, g10618, I14351, g27693, I11864;
wire g34220, g28363, g17568, g14279, g7887, I13749, g13886, g7228, g11994, g15723, g23978;
wire g13967, I12345, I14790, I14516, g23590, I12849, g12008, g17814, g22638, I12848, g12476;
wire g13459, g21384, I23587, g8889, g14038, g23067, g10601, g13918, g16925, g14601, I18538;
wire g8871, I15079, g14677, I12263, g11545, g11444, g13079, I15078, g12239, g20201, g8500;
wire g14937, g26025, g13086, g16681, g17578, g12941, g19795, g12185, g21402, g17586, g11977;
wire g13977, I14530, g8737, g15011, g34227, g14015, g11561, g25172, I22872, g25996, g20170;
wire g10556, g13823, I13454, I21992, g14223, g17493, g15959, g27577, I15364, g12577, g14110;
wire g9246, g15742, I23586, g9203, g14740, I13382, I15289, g19358, I13519, g16299, g31003;
wire g14953, I15288, I13518, g12083, I15308, g11224, g13288, g15730, g14800, I24414, g29046;
wire g13495, I29261, g24809, I22846, g24808, I13729, g10587, g11374, g28391, g12415, g21287;
wire g19506, g10909, g20733, g21307, g15002, I25243, g13260, g14908, g10569, I22929, I15195;
wire I17405, I12344, g14569, g11489, g10568, g25895, g16316, g11559, g11424, I13566, g23655;
wire I29271, g9883, g14123, g15737, g14807, g19903, g12115, g14974, g17790, g17137, I13139;
wire g11544, g13544, g24570, g12052, g14638, I15042, I15255, I13852, g14841, g25385, g24567;
wire g11189, g11679, I23600, g29778, g13124, g25888, g31971, g23210, g16696, g20185, g10578;
wire g20675, g20092, g14014, g11938, g10586, g13093, g8873, g8632, g9538, I20221, I12240;
wire g9509, g23286, g25426, g29672, g17593, g14116, I32185, I14509, g10041, g14720, I32518;
wire g16259, I14508, g16225, g14041, g21187, I22710, g12207, g23975, g12539, I24463, g15753;
wire g12538, I12262, I13184, I14213, g15736, g17635, g16069, g13915, I22945, g14142, g33925;
wire g16657, I14205, g15843, g14517, g24906, g26714, g23666, I26417, g21363, I32439, g12100;
wire I17380, g24566, g22711, g14130, I18682, g17474, g28516, g11419, g29097, g15709, g27882;
wire g11155, I14350, g15708, g12414, g13822, g13266, g25527, I12098, g14727, I12251, I22717;
wire g17492, I17448, I15167, I15194, I17404, I31985, g21186, g23685, g7223, g14600, g14781;
wire g24576, g13119, g21417, g11118, g12114, g13118, g21334, g24609, g20200, I29295, g22663;
wire g33299, g23762, I15053, I15254, g27141, I25909, g24798, g14422, g24973, g20184, g23909;
wire I25908, g22757, g12332, g25019, g25018, I18633, g14542, g14021, g24934, I25242, g17757;
wire g10726, g23747, g10614, g27833, g12049, g10905, I15166, g14905, g12048, g20214, g28109;
wire g12221, g27613, g11892, g13892, g13476, g21416, I13141, I14249, I17379, I17925, I23949;
wire g14797, g27273, I14482, g16687, g13712, g17634, g11914, g17872, g12947, I14248, I22944;
wire g8728, I14204, g25300, g27463, g13907, g28381, g29057, g12463, g14136, g14408, g12972;
wire g28174, g28796, g31753, I22793, g16260, g7823, g28840, g11382, I15176, I12203, g19632;
wire I24440, g11675, g13176, g13092, g26269, g34550, g11154, g29737, g28522, g8678, g17592;
wire g16893, g10537, I14331, g8105, I31984, g16713, I20462, I29255, I24462, g17820, g31709;
wire g15752, I29270, g28949, I13463, g31708, g17846, g17396, g14750, g24584, I14212, g7167;
wire g10796, g20107, g11906, I12403, g16093, g12344, g13083, I32441, g13284, g7549, g25341;
wire g29722, g25268, g16875, g7598, I32758, g14663, g24804, g24652, g13139, g15713, I14369;
wire g34469, I15333, g19546, g8227, I14368, g12028, g15042, g21253, I29277, g23781, g13963;
wire g17640, I14229, g21351, g26666, I14228, g15030, g27903, g13554, I17924, g12491, g28780;
wire I22753, g11312, g11200, g25038, g13115, I15052, g14933, I14925, g16155, g17662, g28820;
wire I12546, I17461, g14851, g27767, g9775, g20371, g24951, g24972, g12767, g13798, g11973;
wire g30580, g29657, g17779, g11674, g7879, g23726, I20203, g16524, g26685, I14429, g14574;
wire g12191, g14452, g11934, g16119, I14428, g12521, g17647, I29313, g8609, g19450, I14765;
wire g11761, g22651, I29285, g14051, g14072, g16749, g20163, g15782, I29254, I15214, g14780;
wire g12045, g10820, g14820, g17513, g28827, g25531, g15853, I15241, g12462, g13241, g25186;
wire g14691, g25953, g8803, g9954, I22792, I22967, g13100, g23575, g20173, g10929, g31669;
wire g15864, g33669, g25334, g17723, g10583, g10928, g15748, g21283, g9912, I13045, g20134;
wire g13515, g13882, g24760, I23961, g25216, g14113, I24385, g15036, g19597, g12629, I12877;
wire I13462, g8847, g12628, g22850, g11441, I13140, I22901, g28786, g11206, g16238, I14499;
wire g17412, I18625, g14768, g28945, g14803, I14498, g33679, g12147, I12402, I15107, I22823;
wire I14611, I14924, g12370, g25974, g17716, g15008, I23971, g25293, g12151, g19854, g13940;
wire I22966, g23949, g28448, I15263, g10552, g8751, g15907, g22681, g11135, I14330, g19916;
wire g16728, g12227, I14764, g11962, I29284, I31973, I29304, I18581, I26051, I25847, I26072;
wire I11825, I12876, g14999, g16304, g12044, I15004, g21509, g17765, I14259, I17495, g27377;
wire g24926, g25275, g12301, I14258, g12120, g27738, I32440, g25237, I15106, g13273, g19335;
wire g10961, g29679, g15729, g14505, I12287, I14955, g19965, g11951, g15728, g13951, I12076;
wire g23047, g13795, g28896, I14171, g20871, I22893, I12269, I13044, g17775, I22865, g23756;
wire g14723, g23780, g14433, I24384, g21350, g16312, g14104, I25846, g14343, g10971, g28958;
wire g14971, g16745, g31748, g26208, g16813, I22938, g27824, g13920, I17460, g24591, g24776;
wire I14817, g25236, I15121, g34422, g28857, g14133, I12279, I14532, g13121, g28793, I13403;
wire I12278, g24950, I12469, g27931, g28765, g7611, g14011, g20151, g20172, I12468, g13291;
wire g11173, g12190, g22753, g28504, g21357, g31009, g14627, g23357, g14959, g14379, g22650;
wire g11134, g23105, g13134, g14378, g7209, g12024, g17650, g10603, g17736, g15798, g25021;
wire I11824, g15674, g9310, I14289, g28298, g9663, g13927, I17494, g29118, I12217, g14730;
wire g22709, I22822, g13240, g24957, g11491, g12644, g11903, I14816, I32203, g23890, g12969;
wire I13520, g20645, g28856, g14548, g17225, g17708, g12197, g8434, g28512, g23552, g15005;
wire g14317, g12411, g8347, I15262, g23778, g11395, I13497, g11990, g13990, g23786, I18487;
wire g13898, I22864, g21356, I12373, g14626, g24661, g24547, I31972, g12450, g10775, g9295;
wire g12819, g12910, g34174, g17792, I22900, g10737, g25537, g12111, g28271, g13861, g21331;
wire g13573, g23932, I14713, g12590, g33083, g11389, g25492, g14697, g9966, g7184, g9705;
wire I14610, I26368, I29263, g11534, I23602, g20784, g28736, g19265, g13098, I20487, g11251;
wire g25381, I23970, g13462, g28843, g19510, g20181, g12019, g17598, g12196, g11997, I20469;
wire I21994, I12242, g12526, g15725, I20468, g29154, g21433, I22892, g19442, g12402, g10611;
wire I13111, g13871, I23919, I18486, g28259, g14924, I22712, g17656, I20187, g15744, I17476;
wire I23918, I18580, I26050, I13384, g12001, I13067, I12841, I11877, g10529, g13628, g23850;
wire g13911, I18531, g17364, g28955, I14277, I21977, g14696, I24363, g8163, g15962, g14764;
wire g11591, g21011, I15147, g12066, I20486, g24943, g20644, g27876, g15833, I13402, g11355;
wire g28994, g14868, g17571, I11866, g27854, g25062, I20223, g16507, g11858, I14352, I17883;
wire g11172, g12511, g22687, g7885, g11996, g17495, g23379, I14170, I13077, g23112, g20870;
wire g17816, g14258, g11394, g22643, g34051, g21386, I18587, g21603, I14853, g27550, g9485;
wire g14069, g22668, g10602, g11446, g14810, g15033, g12287, g21429, g17669, g12307, g14879;
wire I13066, g17668, g23428, g13058, g28977, g12431, g20979, g28783, g20055, g20111, g17525;
wire I13511, g12341, g28823, I14276, I21976, g16291, I23985, g13281, g27670, g22713, g11957;
wire g28336, I32202, g13739, g25396, g28966, g14918, g20150, g14079, g17705, g8292, g14599;
wire I12253, g17679, g7869, g10598, g15788, I18579, g14598, I14733, g15829, g17686, I12372;
wire g14817, g28288, g19913, g19614, g22875, g25020, g7442, g24917, g10561, g27468, I22921;
wire g27306, g19530, g12286, g14656, g9177, g22837, g12306, I26461, I24416, g16604, I22799;
wire g13551, g10336, g28976, I14712, I13335, g16770, g8561, I22973, g26248, g12187, I29262;
wire g11490, I26393, g30249, g33141, g13824, g27479, g12479, g20854, g33135, g7675, g12486;
wire g9694, g8906, g14816, g12223, g14687, g14752, g16272, g22524, g25778, g26212, g17194;
wire g14392, g13700, g11658, g15718, g10488, g29107, g10893, g25932, g29141, g14713, g31507;
wire g15099, g11527, g32715, g15098, g30148, g23602, g28470, g16220, g14679, g23955, g33163;
wire g24619, g14188, g14124, g14678, g16246, g12117, g29361, g15140, g14093, g15061, g13910;
wire g13202, g12123, g27772, g12772, g31121, g23918, g15162, g11384, g23079, g29106, g13094;
wire g26603, g29033, g15628, g32520, g17239, g31134, g33134, g16227, g27007, g31506, g15071;
wire g15147, g15754, g14037, g15825, g16044, g27720, g14419, g29012, g15151, g14418, g10266;
wire g25958, g32296, g31491, g11280, g25944, g29359, g12806, g14194, g19413, g24953, g15059;
wire g26298, g30129, g15058, g11231, g17284, g12193, g11885, g29173, g14313, g28476, g16226;
wire g11763, g25504, g15120, g32910, g25317, g10808, g15146, g14036, g34737, g12437, g27703;
wire g20000, g13480, g14642, g12347, g14064, g13076, g33098, g28519, g12821, g27063, g24751;
wire g29903, g11773, g27516, g33140, g13341, g12137, g13670, g10555, g20841, g23042, g14712;
wire g13335, g19890, g14914, g24391, g15127, g30271, g23124, g23678, g16024, g12208, g33447;
wire g26330, g23686, g20014, g33162, g29898, g12453, g15095, g29191, g19778, g11618, g14382;
wire g14176, g14092, g19999, g22400, g20720, g11469, g12593, g12346, g24720, g11039, g11306;
wire g30132, g22539, g8958, g33147, g9061, g19932, g25887, g15089, g15088, g13937, g21277;
wire g29032, g15126, g11666, g16581, g11363, g11217, g31318, g12711, g8177, g30171, g17515;
wire g15060, g12492, g26545, g27982, g27381, g14415, g13110, g26598, g33146, g29071, g29370;
wire g33427, g22399, g10312, g15055, g15070, g30159, g23560, g12483, g11216, g10799, g12553;
wire g23642, g15067, g15094, g30144, g24453, g15150, g31127, g13908, g12252, g26309, g11747;
wire g13568, g16066, g16231, g33103, g19793, g33095, g12847, g25144, g13772, g28515, g28414;
wire g30288, g26976, g29146, g12851, g14539, g9649, g14538, g28584, g16287, g33089, g15102;
wire g15157, g33088, g22514, g12311, g15066, g24575, g30260, g23883, g26865, g31126, g16268;
wire g12780, g14515, g14414, g11493, g25954, g23729, g20982, g19880, g27731, g12846, g22535;
wire g13806, g29889, g26686, g13517, g20390, g29181, g21284, g26267, g12405, g16210, g15054;
wire g27046, g15156, g30294, g12046, g14399, g11006, g12113, g28106, g25189, g27827, g9586;
wire g19887, g29497, g27769, g15131, g27768, g30160, g33094, g14361, g20183, g28514, g22491;
wire g16479, g27027, g24508, g23052, g12662, g25160, g12249, g11834, g12204, g15143, g30170;
wire g29503, g14033, g12081, g13021, g22521, g27647, g11913, g13913, g27356, g7601, g15168;
wire g27826, g29910, g11607, g14514, g11346, g29070, g12651, g10421, g30119, g14163, g11797;
wire g19919, g30276, g30285, g19444, g12505, g27717, g9100, g12026, g8984, g14121, g25022;
wire g11891, g16242, g28491, g33085, g14291, g11537, g27343, g28981, g29077, g12646, g11283;
wire g10760, g11303, g31942, g27368, g21206, g12850, g13796, g28521, g31965, g33131, g12228;
wire g10649, g12716, g15123, g10491, g20027, g21652, g27379, g11483, g31469, g11862, g12050;
wire g24779, g16237, g29916, g23135, g15992, g28462, g13326, g14767, g14395, g17420, g10899;
wire g22540, g11252, g11621, g15578, g20998, g33143, g7661, g29180, g14247, g13872, g25501;
wire g20717, g14272, g12129, g12002, g11213, g15142, g33084, g20149, g26609, g15130, g24148;
wire g15165, g31373, g11780, g14360, g9835, g14447, g12856, g29187, g11846, g16209, g14911;
wire g27499, g28540, g15372, g14754, g27722, g31117, g27924, g33117, g22190, g8720, g15063;
wire g30934, g19984, g15137, g12432, g24959, g17190, g14394, g14367, g16292, g11357, g29179;
wire g14420, g12198, g19853, g27528, g10318, g14446, g14227, g20857, g27960, g14540, g19401;
wire g17700, g17625, g15073, g28481, g10281, g15122, g26515, g12708, g25005, g10699, g15153;
wire g31116, g11248, g32780, g15136, g29908, g27879, g22450, g12970, g27878, g27337, g15164;
wire g11945, g11999, g10715, g21389, g20995, g28520, g25407, g27010, g11932, g33130, g11448;
wire g14490, g19907, g21140, g15091, g33437, g29007, g10671, g14181, g23871, g27353, g16183;
wire g27823, g11148, g12680, g19935, g31372, g25141, g33175, g24145, g27966, g13971, g29035;
wire g14211, g27364, g33137, g12017, g12364, g30613, g29142, g14497, g30273, g30106, g12288;
wire g29193, g19906, g12571, g12308, g25004, g28496, g29165, g14339, g16072, g10338, g15062;
wire g28986, g29006, g25947, g15508, g13959, g27954, g12752, g11958, g12374, g13378, g14411;
wire g13603, g13944, g14867, g14450, g29175, g10819, g13730, g34359, g14707, g28457, g32212;
wire g12558, g13765, g15051, g15072, g7192, g29873, g17180, g22993, g14094, g15152, g33109;
wire g12189, g13129, g10801, g17694, g33108, g30134, g11626, g10695, g27093, g17619, g12093;
wire g26649, g27875, g33174, g11232, g29034, g19400, g21127, g11697, g11995, g16027, g11261;
wire g14001, g30240, g24631, g12160, g13512, g28480, g23956, g8933, g31483, g13831, g12201;
wire g29164, g12467, g30262, g13989, g13056, g16090, g26573, g11924, g29109, g27352, g26247;
wire g7781, g12419, g25770, g29108, g24976, g12418, g12170, g26098, g23024, g13342, g13031;
wire g12853, g33851, g29174, g21250, g21658, g22654, g25521, g11869, g15647, g28469, g15090;
wire g28468, g10341, g25247, g27704, g11225, g26162, g16646, g12466, g25777, g14335, g12101;
wire g26628, g29040, g30162, g8864, g24383, g27733, g13970, g11171, g29183, g24875, g12166;
wire g14278, g13994, g15149, g25447, g14306, g29933, g15148, g15097, g30147, g13919, g9755;
wire g13078, g23695, g19951, g25776, g25785, g10884, g27382, g28953, g24494, g15133, g32650;
wire g13125, g10666, g25950, g7142, g12154, g29072, g9602, g14556, g26645, g13336, g21256;
wire g22983, g9015, g15050, g12729, g13631, g10922, g25446, g22517, g10179, g9664, g15096;
wire g30146, g25540, g14178, g31482, g30290, g28568, g25203, g11309, g11571, g22523, g14417;
wire g12622, g26715, g23763, g14334, g16232, g11976, g33090, g31233, g17727, g11954, g13954;
wire g28510, g12333, g26297, g15129, g12852, g15057, g11669, g15128, g14000, g33449, g33448;
wire g14568, g17175, g10123, g21655, g34354, g12609, g14751, g14772, g8182, g28493, g26546;
wire g19981, g28340, g14416, g11610, g25784, g27973, g33148, g25956, g11255, g33097, g14391;
wire g12798, g10510, g11270, g16198, g7352, g26625, g27732, g13939, g32017, g26296, g26338;
wire g15056, g27400, g10615, g31133, g33133, g28475, g21143, g19388, g15145, g24439, g9700;
wire g11201, g33112, g27771, g19140, g19997, g15132, g12235, g33096, g14362, g22537, g15161;
wire g14165, g29104, g12515, g15087, g32424, g34496, g14437, g11194, g15069, g14347, g14253;
wire g15068, g17174, g34067, g11119, g30150, g33129, g10821, g12435, g33128, g14821, g22522;
wire g11313, g27345, g12744, g14516, g11276, g12849, g17663, g12848, g27652, g26256, g22536;
wire g15086, g12361, g14726, g30280, g32455, g15159, g16288, g14320, g15158, g30157, g14122;
wire g15144, g31498, g28492, g8086, g11907, g33432, g26314, g12371, g23835, g11238, g17213;
wire g12234, g23586, g33145, g14164, g11185, g13518, g16488, g16424, g26268, g14575, g11935;
wire g8131, g27012, g13883, g33132, g12163, g28483, g26993, g33161, g26667, g30156, g11729;
wire g13501, g27829, g14091, g27828, g22405, g15669, g12358, g27344, g12121, g21193, g22929;
wire g31068, g11566, g13622, g31970, g12173, g28509, g16219, g14522, g11653, g22357, g29145;
wire g12029, g10862, g11415, g29198, g13852, g30601, g28452, g27927, g16201, g15093, g30143;
wire g23063, g15065, g30169, g14397, g12604, g27770, g19338, g12755, g33125, g21209, g14872;
wire g19968, g23208, g15160, g13799, g17482, g33144, g33823, g20234, g29069, g11184, g7158;
wire g10205, g24514, g30922, g29886, g11692, g16313, g27926, g13013, g19070, g22513, g15155;
wire g11207, g15170, g22448, g13539, g13005, g25321, g14396, g14731, g15167, g14413, g28803;
wire g11771, g25800, g27766, g23711, g30117, g29144, g19402, g23108, g17148, g11414, g16476;
wire g32585, g15053, g28482, g30123, g27629, g28552, g15101, g12246, g11584, g30265, g14640;
wire g15064, g10803, g12591, g12785, g27355, g13114, g27825, g11435, g11107, g15166, g12858;
wire g11345, g33093, g31294, g11940, g27367, g14027, g11804, g15570, g14248, g16215, g24990;
wire g14003, g15074, g12318, g27059, g15594, g12059, g12025, g33160, g12540, g13500, g15092;
wire g28149, g15154, g21062, g14090, g13004, g33075, g19268, g12377, g12739, g30130, g24701;
wire g12146, g12645, g13947, g11273, g14513, g29705, g14449, g29189, g33419, g14448, g11972;
wire g27366, g7567, g14212, g12632, g24766, g23051, g34703, g11514, g12226, g31119, g26873;
wire g11012, g15139, g26209, g15138, g11473, g29915, g27354, g12297, g13325, g12980, g12824;
wire g25952, g13946, g25175, g14228, g15585, g26346, g15608, g15052, g12211, g31008, g31476;
wire g29167, g17198, g27659, g17393, g12700, g12659, g12126, g30136, g19953, g10793, g14793;
wire g27338, g12296, g9762, g23662, g27969, g14549, g11755, g29900, g33092, g11563, g12855;
wire g31935, g23204, g14002, g17657, g11191, g28498, g15100, g12581, g33439, g7175, g33438;
wire g7139, g22545, g28031, g12067, g14512, g27735, g27877, g28529, g12150, g33139, g10831;
wire g13032, g33138, g14445, g12695, g29675, g26183, g30252, g7304, g14611, g7499, g14988;
wire g11360, g26872, g14271, g30183, g19430, g15141, g14145, g12256, g25948, g24497, g14529;
wire g27102, g15135, g26574, g14393, g14365, g32845, g17309, g15049, g11950, g10709, g27511;
wire g12854, g28425, g34912, g25851, g13996, g28444, g15106, g17954, g12550, g12314, g14602;
wire g27721, g12085, g22488, g14337, g11203, g13044, g14792, g28353, g29200, g9640, g19063;
wire g33100, g13377, g14425, g27734, g15163, g30929, g19873, g10918, g19422, g14444, g12667;
wire g19209, g13698, g31515, g29184, g23626, g15724, g24018, g30282, g19453, g15121, g12443;
wire g19436, g13661, g11715, g29005, g33107, g12601, g15134, g14364, g25769, g11385;
wire line1, line2, line3, line4, line5, line6, line7, line8, line9, line10, line11;
wire line12, line13, line14, line15, line16, line17, line18, line19, line20, line21, line22;
wire line23, line24, line25, line26, line27, line28, line29, line30, line31, line32, line33;
wire line34, line35, line36, line37, line38, line39, line40, line41, line42, line43, line44;
wire line45, line46, line47, line48, line49, line50, line51, line52, line53, line54, line55;
wire line56, line57, line58, line59, line60, line61, line62, line63, line64, line65, line66;
wire line67, line68, line69, line70, line71, line72, line73, line74, line75, line76, line77;
wire line78, line79, line80, line81, line82, line83, line84, line85, line86, line87, line88;
wire line89, line90, line91, line92, line93, line94, line95, line96, line97, line98, line99;
wire line100, line101, line102, line103, line104, line105, line106, line107, line108, line109, line110;
wire line111, line112, line113, line114, line115, line116, line117, line118, line119, line120, line121;
wire line122, line123, line124, line125, line126, line127, line128, line129, line130, line131, line132;
wire line133, line134, line135, line136, line137, line138, line139, line140, line141, line142, line143;
wire line144, line145, line146, line147, line148, line149, line150, line151, line152, line153, line154;
wire line155, line156, line157, line158, line159, line160, line161, line162, line163, line164, line165;
wire line166, line167, line168, line169, line170, line171, line172, line173, line174, line175, line176;
wire line177, line178, line179, line180, line181, line182, line183, line184, line185, line186, line187;
wire line188, line189, line190, line191, line192, line193, line194, line195, line196, line197, line198;
wire line199, line200, line201, line202, line203, line204, line205, line206, line207, line208, line209;
wire line210, line211, line212, line213, line214, line215, line216, line217, line218, line219, line220;
wire line221, line222, line223, line224, line225, line226, line227, line228, line229, line230, line231;
wire line232, line233, line234, line235, line236, line237, line238, line239, line240, line241, line242;
wire line243, line244, line245, line246, line247, line248, line249, line250, line251, line252, line253;
wire line254, line255, line256, line257, line258, line259, line260, line261, line262, line263, line264;
wire line265, line266, line267, line268, line269, line270, line271, line272, line273, line274, line275;
wire line276, line277, line278, line279, line280, line281, line282, line283, line284, line285, line286;
wire line287, line288, line289, line290, line291, line292, line293, line294, line295, line296, line297;
wire line298, line299, line300, line301, line302, line303, line304, line305, line306, line307, line308;
wire line309, line310, line311, line312, line313, line314, line315, line316, line317, line318, line319;
wire line320, line321, line322, line323, line324, line325, line326, line327, line328, line329, line330;
wire line331, line332, line333, line334, line335, line336, line337, line338, line339, line340, line341;
wire line342, line343, line344, line345, line346, line347, line348, line349, line350, line351, line352;
wire line353, line354, line355, line356, line357, line358, line359, line360, line361, line362, line363;
wire line364, line365, line366, line367, line368, line369, line370, line371, line372, line373, line374;
wire line375, line376, line377, line378, line379, line380, line381, line382, line383, line384, line385;
wire line386, line387, line388, line389, line390, line391, line392, line393, line394, line395, line396;
wire line397, line398, line399, line400, line401, line402, line403, line404, line405, line406, line407;
wire line408, line409, line410, line411, line412, line413, line414, line415, line416, line417, line418;
wire line419, line420, line421, line422, line423, line424, line425, line426, line427, line428, line429;
wire line430, line431, line432, line433, line434, line435, line436, line437, line438, line439, line440;
wire line441, line442, line443, line444, line445, line446, line447, line448, line449, line450, line451;
wire line452, line453, line454, line455, line456, line457, line458, line459, line460, line461, line462;
wire line463, line464, line465, line466, line467, line468, line469, line470, line471, line472, line473;
wire line474, line475, line476, line477, line478, line479, line480, line481, line482, line483, line484;
wire line485, line486, line487, line488, line489, line490, line491, line492, line493, line494, line495;
wire line496, line497, line498, line499, line500, line501, line502, line503, line504, line505, line506;
wire line507, line508, line509, line510, line511, line512, line513, line514, line515, line516, line517;
wire line518, line519, line520, line521, line522, line523, line524, line525, line526, line527, line528;
wire line529, line530, line531, line532, line533, line534, line535, line536, line537, line538, line539;
wire line540, line541, line542, line543, line544, line545, line546, line547, line548, line549, line550;
wire line551, line552, line553, line554, line555, line556, line557, line558, line559, line560, line561;
wire line562, line563, line564, line565, line566, line567, line568, line569, line570, line571, line572;
wire line573, line574, line575, line576, line577, line578, line579, line580, line581, line582, line583;
wire line584, line585, line586, line587, line588, line589, line590, line591, line592, line593, line594;
wire line595, line596, line597, line598, line599, line600, line601, line602, line603, line604, line605;
wire line606, line607, line608, line609, line610, line611, line612, line613, line614, line615, line616;
wire line617, line618, line619, line620, line621, line622, line623, line624, line625, line626, line627;
wire line628, line629, line630, line631, line632, line633, line634, line635, line636, line637, line638;
wire line639, line640, line641, line642, line643, line644, line645, line646, line647, line648, line649;
wire line650, line651, line652, line653, line654, line655, line656, line657, line658, line659, line660;
wire line661, line662, line663, line664, line665, line666, line667, line668, line669, line670, line671;
wire line672, line673, line674, line675, line676, line677, line678, line679, line680, line681, line682;
wire line683, line684, line685, line686, line687, line688, line689, line690, line691, line692, line693;
wire line694, line695, line696, line697, line698, line699, line700, line701, line702, line703, line704;
wire line705, line706, line707, line708, line709, line710, line711, line712, line713, line714, line715;
wire line716, line717, line718, line719, line720, line721, line722, line723, line724, line725, line726;
wire line727, line728, line729, line730, line731, line732, line733, line734, line735, line736, line737;
wire line738, line739, line740, line741, line742, line743, line744, line745, line746, line747, line748;
wire line749, line750, line751, line752, line753, line754, line755, line756, line757, line758, line759;
wire line760, line761, line762, line763, line764, line765, line766, line767, line768, line769, line770;
wire line771, line772, line773, line774, line775, line776, line777, line778, line779, line780, line781;
wire line782, line783, line784, line785, line786, line787, line788, line789, line790, line791, line792;
wire line793, line794, line795, line796, line797, line798, line799, line800, line801, line802, line803;
wire line804, line805, line806, line807, line808, line809, line810, line811, line812, line813, line814;
wire line815, line816, line817, line818, line819, line820, line821, line822, line823, line824, line825;
wire line826, line827, line828, line829, line830, line831, line832, line833, line834, line835, line836;
wire line837, line838, line839, line840, line841, line842, line843, line844, line845, line846, line847;
wire line848, line849, line850, line851, line852, line853, line854, line855, line856, line857, line858;
wire line859, line860, line861, line862, line863, line864, line865, line866, line867, line868, line869;
wire line870, line871, line872, line873, line874, line875, line876, line877, line878, line879, line880;
wire line881, line882, line883, line884, line885, line886, line887, line888, line889, line890, line891;
wire line892, line893, line894, line895, line896, line897, line898, line899, line900, line901, line902;
wire line903, line904, line905, line906, line907, line908, line909, line910, line911, line912, line913;
wire line914, line915, line916, line917, line918, line919, line920, line921, line922, line923, line924;
wire line925, line926, line927, line928, line929, line930, line931, line932, line933, line934, line935;
wire line936, line937, line938, line939, line940, line941, line942, line943, line944, line945, line946;
wire line947, line948, line949, line950, line951, line952, line953, line954, line955, line956, line957;
wire line958, line959, line960, line961, line962, line963, line964, line965, line966, line967, line968;
wire line969, line970, line971, line972, line973, line974, line975, line976, line977, line978, line979;
wire line980, line981, line982, line983, line984, line985, line986, line987, line988, line989, line990;
wire line991, line992, line993, line994, line995, line996, line997, line998, line999, line1000, line1001;
wire line1002, line1003, line1004, line1005, line1006, line1007, line1008, line1009, line1010, line1011, line1012;
wire line1013, line1014, line1015, line1016, line1017, line1018, line1019, line1020, line1021, line1022, line1023;
wire line1024, line1025, line1026, line1027, line1028, line1029, line1030, line1031, line1032, line1033, line1034;
wire line1035, line1036, line1037, line1038, line1039, line1040, line1041, line1042, line1043, line1044, line1045;
wire line1046, line1047, line1048, line1049, line1050, line1051, line1052, line1053, line1054, line1055, line1056;
wire line1057, line1058, line1059, line1060, line1061, line1062, line1063, line1064, line1065, line1066, line1067;
wire line1068, line1069, line1070, line1071, line1072, line1073, line1074, line1075, line1076, line1077, line1078;
wire line1079, line1080, line1081, line1082, line1083, line1084, line1085, line1086, line1087, line1088, line1089;
wire line1090, line1091, line1092, line1093, line1094, line1095, line1096, line1097, line1098, line1099, line1100;
wire line1101, line1102, line1103, line1104, line1105, line1106, line1107, line1108, line1109, line1110, line1111;
wire line1112, line1113, line1114, line1115, line1116, line1117, line1118, line1119, line1120, line1121, line1122;
wire line1123, line1124, line1125, line1126, line1127, line1128, line1129, line1130, line1131, line1132, line1133;
wire line1134, line1135, line1136, line1137, line1138, line1139, line1140, line1141, line1142, line1143, line1144;
wire line1145, line1146, line1147, line1148, line1149, line1150, line1151, line1152, line1153, line1154, line1155;
wire line1156, line1157, line1158, line1159, line1160, line1161, line1162, line1163, line1164, line1165, line1166;
wire line1167, line1168, line1169, line1170, line1171, line1172, line1173, line1174, line1175, line1176, line1177;
wire line1178, line1179, line1180, line1181, line1182, line1183, line1184, line1185, line1186, line1187, line1188;
wire line1189, line1190, line1191, line1192, line1193, line1194, line1195, line1196, line1197, line1198, line1199;
wire line1200, line1201, line1202, line1203, line1204, line1205, line1206, line1207, line1208, line1209, line1210;
wire line1211, line1212, line1213, line1214, line1215, line1216, line1217, line1218, line1219, line1220, line1221;
wire line1222, line1223, line1224, line1225, line1226, line1227, line1228, line1229, line1230, line1231, line1232;
wire line1233, line1234, line1235, line1236, line1237, line1238, line1239, line1240, line1241, line1242, line1243;
wire line1244, line1245, line1246, line1247, line1248, line1249, line1250, line1251, line1252, line1253, line1254;
wire line1255, line1256, line1257, line1258, line1259, line1260, line1261, line1262, line1263, line1264, line1265;
wire line1266, line1267, line1268, line1269, line1270, line1271, line1272, line1273, line1274, line1275, line1276;
wire line1277, line1278, line1279, line1280, line1281, line1282, line1283, line1284, line1285, line1286, line1287;
wire line1288, line1289, line1290, line1291, line1292, line1293, line1294, line1295, line1296, line1297, line1298;
wire line1299, line1300, line1301, line1302, line1303, line1304, line1305, line1306, line1307, line1308, line1309;
wire line1310, line1311, line1312, line1313, line1314, line1315, line1316, line1317, line1318, line1319, line1320;
wire line1321, line1322, line1323, line1324, line1325, line1326, line1327, line1328, line1329, line1330, line1331;
wire line1332, line1333, line1334, line1335, line1336, line1337, line1338, line1339, line1340, line1341, line1342;
wire line1343, line1344, line1345, line1346, line1347, line1348, line1349, line1350, line1351, line1352, line1353;
wire line1354, line1355, line1356, line1357, line1358, line1359, line1360, line1361, line1362, line1363, line1364;
wire line1365, line1366, line1367, line1368, line1369, line1370, line1371, line1372, line1373, line1374, line1375;
wire line1376, line1377, line1378, line1379, line1380, line1381, line1382, line1383, line1384, line1385, line1386;
wire line1387, line1388, line1389, line1390, line1391, line1392, line1393, line1394, line1395, line1396, line1397;
wire line1398, line1399, line1400, line1401, line1402, line1403, line1404, line1405, line1406, line1407, line1408;
wire line1409, line1410, line1411, line1412, line1413, line1414, line1415, line1416, line1417, line1418, line1419;
wire line1420, line1421, line1422, line1423, line1424, line1425, line1426;
DFFX1 gate1(.Q (g5057), .QB (line1), .D(g33046), .CK(clk));
DFFX1 gate2(.Q (g2771), .QB (line2), .D(g34441), .CK(clk));
DFFX1 gate3(.Q (g1882), .QB (line3), .D(g33982), .CK(clk));
DFFX1 gate4(.Q (g6462), .QB (line4), .D(g25751), .CK(clk));
DFFX1 gate5(.Q (g2299), .QB (line5), .D(g34007), .CK(clk));
DFFX1 gate6(.Q (g4040), .QB (line6), .D(g24276), .CK(clk));
DFFX1 gate7(.Q (g2547), .QB (line7), .D(g30381), .CK(clk));
DFFX1 gate8(.Q (g559), .QB (line8), .D(g640), .CK(clk));
DFFX1 gate9(.Q (g3017), .QB (line9), .D(g31877), .CK(clk));
DFFX1 gate10(.Q (g3243), .QB (line10), .D(g30405), .CK(clk));
DFFX1 gate11(.Q (g452), .QB (line11), .D(g25604), .CK(clk));
DFFX1 gate12(.Q (g464), .QB (line12), .D(g25607), .CK(clk));
DFFX1 gate13(.Q (g3542), .QB (line13), .D(g30416), .CK(clk));
DFFX1 gate14(.Q (g5232), .QB (line14), .D(g30466), .CK(clk));
DFFX1 gate15(.Q (g5813), .QB (line15), .D(g25736), .CK(clk));
DFFX1 gate16(.Q (g2907), .QB (line16), .D(g34617), .CK(clk));
DFFX1 gate17(.Q (g1744), .QB (line17), .D(g33974), .CK(clk));
DFFX1 gate18(.Q (g5909), .QB (line18), .D(g30505), .CK(clk));
DFFX1 gate19(.Q (g1802), .QB (line19), .D(g33554), .CK(clk));
DFFX1 gate20(.Q (g3554), .QB (line20), .D(g30432), .CK(clk));
DFFX1 gate21(.Q (g6219), .QB (line21), .D(g33064), .CK(clk));
DFFX1 gate22(.Q (g807), .QB (line22), .D(g34881), .CK(clk));
DFFX1 gate23(.Q (g6031), .QB (line23), .D(g6027), .CK(clk));
DFFX1 gate24(.Q (g847), .QB (line24), .D(g24216), .CK(clk));
DFFX1 gate25(.Q (g976), .QB (line25), .D(g24232), .CK(clk));
DFFX1 gate26(.Q (g4172), .QB (line26), .D(g34733), .CK(clk));
DFFX1 gate27(.Q (g4372), .QB (line27), .D(g34882), .CK(clk));
DFFX1 gate28(.Q (g3512), .QB (line28), .D(g33026), .CK(clk));
DFFX1 gate29(.Q (g749), .QB (line29), .D(g31867), .CK(clk));
DFFX1 gate30(.Q (g3490), .QB (line30), .D(g25668), .CK(clk));
DFFX1 gate31(.Q (g6005), .QB (line31), .D(g24344), .CK(clk));
DFFX1 gate32(.Q (g4235), .QB (line32), .D(g4232), .CK(clk));
DFFX1 gate33(.Q (g1600), .QB (line33), .D(g33966), .CK(clk));
DFFX1 gate34(.Q (g1714), .QB (line34), .D(g33550), .CK(clk));
DFFX1 gate35(.Q (g3649), .QB (line35), .D(g3625), .CK(clk));
DFFX1 gate36(.Q (g3155), .QB (line36), .D(g30393), .CK(clk));
DFFX1 gate37(.Q (g3355), .QB (line37), .D(g31880), .CK(clk));
DFFX1 gate38(.Q (g2236), .QB (line38), .D(g29248), .CK(clk));
DFFX1 gate39(.Q (g4555), .QB (line39), .D(g4571), .CK(clk));
DFFX1 gate40(.Q (g3698), .QB (line40), .D(g24274), .CK(clk));
DFFX1 gate41(.Q (g6073), .QB (line41), .D(g31920), .CK(clk));
DFFX1 gate42(.Q (g1736), .QB (line42), .D(g33973), .CK(clk));
DFFX1 gate43(.Q (g1968), .QB (line43), .D(g30360), .CK(clk));
DFFX1 gate44(.Q (g4621), .QB (line44), .D(g34460), .CK(clk));
DFFX1 gate45(.Q (g5607), .QB (line45), .D(g30494), .CK(clk));
DFFX1 gate46(.Q (g2657), .QB (line46), .D(g30384), .CK(clk));
DFFX1 gate47(.Q (g5659), .QB (line47), .D(g24340), .CK(clk));
DFFX1 gate48(.Q (g490), .QB (line48), .D(g29223), .CK(clk));
DFFX1 gate49(.Q (g311), .QB (line49), .D(g26881), .CK(clk));
DFFX1 gate50(.Q (g6069), .QB (line50), .D(g31925), .CK(clk));
DFFX1 gate51(.Q (g772), .QB (line51), .D(g34252), .CK(clk));
DFFX1 gate52(.Q (g5587), .QB (line52), .D(g30489), .CK(clk));
DFFX1 gate53(.Q (g6177), .QB (line53), .D(g29301), .CK(clk));
DFFX1 gate54(.Q (g6377), .QB (line54), .D(g6373), .CK(clk));
DFFX1 gate55(.Q (g3167), .QB (line55), .D(g33022), .CK(clk));
DFFX1 gate56(.Q (g5615), .QB (line56), .D(g30496), .CK(clk));
DFFX1 gate57(.Q (g4567), .QB (line57), .D(g33043), .CK(clk));
DFFX1 gate58(.Q (g3057), .QB (line58), .D(g28062), .CK(clk));
DFFX1 gate59(.Q (g3457), .QB (line59), .D(g29263), .CK(clk));
DFFX1 gate60(.Q (g6287), .QB (line60), .D(g30533), .CK(clk));
DFFX1 gate61(.Q (g1500), .QB (line61), .D(g24256), .CK(clk));
DFFX1 gate62(.Q (g2563), .QB (line62), .D(g34015), .CK(clk));
DFFX1 gate63(.Q (g4776), .QB (line63), .D(g34031), .CK(clk));
DFFX1 gate64(.Q (g4593), .QB (line64), .D(g34452), .CK(clk));
DFFX1 gate65(.Q (g6199), .QB (line65), .D(g34646), .CK(clk));
DFFX1 gate66(.Q (g2295), .QB (line66), .D(g34001), .CK(clk));
DFFX1 gate67(.Q (g1384), .QB (line67), .D(g25633), .CK(clk));
DFFX1 gate68(.Q (g1339), .QB (line68), .D(g24259), .CK(clk));
DFFX1 gate69(.Q (g5180), .QB (line69), .D(g33049), .CK(clk));
DFFX1 gate70(.Q (g2844), .QB (line70), .D(g34609), .CK(clk));
DFFX1 gate71(.Q (g1024), .QB (line71), .D(g31869), .CK(clk));
DFFX1 gate72(.Q (g5591), .QB (line72), .D(g30490), .CK(clk));
DFFX1 gate73(.Q (g3598), .QB (line73), .D(g30427), .CK(clk));
DFFX1 gate74(.Q (g4264), .QB (line74), .D(g21894), .CK(clk));
DFFX1 gate75(.Q (g767), .QB (line75), .D(g33965), .CK(clk));
DFFX1 gate76(.Q (g5853), .QB (line76), .D(g34645), .CK(clk));
DFFX1 gate77(.Q (g3321), .QB (line77), .D(g3317), .CK(clk));
DFFX1 gate78(.Q (g2089), .QB (line78), .D(g33571), .CK(clk));
DFFX1 gate79(.Q (g4933), .QB (line79), .D(g34267), .CK(clk));
DFFX1 gate80(.Q (g4521), .QB (line80), .D(g26971), .CK(clk));
DFFX1 gate81(.Q (g5507), .QB (line81), .D(g34644), .CK(clk));
DFFX1 gate82(.Q (g3625), .QB (line82), .D(g3618), .CK(clk));
DFFX1 gate83(.Q (g6291), .QB (line83), .D(g30534), .CK(clk));
DFFX1 gate84(.Q (g294), .QB (line84), .D(g33535), .CK(clk));
DFFX1 gate85(.Q (g5559), .QB (line85), .D(g30498), .CK(clk));
DFFX1 gate86(.Q (g5794), .QB (line86), .D(g25728), .CK(clk));
DFFX1 gate87(.Q (g6144), .QB (line87), .D(g25743), .CK(clk));
DFFX1 gate88(.Q (g3813), .QB (line88), .D(g25684), .CK(clk));
DFFX1 gate89(.Q (g562), .QB (line89), .D(g25613), .CK(clk));
DFFX1 gate90(.Q (g608), .QB (line90), .D(g34438), .CK(clk));
DFFX1 gate91(.Q (g1205), .QB (line91), .D(g24244), .CK(clk));
DFFX1 gate92(.Q (g3909), .QB (line92), .D(g30439), .CK(clk));
DFFX1 gate93(.Q (g6259), .QB (line93), .D(g30541), .CK(clk));
DFFX1 gate94(.Q (g5905), .QB (line94), .D(g30519), .CK(clk));
DFFX1 gate95(.Q (g921), .QB (line95), .D(g25621), .CK(clk));
DFFX1 gate96(.Q (g2955), .QB (line96), .D(g34807), .CK(clk));
DFFX1 gate97(.Q (g203), .QB (line97), .D(g25599), .CK(clk));
DFFX1 gate98(.Q (g6088), .QB (line98), .D(g31924), .CK(clk));
DFFX1 gate99(.Q (g1099), .QB (line99), .D(g24235), .CK(clk));
DFFX1 gate100(.Q (g4878), .QB (line100), .D(g34036), .CK(clk));
DFFX1 gate101(.Q (g5204), .QB (line101), .D(g30476), .CK(clk));
DFFX1 gate102(.Q (g5630), .QB (line102), .D(g5623), .CK(clk));
DFFX1 gate103(.Q (g3606), .QB (line103), .D(g30429), .CK(clk));
DFFX1 gate104(.Q (g1926), .QB (line104), .D(g32997), .CK(clk));
DFFX1 gate105(.Q (g6215), .QB (line105), .D(g33063), .CK(clk));
DFFX1 gate106(.Q (g3586), .QB (line106), .D(g30424), .CK(clk));
DFFX1 gate107(.Q (g291), .QB (line107), .D(g32977), .CK(clk));
DFFX1 gate108(.Q (g4674), .QB (line108), .D(g34026), .CK(clk));
DFFX1 gate109(.Q (g3570), .QB (line109), .D(g30420), .CK(clk));
DFFX1 gate110(.Q (g640), .QB (line110), .D(g637), .CK(clk));
DFFX1 gate111(.Q (g5969), .QB (line111), .D(g6012), .CK(clk));
DFFX1 gate112(.Q (g1862), .QB (line112), .D(g33560), .CK(clk));
DFFX1 gate113(.Q (g676), .QB (line113), .D(g29226), .CK(clk));
DFFX1 gate114(.Q (g843), .QB (line114), .D(g25619), .CK(clk));
DFFX1 gate115(.Q (g4132), .QB (line115), .D(g28076), .CK(clk));
DFFX1 gate116(.Q (g4332), .QB (line116), .D(g34455), .CK(clk));
DFFX1 gate117(.Q (g4153), .QB (line117), .D(g30457), .CK(clk));
DFFX1 gate118(.Q (g5666), .QB (line118), .D(g5637), .CK(clk));
DFFX1 gate119(.Q (g6336), .QB (line119), .D(g33625), .CK(clk));
DFFX1 gate120(.Q (g622), .QB (line120), .D(g34790), .CK(clk));
DFFX1 gate121(.Q (g3506), .QB (line121), .D(g30414), .CK(clk));
DFFX1 gate122(.Q (g4558), .QB (line122), .D(g26966), .CK(clk));
DFFX1 gate123(.Q (g6065), .QB (line123), .D(g31923), .CK(clk));
DFFX1 gate124(.Q (g6322), .QB (line124), .D(g6315), .CK(clk));
DFFX1 gate125(.Q (g3111), .QB (line125), .D(g25656), .CK(clk));
DFFX1 gate126(.Q (g117), .QB (line126), .D(g30390), .CK(clk));
DFFX1 gate127(.Q (g2837), .QB (line127), .D(g26935), .CK(clk));
DFFX1 gate128(.Q (g939), .QB (line128), .D(g34727), .CK(clk));
DFFX1 gate129(.Q (g278), .QB (line129), .D(g25594), .CK(clk));
DFFX1 gate130(.Q (g4492), .QB (line130), .D(g26963), .CK(clk));
DFFX1 gate131(.Q (g4864), .QB (line131), .D(g34034), .CK(clk));
DFFX1 gate132(.Q (g1036), .QB (line132), .D(g33541), .CK(clk));
DFFX1 gate133(.Q (g128), .QB (line133), .D(g28093), .CK(clk));
DFFX1 gate134(.Q (g1178), .QB (line134), .D(g24236), .CK(clk));
DFFX1 gate135(.Q (g3239), .QB (line135), .D(g30404), .CK(clk));
DFFX1 gate136(.Q (g718), .QB (line136), .D(g28051), .CK(clk));
DFFX1 gate137(.Q (g6195), .QB (line137), .D(g29303), .CK(clk));
DFFX1 gate138(.Q (g1135), .QB (line138), .D(g26917), .CK(clk));
DFFX1 gate139(.Q (g6137), .QB (line139), .D(g25741), .CK(clk));
DFFX1 gate140(.Q (g6395), .QB (line140), .D(g33624), .CK(clk));
DFFX1 gate141(.Q (g3380), .QB (line141), .D(g31882), .CK(clk));
DFFX1 gate142(.Q (g5343), .QB (line142), .D(g24337), .CK(clk));
DFFX1 gate143(.Q (g554), .QB (line143), .D(g34911), .CK(clk));
DFFX1 gate144(.Q (g496), .QB (line144), .D(g33963), .CK(clk));
DFFX1 gate145(.Q (g3853), .QB (line145), .D(g34627), .CK(clk));
DFFX1 gate146(.Q (g5134), .QB (line146), .D(g29282), .CK(clk));
DFFX1 gate147(.Q (g1422), .QB (line147), .D(g1418), .CK(clk));
DFFX1 gate148(.Q (g3794), .QB (line148), .D(g25676), .CK(clk));
DFFX1 gate149(.Q (g2485), .QB (line149), .D(g33013), .CK(clk));
DFFX1 gate150(.Q (g925), .QB (line150), .D(g32981), .CK(clk));
DFFX1 gate151(.Q (g48), .QB (line151), .D(g34993), .CK(clk));
DFFX1 gate152(.Q (g5555), .QB (line152), .D(g30483), .CK(clk));
DFFX1 gate153(.Q (g878), .QB (line153), .D(g875), .CK(clk));
DFFX1 gate154(.Q (g1798), .QB (line154), .D(g32994), .CK(clk));
DFFX1 gate155(.Q (g4076), .QB (line155), .D(g28070), .CK(clk));
DFFX1 gate156(.Q (g2941), .QB (line156), .D(g34806), .CK(clk));
DFFX1 gate157(.Q (g3905), .QB (line157), .D(g30453), .CK(clk));
DFFX1 gate158(.Q (g763), .QB (line158), .D(g33539), .CK(clk));
DFFX1 gate159(.Q (g6255), .QB (line159), .D(g30526), .CK(clk));
DFFX1 gate160(.Q (g4375), .QB (line160), .D(g26951), .CK(clk));
DFFX1 gate161(.Q (g4871), .QB (line161), .D(g34035), .CK(clk));
DFFX1 gate162(.Q (g4722), .QB (line162), .D(g34636), .CK(clk));
DFFX1 gate163(.Q (g590), .QB (line163), .D(g32978), .CK(clk));
DFFX1 gate164(.Q (g6692), .QB (line164), .D(g6668), .CK(clk));
DFFX1 gate165(.Q (g1632), .QB (line165), .D(g30348), .CK(clk));
DFFX1 gate166(.Q (g5313), .QB (line166), .D(g24336), .CK(clk));
DFFX1 gate167(.Q (g3100), .QB (line167), .D(g3092), .CK(clk));
DFFX1 gate168(.Q (g1495), .QB (line168), .D(g24250), .CK(clk));
DFFX1 gate169(.Q (g6497), .QB (line169), .D(g6490), .CK(clk));
DFFX1 gate170(.Q (g1437), .QB (line170), .D(g29236), .CK(clk));
DFFX1 gate171(.Q (g6154), .QB (line171), .D(g29298), .CK(clk));
DFFX1 gate172(.Q (g1579), .QB (line172), .D(g1576), .CK(clk));
DFFX1 gate173(.Q (g5567), .QB (line173), .D(g30499), .CK(clk));
DFFX1 gate174(.Q (g1752), .QB (line174), .D(g33976), .CK(clk));
DFFX1 gate175(.Q (g1917), .QB (line175), .D(g32996), .CK(clk));
DFFX1 gate176(.Q (g744), .QB (line176), .D(g30335), .CK(clk));
DFFX1 gate177(.Q (g3040), .QB (line177), .D(g31878), .CK(clk));
DFFX1 gate178(.Q (g4737), .QB (line178), .D(g34637), .CK(clk));
DFFX1 gate179(.Q (g4809), .QB (line179), .D(g25693), .CK(clk));
DFFX1 gate180(.Q (g6267), .QB (line180), .D(g30528), .CK(clk));
DFFX1 gate181(.Q (g3440), .QB (line181), .D(g25661), .CK(clk));
DFFX1 gate182(.Q (g3969), .QB (line182), .D(g4012), .CK(clk));
DFFX1 gate183(.Q (g1442), .QB (line183), .D(g24251), .CK(clk));
DFFX1 gate184(.Q (g5965), .QB (line184), .D(g30521), .CK(clk));
DFFX1 gate185(.Q (g4477), .QB (line185), .D(g26960), .CK(clk));
DFFX1 gate186(.Q (g1233), .QB (line186), .D(g24239), .CK(clk));
DFFX1 gate187(.Q (g4643), .QB (line187), .D(g34259), .CK(clk));
DFFX1 gate188(.Q (g5264), .QB (line188), .D(g30474), .CK(clk));
DFFX1 gate189(.Q (g6329), .QB (line189), .D(g6351), .CK(clk));
DFFX1 gate190(.Q (g2610), .QB (line190), .D(g33016), .CK(clk));
DFFX1 gate191(.Q (g5160), .QB (line191), .D(g34643), .CK(clk));
DFFX1 gate192(.Q (g5360), .QB (line192), .D(g31905), .CK(clk));
DFFX1 gate193(.Q (g5933), .QB (line193), .D(g30510), .CK(clk));
DFFX1 gate194(.Q (g1454), .QB (line194), .D(g29239), .CK(clk));
DFFX1 gate195(.Q (g753), .QB (line195), .D(g26897), .CK(clk));
DFFX1 gate196(.Q (g1296), .QB (line196), .D(g34729), .CK(clk));
DFFX1 gate197(.Q (g3151), .QB (line197), .D(g34625), .CK(clk));
DFFX1 gate198(.Q (g2980), .QB (line198), .D(g34800), .CK(clk));
DFFX1 gate199(.Q (g6727), .QB (line199), .D(g24353), .CK(clk));
DFFX1 gate200(.Q (g3530), .QB (line200), .D(g33029), .CK(clk));
DFFX1 gate201(.Q (g4742), .QB (line201), .D(g21903), .CK(clk));
DFFX1 gate202(.Q (g4104), .QB (line202), .D(g33615), .CK(clk));
DFFX1 gate203(.Q (g1532), .QB (line203), .D(g24253), .CK(clk));
DFFX1 gate204(.Q (g4304), .QB (line204), .D(g24281), .CK(clk));
DFFX1 gate205(.Q (g2177), .QB (line205), .D(g33997), .CK(clk));
DFFX1 gate206(.Q (g3010), .QB (line206), .D(g25651), .CK(clk));
DFFX1 gate207(.Q (g52), .QB (line207), .D(g34997), .CK(clk));
DFFX1 gate208(.Q (g4754), .QB (line208), .D(g34263), .CK(clk));
DFFX1 gate209(.Q (g1189), .QB (line209), .D(g24237), .CK(clk));
DFFX1 gate210(.Q (g2287), .QB (line210), .D(g33584), .CK(clk));
DFFX1 gate211(.Q (g4273), .QB (line211), .D(g24280), .CK(clk));
DFFX1 gate212(.Q (g1389), .QB (line212), .D(g26920), .CK(clk));
DFFX1 gate213(.Q (g1706), .QB (line213), .D(g33548), .CK(clk));
DFFX1 gate214(.Q (g5835), .QB (line214), .D(g29296), .CK(clk));
DFFX1 gate215(.Q (g1171), .QB (line215), .D(g30338), .CK(clk));
DFFX1 gate216(.Q (g4269), .QB (line216), .D(g21895), .CK(clk));
DFFX1 gate217(.Q (g2399), .QB (line217), .D(g33588), .CK(clk));
DFFX1 gate218(.Q (g3372), .QB (line218), .D(g31886), .CK(clk));
DFFX1 gate219(.Q (g4983), .QB (line219), .D(g34041), .CK(clk));
DFFX1 gate220(.Q (g5611), .QB (line220), .D(g30495), .CK(clk));
DFFX1 gate221(.Q (g3618), .QB (line221), .D(g3661), .CK(clk));
DFFX1 gate222(.Q (g4572), .QB (line222), .D(g29279), .CK(clk));
DFFX1 gate223(.Q (g3143), .QB (line223), .D(g25655), .CK(clk));
DFFX1 gate224(.Q (g2898), .QB (line224), .D(g34795), .CK(clk));
DFFX1 gate225(.Q (g3343), .QB (line225), .D(g24269), .CK(clk));
DFFX1 gate226(.Q (g3235), .QB (line226), .D(g30403), .CK(clk));
DFFX1 gate227(.Q (g4543), .QB (line227), .D(g33042), .CK(clk));
DFFX1 gate228(.Q (g3566), .QB (line228), .D(g30419), .CK(clk));
DFFX1 gate229(.Q (g4534), .QB (line229), .D(g34023), .CK(clk));
DFFX1 gate230(.Q (g4961), .QB (line230), .D(g28090), .CK(clk));
DFFX1 gate231(.Q (g6398), .QB (line231), .D(g31926), .CK(clk));
DFFX1 gate232(.Q (g4927), .QB (line232), .D(g34642), .CK(clk));
DFFX1 gate233(.Q (g2259), .QB (line233), .D(g30370), .CK(clk));
DFFX1 gate234(.Q (g2819), .QB (line234), .D(g34448), .CK(clk));
DFFX1 gate235(.Q (g4414), .QB (line235), .D(g26946), .CK(clk));
DFFX1 gate236(.Q (g5802), .QB (line236), .D(g5794), .CK(clk));
DFFX1 gate237(.Q (g2852), .QB (line237), .D(g34610), .CK(clk));
DFFX1 gate238(.Q (g417), .QB (line238), .D(g24209), .CK(clk));
DFFX1 gate239(.Q (g681), .QB (line239), .D(g28047), .CK(clk));
DFFX1 gate240(.Q (g437), .QB (line240), .D(g24206), .CK(clk));
DFFX1 gate241(.Q (g351), .QB (line241), .D(g26891), .CK(clk));
DFFX1 gate242(.Q (g5901), .QB (line242), .D(g30504), .CK(clk));
DFFX1 gate243(.Q (g2886), .QB (line243), .D(g34798), .CK(clk));
DFFX1 gate244(.Q (g3494), .QB (line244), .D(g25669), .CK(clk));
DFFX1 gate245(.Q (g5511), .QB (line245), .D(g30480), .CK(clk));
DFFX1 gate246(.Q (g3518), .QB (line246), .D(g33027), .CK(clk));
DFFX1 gate247(.Q (g1604), .QB (line247), .D(g33972), .CK(clk));
DFFX1 gate248(.Q (g4135), .QB (line248), .D(g28077), .CK(clk));
DFFX1 gate249(.Q (g5092), .QB (line249), .D(g25697), .CK(clk));
DFFX1 gate250(.Q (g4831), .QB (line250), .D(g28099), .CK(clk));
DFFX1 gate251(.Q (g4382), .QB (line251), .D(g26947), .CK(clk));
DFFX1 gate252(.Q (g6386), .QB (line252), .D(g24350), .CK(clk));
DFFX1 gate253(.Q (g479), .QB (line253), .D(g24210), .CK(clk));
DFFX1 gate254(.Q (g3965), .QB (line254), .D(g30455), .CK(clk));
DFFX1 gate255(.Q (g4749), .QB (line255), .D(g28084), .CK(clk));
DFFX1 gate256(.Q (g2008), .QB (line256), .D(g33993), .CK(clk));
DFFX1 gate257(.Q (g736), .QB (line257), .D(g802), .CK(clk));
DFFX1 gate258(.Q (g3933), .QB (line258), .D(g30444), .CK(clk));
DFFX1 gate259(.Q (g222), .QB (line259), .D(g33537), .CK(clk));
DFFX1 gate260(.Q (g3050), .QB (line260), .D(g25650), .CK(clk));
DFFX1 gate261(.Q (g5736), .QB (line261), .D(g31915), .CK(clk));
DFFX1 gate262(.Q (g1052), .QB (line262), .D(g25625), .CK(clk));
DFFX1 gate263(.Q (g58), .QB (line263), .D(g30328), .CK(clk));
DFFX1 gate264(.Q (g5623), .QB (line264), .D(g5666), .CK(clk));
DFFX1 gate265(.Q (g2122), .QB (line265), .D(g30366), .CK(clk));
DFFX1 gate266(.Q (g2465), .QB (line266), .D(g33593), .CK(clk));
DFFX1 gate267(.Q (g6483), .QB (line267), .D(g25755), .CK(clk));
DFFX1 gate268(.Q (g5889), .QB (line268), .D(g30502), .CK(clk));
DFFX1 gate269(.Q (g4495), .QB (line269), .D(g33036), .CK(clk));
DFFX1 gate270(.Q (g365), .QB (line270), .D(g25595), .CK(clk));
DFFX1 gate271(.Q (g4653), .QB (line271), .D(g34462), .CK(clk));
DFFX1 gate272(.Q (g3179), .QB (line272), .D(g33024), .CK(clk));
DFFX1 gate273(.Q (g1728), .QB (line273), .D(g33552), .CK(clk));
DFFX1 gate274(.Q (g2433), .QB (line274), .D(g34014), .CK(clk));
DFFX1 gate275(.Q (g3835), .QB (line275), .D(g29273), .CK(clk));
DFFX1 gate276(.Q (g6187), .QB (line276), .D(g25748), .CK(clk));
DFFX1 gate277(.Q (g4917), .QB (line277), .D(g34638), .CK(clk));
DFFX1 gate278(.Q (g1070), .QB (line278), .D(g30341), .CK(clk));
DFFX1 gate279(.Q (g822), .QB (line279), .D(g26899), .CK(clk));
DFFX1 gate280(.Q (g6027), .QB (line280), .D(g6023), .CK(clk));
DFFX1 gate281(.Q (g914), .QB (line281), .D(g30336), .CK(clk));
DFFX1 gate282(.Q (g5339), .QB (line282), .D(g5335), .CK(clk));
DFFX1 gate283(.Q (g4164), .QB (line283), .D(g26940), .CK(clk));
DFFX1 gate284(.Q (g969), .QB (line284), .D(g25622), .CK(clk));
DFFX1 gate285(.Q (g2807), .QB (line285), .D(g34447), .CK(clk));
DFFX1 gate286(.Q (g5424), .QB (line286), .D(g25709), .CK(clk));
DFFX1 gate287(.Q (g4054), .QB (line287), .D(g33613), .CK(clk));
DFFX1 gate288(.Q (g6191), .QB (line288), .D(g25749), .CK(clk));
DFFX1 gate289(.Q (g5077), .QB (line289), .D(g25704), .CK(clk));
DFFX1 gate290(.Q (g5523), .QB (line290), .D(g33053), .CK(clk));
DFFX1 gate291(.Q (g3680), .QB (line291), .D(g3676), .CK(clk));
DFFX1 gate292(.Q (g6637), .QB (line292), .D(g30555), .CK(clk));
DFFX1 gate293(.Q (g174), .QB (line293), .D(g25601), .CK(clk));
DFFX1 gate294(.Q (g1682), .QB (line294), .D(g33971), .CK(clk));
DFFX1 gate295(.Q (g355), .QB (line295), .D(g26892), .CK(clk));
DFFX1 gate296(.Q (g1087), .QB (line296), .D(g1083), .CK(clk));
DFFX1 gate297(.Q (g1105), .QB (line297), .D(g26915), .CK(clk));
DFFX1 gate298(.Q (g2342), .QB (line298), .D(g33008), .CK(clk));
DFFX1 gate299(.Q (g6307), .QB (line299), .D(g30538), .CK(clk));
DFFX1 gate300(.Q (g3802), .QB (line300), .D(g3794), .CK(clk));
DFFX1 gate301(.Q (g6159), .QB (line301), .D(g25750), .CK(clk));
DFFX1 gate302(.Q (g2255), .QB (line302), .D(g30369), .CK(clk));
DFFX1 gate303(.Q (g2815), .QB (line303), .D(g34446), .CK(clk));
DFFX1 gate304(.Q (g911), .QB (line304), .D(g29230), .CK(clk));
DFFX1 gate305(.Q (g43), .QB (line305), .D(g34789), .CK(clk));
DFFX1 gate306(.Q (g4012), .QB (line306), .D(g3983), .CK(clk));
DFFX1 gate307(.Q (g1748), .QB (line307), .D(g33975), .CK(clk));
DFFX1 gate308(.Q (g5551), .QB (line308), .D(g30497), .CK(clk));
DFFX1 gate309(.Q (g5742), .QB (line309), .D(g31917), .CK(clk));
DFFX1 gate310(.Q (g3558), .QB (line310), .D(g30418), .CK(clk));
DFFX1 gate311(.Q (g5499), .QB (line311), .D(g25721), .CK(clk));
DFFX1 gate312(.Q (g2960), .QB (line312), .D(g34622), .CK(clk));
DFFX1 gate313(.Q (g3901), .QB (line313), .D(g30438), .CK(clk));
DFFX1 gate314(.Q (g4888), .QB (line314), .D(g34266), .CK(clk));
DFFX1 gate315(.Q (g6251), .QB (line315), .D(g30540), .CK(clk));
DFFX1 gate316(.Q (g6315), .QB (line316), .D(g6358), .CK(clk));
DFFX1 gate317(.Q (g1373), .QB (line317), .D(g32986), .CK(clk));
DFFX1 gate318(.Q (g3092), .QB (line318), .D(g25648), .CK(clk));
DFFX1 gate319(.Q (g157), .QB (line319), .D(g33960), .CK(clk));
DFFX1 gate320(.Q (g2783), .QB (line320), .D(g34442), .CK(clk));
DFFX1 gate321(.Q (g4281), .QB (line321), .D(g4277), .CK(clk));
DFFX1 gate322(.Q (g3574), .QB (line322), .D(g30421), .CK(clk));
DFFX1 gate323(.Q (g2112), .QB (line323), .D(g33573), .CK(clk));
DFFX1 gate324(.Q (g1283), .QB (line324), .D(g34730), .CK(clk));
DFFX1 gate325(.Q (g433), .QB (line325), .D(g24205), .CK(clk));
DFFX1 gate326(.Q (g4297), .QB (line326), .D(g4294), .CK(clk));
DFFX1 gate327(.Q (g5983), .QB (line327), .D(g6005), .CK(clk));
DFFX1 gate328(.Q (g1459), .QB (line328), .D(g1399), .CK(clk));
DFFX1 gate329(.Q (g758), .QB (line329), .D(g32979), .CK(clk));
DFFX1 gate330(.Q (g5712), .QB (line330), .D(g25731), .CK(clk));
DFFX1 gate331(.Q (g4138), .QB (line331), .D(g28078), .CK(clk));
DFFX1 gate332(.Q (g4639), .QB (line332), .D(g34025), .CK(clk));
DFFX1 gate333(.Q (g6537), .QB (line333), .D(g25763), .CK(clk));
DFFX1 gate334(.Q (g5543), .QB (line334), .D(g30481), .CK(clk));
DFFX1 gate335(.Q (g1582), .QB (line335), .D(g1500), .CK(clk));
DFFX1 gate336(.Q (g3736), .QB (line336), .D(g31890), .CK(clk));
DFFX1 gate337(.Q (g5961), .QB (line337), .D(g30517), .CK(clk));
DFFX1 gate338(.Q (g6243), .QB (line338), .D(g30539), .CK(clk));
DFFX1 gate339(.Q (g632), .QB (line339), .D(g34880), .CK(clk));
DFFX1 gate340(.Q (g1227), .QB (line340), .D(g24242), .CK(clk));
DFFX1 gate341(.Q (g3889), .QB (line341), .D(g30436), .CK(clk));
DFFX1 gate342(.Q (g3476), .QB (line342), .D(g29265), .CK(clk));
DFFX1 gate343(.Q (g1664), .QB (line343), .D(g32990), .CK(clk));
DFFX1 gate344(.Q (g1246), .QB (line344), .D(g24245), .CK(clk));
DFFX1 gate345(.Q (g6128), .QB (line345), .D(g25739), .CK(clk));
DFFX1 gate346(.Q (g6629), .QB (line346), .D(g30553), .CK(clk));
DFFX1 gate347(.Q (g246), .QB (line347), .D(g26907), .CK(clk));
DFFX1 gate348(.Q (g4049), .QB (line348), .D(g24278), .CK(clk));
DFFX1 gate349(.Q (g4449), .QB (line349), .D(g26955), .CK(clk));
DFFX1 gate350(.Q (g2932), .QB (line350), .D(g24282), .CK(clk));
DFFX1 gate351(.Q (g4575), .QB (line351), .D(g29276), .CK(clk));
DFFX1 gate352(.Q (g4098), .QB (line352), .D(g31894), .CK(clk));
DFFX1 gate353(.Q (g4498), .QB (line353), .D(g33037), .CK(clk));
DFFX1 gate354(.Q (g528), .QB (line354), .D(g26894), .CK(clk));
DFFX1 gate355(.Q (g5436), .QB (line355), .D(g25711), .CK(clk));
DFFX1 gate356(.Q (g16), .QB (line356), .D(g34593), .CK(clk));
DFFX1 gate357(.Q (g3139), .QB (line357), .D(g25654), .CK(clk));
DFFX1 gate358(.Q (g102), .QB (line358), .D(g33962), .CK(clk));
DFFX1 gate359(.Q (g4584), .QB (line359), .D(g34451), .CK(clk));
DFFX1 gate360(.Q (g142), .QB (line360), .D(g34250), .CK(clk));
DFFX1 gate361(.Q (g5335), .QB (line361), .D(g5331), .CK(clk));
DFFX1 gate362(.Q (g5831), .QB (line362), .D(g29295), .CK(clk));
DFFX1 gate363(.Q (g239), .QB (line363), .D(g26905), .CK(clk));
DFFX1 gate364(.Q (g1216), .QB (line364), .D(g25629), .CK(clk));
DFFX1 gate365(.Q (g2848), .QB (line365), .D(g34792), .CK(clk));
DFFX1 gate366(.Q (g5805), .QB (line366), .D(g5798), .CK(clk));
DFFX1 gate367(.Q (g5022), .QB (line367), .D(g25703), .CK(clk));
DFFX1 gate368(.Q (g4019), .QB (line368), .D(g4000), .CK(clk));
DFFX1 gate369(.Q (g1030), .QB (line369), .D(g32983), .CK(clk));
DFFX1 gate370(.Q (g3672), .QB (line370), .D(g3668), .CK(clk));
DFFX1 gate371(.Q (g3231), .QB (line371), .D(g30402), .CK(clk));
DFFX1 gate372(.Q (g6490), .QB (line372), .D(g25757), .CK(clk));
DFFX1 gate373(.Q (g1430), .QB (line373), .D(g1426), .CK(clk));
DFFX1 gate374(.Q (g4452), .QB (line374), .D(g4446), .CK(clk));
DFFX1 gate375(.Q (g2241), .QB (line375), .D(g33999), .CK(clk));
DFFX1 gate376(.Q (g1564), .QB (line376), .D(g24262), .CK(clk));
DFFX1 gate377(.Q (g5798), .QB (line377), .D(g25729), .CK(clk));
DFFX1 gate378(.Q (g6148), .QB (line378), .D(g6140), .CK(clk));
DFFX1 gate379(.Q (g6649), .QB (line379), .D(g30558), .CK(clk));
DFFX1 gate380(.Q (g110), .QB (line380), .D(g34848), .CK(clk));
DFFX1 gate381(.Q (g884), .QB (line381), .D(g881), .CK(clk));
DFFX1 gate382(.Q (g3742), .QB (line382), .D(g31892), .CK(clk));
DFFX1 gate383(.Q (g225), .QB (line383), .D(g26901), .CK(clk));
DFFX1 gate384(.Q (g4486), .QB (line384), .D(g26961), .CK(clk));
DFFX1 gate385(.Q (g4504), .QB (line385), .D(g33039), .CK(clk));
DFFX1 gate386(.Q (g5873), .QB (line386), .D(g33059), .CK(clk));
DFFX1 gate387(.Q (g5037), .QB (line387), .D(g31899), .CK(clk));
DFFX1 gate388(.Q (g2319), .QB (line388), .D(g33007), .CK(clk));
DFFX1 gate389(.Q (g5495), .QB (line389), .D(g25720), .CK(clk));
DFFX1 gate390(.Q (g4185), .QB (line390), .D(g21891), .CK(clk));
DFFX1 gate391(.Q (g5208), .QB (line391), .D(g30462), .CK(clk));
DFFX1 gate392(.Q (g2152), .QB (line392), .D(g18422), .CK(clk));
DFFX1 gate393(.Q (g5579), .QB (line393), .D(g30487), .CK(clk));
DFFX1 gate394(.Q (g5869), .QB (line394), .D(g33058), .CK(clk));
DFFX1 gate395(.Q (g5719), .QB (line395), .D(g31916), .CK(clk));
DFFX1 gate396(.Q (g1589), .QB (line396), .D(g24261), .CK(clk));
DFFX1 gate397(.Q (g5752), .QB (line397), .D(g25730), .CK(clk));
DFFX1 gate398(.Q (g6279), .QB (line398), .D(g30531), .CK(clk));
DFFX1 gate399(.Q (g5917), .QB (line399), .D(g30506), .CK(clk));
DFFX1 gate400(.Q (g2975), .QB (line400), .D(g34804), .CK(clk));
DFFX1 gate401(.Q (g6167), .QB (line401), .D(g25747), .CK(clk));
DFFX1 gate402(.Q (g3983), .QB (line402), .D(g4005), .CK(clk));
DFFX1 gate403(.Q (g2599), .QB (line403), .D(g33601), .CK(clk));
DFFX1 gate404(.Q (g1448), .QB (line404), .D(g26922), .CK(clk));
DFFX1 gate405(.Q (g881), .QB (line405), .D(g878), .CK(clk));
DFFX1 gate406(.Q (g3712), .QB (line406), .D(g25679), .CK(clk));
DFFX1 gate407(.Q (g2370), .QB (line407), .D(g29250), .CK(clk));
DFFX1 gate408(.Q (g5164), .QB (line408), .D(g30459), .CK(clk));
DFFX1 gate409(.Q (g1333), .QB (line409), .D(g1582), .CK(clk));
DFFX1 gate410(.Q (g153), .QB (line410), .D(g33534), .CK(clk));
DFFX1 gate411(.Q (g6549), .QB (line411), .D(g30543), .CK(clk));
DFFX1 gate412(.Q (g4087), .QB (line412), .D(g29275), .CK(clk));
DFFX1 gate413(.Q (g4801), .QB (line413), .D(g34030), .CK(clk));
DFFX1 gate414(.Q (g2984), .QB (line414), .D(g34980), .CK(clk));
DFFX1 gate415(.Q (g3961), .QB (line415), .D(g30451), .CK(clk));
DFFX1 gate416(.Q (g5770), .QB (line416), .D(g25723), .CK(clk));
DFFX1 gate417(.Q (g962), .QB (line417), .D(g25627), .CK(clk));
DFFX1 gate418(.Q (g101), .QB (line418), .D(g34787), .CK(clk));
DFFX1 gate419(.Q (g4226), .QB (line419), .D(g4222), .CK(clk));
DFFX1 gate420(.Q (g6625), .QB (line420), .D(g30552), .CK(clk));
DFFX1 gate421(.Q (g51), .QB (line421), .D(g34996), .CK(clk));
DFFX1 gate422(.Q (g1018), .QB (line422), .D(g30337), .CK(clk));
DFFX1 gate423(.Q (g1418), .QB (line423), .D(g24254), .CK(clk));
DFFX1 gate424(.Q (g4045), .QB (line424), .D(g24277), .CK(clk));
DFFX1 gate425(.Q (g1467), .QB (line425), .D(g29237), .CK(clk));
DFFX1 gate426(.Q (g2461), .QB (line426), .D(g30378), .CK(clk));
DFFX1 gate427(.Q (g5706), .QB (line427), .D(g31912), .CK(clk));
DFFX1 gate428(.Q (g457), .QB (line428), .D(g25603), .CK(clk));
DFFX1 gate429(.Q (g2756), .QB (line429), .D(g33019), .CK(clk));
DFFX1 gate430(.Q (g5990), .QB (line430), .D(g33623), .CK(clk));
DFFX1 gate431(.Q (g471), .QB (line431), .D(g25608), .CK(clk));
DFFX1 gate432(.Q (g1256), .QB (line432), .D(g29235), .CK(clk));
DFFX1 gate433(.Q (g5029), .QB (line433), .D(g31902), .CK(clk));
DFFX1 gate434(.Q (g6519), .QB (line434), .D(g29306), .CK(clk));
DFFX1 gate435(.Q (g4169), .QB (line435), .D(g28080), .CK(clk));
DFFX1 gate436(.Q (g1816), .QB (line436), .D(g33978), .CK(clk));
DFFX1 gate437(.Q (g4369), .QB (line437), .D(g26970), .CK(clk));
DFFX1 gate438(.Q (g3436), .QB (line438), .D(g25660), .CK(clk));
DFFX1 gate439(.Q (g5787), .QB (line439), .D(g25726), .CK(clk));
DFFX1 gate440(.Q (g4578), .QB (line440), .D(g29278), .CK(clk));
DFFX1 gate441(.Q (g4459), .QB (line441), .D(g34253), .CK(clk));
DFFX1 gate442(.Q (g3831), .QB (line442), .D(g29272), .CK(clk));
DFFX1 gate443(.Q (g2514), .QB (line443), .D(g33595), .CK(clk));
DFFX1 gate444(.Q (g3288), .QB (line444), .D(g33610), .CK(clk));
DFFX1 gate445(.Q (g2403), .QB (line445), .D(g33589), .CK(clk));
DFFX1 gate446(.Q (g2145), .QB (line446), .D(g34605), .CK(clk));
DFFX1 gate447(.Q (g1700), .QB (line447), .D(g30350), .CK(clk));
DFFX1 gate448(.Q (g513), .QB (line448), .D(g25611), .CK(clk));
DFFX1 gate449(.Q (g2841), .QB (line449), .D(g26936), .CK(clk));
DFFX1 gate450(.Q (g5297), .QB (line450), .D(g33619), .CK(clk));
DFFX1 gate451(.Q (g3805), .QB (line451), .D(g3798), .CK(clk));
DFFX1 gate452(.Q (g2763), .QB (line452), .D(g34022), .CK(clk));
DFFX1 gate453(.Q (g4793), .QB (line453), .D(g34033), .CK(clk));
DFFX1 gate454(.Q (g952), .QB (line454), .D(g34726), .CK(clk));
DFFX1 gate455(.Q (g1263), .QB (line455), .D(g31870), .CK(clk));
DFFX1 gate456(.Q (g1950), .QB (line456), .D(g33985), .CK(clk));
DFFX1 gate457(.Q (g5138), .QB (line457), .D(g29283), .CK(clk));
DFFX1 gate458(.Q (g2307), .QB (line458), .D(g34003), .CK(clk));
DFFX1 gate459(.Q (g5109), .QB (line459), .D(g5101), .CK(clk));
DFFX1 gate460(.Q (g5791), .QB (line460), .D(g25727), .CK(clk));
DFFX1 gate461(.Q (g3798), .QB (line461), .D(g25677), .CK(clk));
DFFX1 gate462(.Q (g4664), .QB (line462), .D(g34463), .CK(clk));
DFFX1 gate463(.Q (g2223), .QB (line463), .D(g33006), .CK(clk));
DFFX1 gate464(.Q (g5808), .QB (line464), .D(g29292), .CK(clk));
DFFX1 gate465(.Q (g6645), .QB (line465), .D(g30557), .CK(clk));
DFFX1 gate466(.Q (g2016), .QB (line466), .D(g33989), .CK(clk));
DFFX1 gate467(.Q (g5759), .QB (line467), .D(g28098), .CK(clk));
DFFX1 gate468(.Q (g3873), .QB (line468), .D(g33033), .CK(clk));
DFFX1 gate469(.Q (g3632), .QB (line469), .D(g3654), .CK(clk));
DFFX1 gate470(.Q (g2315), .QB (line470), .D(g34005), .CK(clk));
DFFX1 gate471(.Q (g2811), .QB (line471), .D(g26932), .CK(clk));
DFFX1 gate472(.Q (g5957), .QB (line472), .D(g30516), .CK(clk));
DFFX1 gate473(.Q (g2047), .QB (line473), .D(g33575), .CK(clk));
DFFX1 gate474(.Q (g3869), .QB (line474), .D(g33032), .CK(clk));
DFFX1 gate475(.Q (g6358), .QB (line475), .D(g6329), .CK(clk));
DFFX1 gate476(.Q (g3719), .QB (line476), .D(g31891), .CK(clk));
DFFX1 gate477(.Q (g5575), .QB (line477), .D(g30486), .CK(clk));
DFFX1 gate478(.Q (g46), .QB (line478), .D(g34991), .CK(clk));
DFFX1 gate479(.Q (g3752), .QB (line479), .D(g25678), .CK(clk));
DFFX1 gate480(.Q (g3917), .QB (line480), .D(g30440), .CK(clk));
DFFX1 gate481(.Q (g4188), .QB (line481), .D(g4191), .CK(clk));
DFFX1 gate482(.Q (g1585), .QB (line482), .D(g1570), .CK(clk));
DFFX1 gate483(.Q (g4388), .QB (line483), .D(g26949), .CK(clk));
DFFX1 gate484(.Q (g6275), .QB (line484), .D(g30530), .CK(clk));
DFFX1 gate485(.Q (g6311), .QB (line485), .D(g30542), .CK(clk));
DFFX1 gate486(.Q (g4216), .QB (line486), .D(g4213), .CK(clk));
DFFX1 gate487(.Q (g1041), .QB (line487), .D(g25624), .CK(clk));
DFFX1 gate488(.Q (g2595), .QB (line488), .D(g30383), .CK(clk));
DFFX1 gate489(.Q (g2537), .QB (line489), .D(g33597), .CK(clk));
DFFX1 gate490(.Q (g136), .QB (line490), .D(g34598), .CK(clk));
DFFX1 gate491(.Q (g4430), .QB (line491), .D(g26957), .CK(clk));
DFFX1 gate492(.Q (g4564), .QB (line492), .D(g26967), .CK(clk));
DFFX1 gate493(.Q (g3454), .QB (line493), .D(g3447), .CK(clk));
DFFX1 gate494(.Q (g4826), .QB (line494), .D(g28102), .CK(clk));
DFFX1 gate495(.Q (g6239), .QB (line495), .D(g30524), .CK(clk));
DFFX1 gate496(.Q (g3770), .QB (line496), .D(g25671), .CK(clk));
DFFX1 gate497(.Q (g232), .QB (line497), .D(g26903), .CK(clk));
DFFX1 gate498(.Q (g5268), .QB (line498), .D(g30475), .CK(clk));
DFFX1 gate499(.Q (g6545), .QB (line499), .D(g34647), .CK(clk));
DFFX1 gate500(.Q (g2417), .QB (line500), .D(g30377), .CK(clk));
DFFX1 gate501(.Q (g1772), .QB (line501), .D(g33553), .CK(clk));
DFFX1 gate502(.Q (g4741), .QB (line502), .D(g21902), .CK(clk));
DFFX1 gate503(.Q (g5052), .QB (line503), .D(g31903), .CK(clk));
DFFX1 gate504(.Q (g5452), .QB (line504), .D(g25715), .CK(clk));
DFFX1 gate505(.Q (g1890), .QB (line505), .D(g33984), .CK(clk));
DFFX1 gate506(.Q (g2629), .QB (line506), .D(g33602), .CK(clk));
DFFX1 gate507(.Q (g572), .QB (line507), .D(g28045), .CK(clk));
DFFX1 gate508(.Q (g2130), .QB (line508), .D(g34603), .CK(clk));
DFFX1 gate509(.Q (g4108), .QB (line509), .D(g33035), .CK(clk));
DFFX1 gate510(.Q (g4308), .QB (line510), .D(g4304), .CK(clk));
DFFX1 gate511(.Q (g475), .QB (line511), .D(g24208), .CK(clk));
DFFX1 gate512(.Q (g990), .QB (line512), .D(g1239), .CK(clk));
DFFX1 gate513(.Q (g31), .QB (line513), .D(g34596), .CK(clk));
DFFX1 gate514(.Q (g3412), .QB (line514), .D(g28064), .CK(clk));
DFFX1 gate515(.Q (g45), .QB (line515), .D(g34990), .CK(clk));
DFFX1 gate516(.Q (g799), .QB (line516), .D(g24213), .CK(clk));
DFFX1 gate517(.Q (g3706), .QB (line517), .D(g31887), .CK(clk));
DFFX1 gate518(.Q (g3990), .QB (line518), .D(g33614), .CK(clk));
DFFX1 gate519(.Q (g5385), .QB (line519), .D(g31907), .CK(clk));
DFFX1 gate520(.Q (g5881), .QB (line520), .D(g33060), .CK(clk));
DFFX1 gate521(.Q (g1992), .QB (line521), .D(g30362), .CK(clk));
DFFX1 gate522(.Q (g3029), .QB (line522), .D(g31875), .CK(clk));
DFFX1 gate523(.Q (g3171), .QB (line523), .D(g33023), .CK(clk));
DFFX1 gate524(.Q (g3787), .QB (line524), .D(g25674), .CK(clk));
DFFX1 gate525(.Q (g812), .QB (line525), .D(g26898), .CK(clk));
DFFX1 gate526(.Q (g832), .QB (line526), .D(g25618), .CK(clk));
DFFX1 gate527(.Q (g5897), .QB (line527), .D(g30518), .CK(clk));
DFFX1 gate528(.Q (g4165), .QB (line528), .D(g28079), .CK(clk));
DFFX1 gate529(.Q (g4571), .QB (line529), .D(g6974), .CK(clk));
DFFX1 gate530(.Q (g3281), .QB (line530), .D(g3303), .CK(clk));
DFFX1 gate531(.Q (g4455), .QB (line531), .D(g26959), .CK(clk));
DFFX1 gate532(.Q (g2902), .QB (line532), .D(g34801), .CK(clk));
DFFX1 gate533(.Q (g333), .QB (line533), .D(g26884), .CK(clk));
DFFX1 gate534(.Q (g168), .QB (line534), .D(g25600), .CK(clk));
DFFX1 gate535(.Q (g2823), .QB (line535), .D(g26933), .CK(clk));
DFFX1 gate536(.Q (g3684), .QB (line536), .D(g28066), .CK(clk));
DFFX1 gate537(.Q (g3639), .QB (line537), .D(g33612), .CK(clk));
DFFX1 gate538(.Q (g5331), .QB (line538), .D(g5327), .CK(clk));
DFFX1 gate539(.Q (g3338), .QB (line539), .D(g24268), .CK(clk));
DFFX1 gate540(.Q (g5406), .QB (line540), .D(g25716), .CK(clk));
DFFX1 gate541(.Q (g3791), .QB (line541), .D(g25675), .CK(clk));
DFFX1 gate542(.Q (g269), .QB (line542), .D(g26906), .CK(clk));
DFFX1 gate543(.Q (g401), .QB (line543), .D(g24203), .CK(clk));
DFFX1 gate544(.Q (g6040), .QB (line544), .D(g24346), .CK(clk));
DFFX1 gate545(.Q (g441), .QB (line545), .D(g24207), .CK(clk));
DFFX1 gate546(.Q (g5105), .QB (line546), .D(g25701), .CK(clk));
DFFX1 gate547(.Q (g3808), .QB (line547), .D(g29269), .CK(clk));
DFFX1 gate548(.Q (g9), .QB (line548), .D(g34592), .CK(clk));
DFFX1 gate549(.Q (g3759), .QB (line549), .D(g28068), .CK(clk));
DFFX1 gate550(.Q (g4467), .QB (line550), .D(g34255), .CK(clk));
DFFX1 gate551(.Q (g3957), .QB (line551), .D(g30450), .CK(clk));
DFFX1 gate552(.Q (g4093), .QB (line552), .D(g30456), .CK(clk));
DFFX1 gate553(.Q (g1760), .QB (line553), .D(g32991), .CK(clk));
DFFX1 gate554(.Q (g6151), .QB (line554), .D(g6144), .CK(clk));
DFFX1 gate555(.Q (g6351), .QB (line555), .D(g24348), .CK(clk));
DFFX1 gate556(.Q (g160), .QB (line556), .D(g34249), .CK(clk));
DFFX1 gate557(.Q (g5445), .QB (line557), .D(g25713), .CK(clk));
DFFX1 gate558(.Q (g5373), .QB (line558), .D(g31909), .CK(clk));
DFFX1 gate559(.Q (g2279), .QB (line559), .D(g30371), .CK(clk));
DFFX1 gate560(.Q (g3498), .QB (line560), .D(g29268), .CK(clk));
DFFX1 gate561(.Q (g586), .QB (line561), .D(g29224), .CK(clk));
DFFX1 gate562(.Q (g869), .QB (line562), .D(g859), .CK(clk));
DFFX1 gate563(.Q (g2619), .QB (line563), .D(g33017), .CK(clk));
DFFX1 gate564(.Q (g1183), .QB (line564), .D(g30339), .CK(clk));
DFFX1 gate565(.Q (g1608), .QB (line565), .D(g33967), .CK(clk));
DFFX1 gate566(.Q (g4197), .QB (line566), .D(g4194), .CK(clk));
DFFX1 gate567(.Q (g5283), .QB (line567), .D(g5276), .CK(clk));
DFFX1 gate568(.Q (g1779), .QB (line568), .D(g33559), .CK(clk));
DFFX1 gate569(.Q (g2652), .QB (line569), .D(g29255), .CK(clk));
DFFX1 gate570(.Q (g5459), .QB (line570), .D(g5452), .CK(clk));
DFFX1 gate571(.Q (g2193), .QB (line571), .D(g30368), .CK(clk));
DFFX1 gate572(.Q (g2393), .QB (line572), .D(g30375), .CK(clk));
DFFX1 gate573(.Q (g5767), .QB (line573), .D(g25732), .CK(clk));
DFFX1 gate574(.Q (g661), .QB (line574), .D(g28052), .CK(clk));
DFFX1 gate575(.Q (g4950), .QB (line575), .D(g28089), .CK(clk));
DFFX1 gate576(.Q (g5535), .QB (line576), .D(g33055), .CK(clk));
DFFX1 gate577(.Q (g2834), .QB (line577), .D(g30392), .CK(clk));
DFFX1 gate578(.Q (g1361), .QB (line578), .D(g30343), .CK(clk));
DFFX1 gate579(.Q (g3419), .QB (line579), .D(g25657), .CK(clk));
DFFX1 gate580(.Q (g6235), .QB (line580), .D(g30523), .CK(clk));
DFFX1 gate581(.Q (g1146), .QB (line581), .D(g24233), .CK(clk));
DFFX1 gate582(.Q (g2625), .QB (line582), .D(g33018), .CK(clk));
DFFX1 gate583(.Q (g150), .QB (line583), .D(g32976), .CK(clk));
DFFX1 gate584(.Q (g1696), .QB (line584), .D(g30349), .CK(clk));
DFFX1 gate585(.Q (g6555), .QB (line585), .D(g33067), .CK(clk));
DFFX1 gate586(.Q (g859), .QB (line586), .D(g26900), .CK(clk));
DFFX1 gate587(.Q (g3385), .QB (line587), .D(g31883), .CK(clk));
DFFX1 gate588(.Q (g3881), .QB (line588), .D(g33034), .CK(clk));
DFFX1 gate589(.Q (g6621), .QB (line589), .D(g30551), .CK(clk));
DFFX1 gate590(.Q (g3470), .QB (line590), .D(g25667), .CK(clk));
DFFX1 gate591(.Q (g3897), .QB (line591), .D(g30452), .CK(clk));
DFFX1 gate592(.Q (g518), .QB (line592), .D(g25612), .CK(clk));
DFFX1 gate593(.Q (g3025), .QB (line593), .D(g31874), .CK(clk));
DFFX1 gate594(.Q (g538), .QB (line594), .D(g34719), .CK(clk));
DFFX1 gate595(.Q (g2606), .QB (line595), .D(g33607), .CK(clk));
DFFX1 gate596(.Q (g1472), .QB (line596), .D(g26923), .CK(clk));
DFFX1 gate597(.Q (g6113), .QB (line597), .D(g25746), .CK(clk));
DFFX1 gate598(.Q (g542), .QB (line598), .D(g24211), .CK(clk));
DFFX1 gate599(.Q (g5188), .QB (line599), .D(g33050), .CK(clk));
DFFX1 gate600(.Q (g5689), .QB (line600), .D(g24341), .CK(clk));
DFFX1 gate601(.Q (g1116), .QB (line601), .D(g1056), .CK(clk));
DFFX1 gate602(.Q (g405), .QB (line602), .D(g24201), .CK(clk));
DFFX1 gate603(.Q (g5216), .QB (line603), .D(g30463), .CK(clk));
DFFX1 gate604(.Q (g6494), .QB (line604), .D(g6486), .CK(clk));
DFFX1 gate605(.Q (g4669), .QB (line605), .D(g34464), .CK(clk));
DFFX1 gate606(.Q (g5428), .QB (line606), .D(g25710), .CK(clk));
DFFX1 gate607(.Q (g996), .QB (line607), .D(g24243), .CK(clk));
DFFX1 gate608(.Q (g4531), .QB (line608), .D(g24335), .CK(clk));
DFFX1 gate609(.Q (g2860), .QB (line609), .D(g34611), .CK(clk));
DFFX1 gate610(.Q (g4743), .QB (line610), .D(g34262), .CK(clk));
DFFX1 gate611(.Q (g6593), .QB (line611), .D(g30546), .CK(clk));
DFFX1 gate612(.Q (g2710), .QB (line612), .D(g18527), .CK(clk));
DFFX1 gate613(.Q (g215), .QB (line613), .D(g25591), .CK(clk));
DFFX1 gate614(.Q (g4411), .QB (line614), .D(g4414), .CK(clk));
DFFX1 gate615(.Q (g1413), .QB (line615), .D(g30347), .CK(clk));
DFFX1 gate616(.Q (g4474), .QB (line616), .D(g10384), .CK(clk));
DFFX1 gate617(.Q (g5308), .QB (line617), .D(g5283), .CK(clk));
DFFX1 gate618(.Q (g6641), .QB (line618), .D(g30556), .CK(clk));
DFFX1 gate619(.Q (g3045), .QB (line619), .D(g33020), .CK(clk));
DFFX1 gate620(.Q (g6), .QB (line620), .D(g34589), .CK(clk));
DFFX1 gate621(.Q (g1936), .QB (line621), .D(g33562), .CK(clk));
DFFX1 gate622(.Q (g55), .QB (line622), .D(g35002), .CK(clk));
DFFX1 gate623(.Q (g504), .QB (line623), .D(g25610), .CK(clk));
DFFX1 gate624(.Q (g2587), .QB (line624), .D(g33015), .CK(clk));
DFFX1 gate625(.Q (g4480), .QB (line625), .D(g31896), .CK(clk));
DFFX1 gate626(.Q (g2311), .QB (line626), .D(g34004), .CK(clk));
DFFX1 gate627(.Q (g3602), .QB (line627), .D(g30428), .CK(clk));
DFFX1 gate628(.Q (g5571), .QB (line628), .D(g30485), .CK(clk));
DFFX1 gate629(.Q (g3578), .QB (line629), .D(g30422), .CK(clk));
DFFX1 gate630(.Q (g468), .QB (line630), .D(g25606), .CK(clk));
DFFX1 gate631(.Q (g5448), .QB (line631), .D(g25714), .CK(clk));
DFFX1 gate632(.Q (g3767), .QB (line632), .D(g25680), .CK(clk));
DFFX1 gate633(.Q (g5827), .QB (line633), .D(g29294), .CK(clk));
DFFX1 gate634(.Q (g3582), .QB (line634), .D(g30423), .CK(clk));
DFFX1 gate635(.Q (g6271), .QB (line635), .D(g30529), .CK(clk));
DFFX1 gate636(.Q (g4688), .QB (line636), .D(g34028), .CK(clk));
DFFX1 gate637(.Q (g5774), .QB (line637), .D(g25724), .CK(clk));
DFFX1 gate638(.Q (g2380), .QB (line638), .D(g33587), .CK(clk));
DFFX1 gate639(.Q (g5196), .QB (line639), .D(g30460), .CK(clk));
DFFX1 gate640(.Q (g5396), .QB (line640), .D(g31910), .CK(clk));
DFFX1 gate641(.Q (g3227), .QB (line641), .D(g30401), .CK(clk));
DFFX1 gate642(.Q (g2020), .QB (line642), .D(g33990), .CK(clk));
DFFX1 gate643(.Q (g4000), .QB (line643), .D(g3976), .CK(clk));
DFFX1 gate644(.Q (g1079), .QB (line644), .D(g1075), .CK(clk));
DFFX1 gate645(.Q (g6541), .QB (line645), .D(g29309), .CK(clk));
DFFX1 gate646(.Q (g3203), .QB (line646), .D(g30411), .CK(clk));
DFFX1 gate647(.Q (g1668), .QB (line647), .D(g33546), .CK(clk));
DFFX1 gate648(.Q (g4760), .QB (line648), .D(g28085), .CK(clk));
DFFX1 gate649(.Q (g262), .QB (line649), .D(g26904), .CK(clk));
DFFX1 gate650(.Q (g1840), .QB (line650), .D(g33556), .CK(clk));
DFFX1 gate651(.Q (g70), .QB (line651), .D(g18093), .CK(clk));
DFFX1 gate652(.Q (g5467), .QB (line652), .D(g25722), .CK(clk));
DFFX1 gate653(.Q (g460), .QB (line653), .D(g25605), .CK(clk));
DFFX1 gate654(.Q (g6209), .QB (line654), .D(g33062), .CK(clk));
DFFX1 gate655(.Q (g74), .QB (line655), .D(g26893), .CK(clk));
DFFX1 gate656(.Q (g5290), .QB (line656), .D(g5313), .CK(clk));
DFFX1 gate657(.Q (g655), .QB (line657), .D(g28050), .CK(clk));
DFFX1 gate658(.Q (g3502), .QB (line658), .D(g34626), .CK(clk));
DFFX1 gate659(.Q (g2204), .QB (line659), .D(g33583), .CK(clk));
DFFX1 gate660(.Q (g5256), .QB (line660), .D(g30472), .CK(clk));
DFFX1 gate661(.Q (g4608), .QB (line661), .D(g34454), .CK(clk));
DFFX1 gate662(.Q (g794), .QB (line662), .D(g34850), .CK(clk));
DFFX1 gate663(.Q (g4023), .QB (line663), .D(g4019), .CK(clk));
DFFX1 gate664(.Q (g4423), .QB (line664), .D(g4537), .CK(clk));
DFFX1 gate665(.Q (g3689), .QB (line665), .D(g24272), .CK(clk));
DFFX1 gate666(.Q (g5381), .QB (line666), .D(g31906), .CK(clk));
DFFX1 gate667(.Q (g5685), .QB (line667), .D(g5681), .CK(clk));
DFFX1 gate668(.Q (g703), .QB (line668), .D(g24214), .CK(clk));
DFFX1 gate669(.Q (g5421), .QB (line669), .D(g25718), .CK(clk));
DFFX1 gate670(.Q (g862), .QB (line670), .D(g26909), .CK(clk));
DFFX1 gate671(.Q (g3247), .QB (line671), .D(g30406), .CK(clk));
DFFX1 gate672(.Q (g2040), .QB (line672), .D(g33569), .CK(clk));
DFFX1 gate673(.Q (g4999), .QB (line673), .D(g25694), .CK(clk));
DFFX1 gate674(.Q (g4146), .QB (line674), .D(g34628), .CK(clk));
DFFX1 gate675(.Q (g4633), .QB (line675), .D(g34458), .CK(clk));
DFFX1 gate676(.Q (g1157), .QB (line676), .D(g24240), .CK(clk));
DFFX1 gate677(.Q (g5723), .QB (line677), .D(g31918), .CK(clk));
DFFX1 gate678(.Q (g4732), .QB (line678), .D(g34634), .CK(clk));
DFFX1 gate679(.Q (g5101), .QB (line679), .D(g25700), .CK(clk));
DFFX1 gate680(.Q (g5817), .QB (line680), .D(g29293), .CK(clk));
DFFX1 gate681(.Q (g2151), .QB (line681), .D(g18421), .CK(clk));
DFFX1 gate682(.Q (g2351), .QB (line682), .D(g33009), .CK(clk));
DFFX1 gate683(.Q (g2648), .QB (line683), .D(g33603), .CK(clk));
DFFX1 gate684(.Q (g6736), .QB (line684), .D(g24355), .CK(clk));
DFFX1 gate685(.Q (g4944), .QB (line685), .D(g34268), .CK(clk));
DFFX1 gate686(.Q (g4072), .QB (line686), .D(g25691), .CK(clk));
DFFX1 gate687(.Q (g344), .QB (line687), .D(g26890), .CK(clk));
DFFX1 gate688(.Q (g4443), .QB (line688), .D(g4449), .CK(clk));
DFFX1 gate689(.Q (g3466), .QB (line689), .D(g29264), .CK(clk));
DFFX1 gate690(.Q (g4116), .QB (line690), .D(g28072), .CK(clk));
DFFX1 gate691(.Q (g5041), .QB (line691), .D(g31900), .CK(clk));
DFFX1 gate692(.Q (g5441), .QB (line692), .D(g25712), .CK(clk));
DFFX1 gate693(.Q (g4434), .QB (line693), .D(g26956), .CK(clk));
DFFX1 gate694(.Q (g3827), .QB (line694), .D(g29271), .CK(clk));
DFFX1 gate695(.Q (g6500), .QB (line695), .D(g29304), .CK(clk));
DFFX1 gate696(.Q (g5673), .QB (line696), .D(g5654), .CK(clk));
DFFX1 gate697(.Q (g3133), .QB (line697), .D(g29261), .CK(clk));
DFFX1 gate698(.Q (g3333), .QB (line698), .D(g28063), .CK(clk));
DFFX1 gate699(.Q (g979), .QB (line699), .D(g1116), .CK(clk));
DFFX1 gate700(.Q (g4681), .QB (line700), .D(g34027), .CK(clk));
DFFX1 gate701(.Q (g298), .QB (line701), .D(g33961), .CK(clk));
DFFX1 gate702(.Q (g3774), .QB (line702), .D(g25672), .CK(clk));
DFFX1 gate703(.Q (g2667), .QB (line703), .D(g33604), .CK(clk));
DFFX1 gate704(.Q (g3396), .QB (line704), .D(g33025), .CK(clk));
DFFX1 gate705(.Q (g4210), .QB (line705), .D(g4207), .CK(clk));
DFFX1 gate706(.Q (g1894), .QB (line706), .D(g32995), .CK(clk));
DFFX1 gate707(.Q (g2988), .QB (line707), .D(g34624), .CK(clk));
DFFX1 gate708(.Q (g3538), .QB (line708), .D(g30415), .CK(clk));
DFFX1 gate709(.Q (g301), .QB (line709), .D(g33536), .CK(clk));
DFFX1 gate710(.Q (g341), .QB (line710), .D(g26888), .CK(clk));
DFFX1 gate711(.Q (g827), .QB (line711), .D(g28055), .CK(clk));
DFFX1 gate712(.Q (g1075), .QB (line712), .D(g24238), .CK(clk));
DFFX1 gate713(.Q (g6077), .QB (line713), .D(g31921), .CK(clk));
DFFX1 gate714(.Q (g2555), .QB (line714), .D(g33600), .CK(clk));
DFFX1 gate715(.Q (g5011), .QB (line715), .D(g28105), .CK(clk));
DFFX1 gate716(.Q (g199), .QB (line716), .D(g34721), .CK(clk));
DFFX1 gate717(.Q (g6523), .QB (line717), .D(g29307), .CK(clk));
DFFX1 gate718(.Q (g1526), .QB (line718), .D(g30345), .CK(clk));
DFFX1 gate719(.Q (g4601), .QB (line719), .D(g34453), .CK(clk));
DFFX1 gate720(.Q (g854), .QB (line720), .D(g32980), .CK(clk));
DFFX1 gate721(.Q (g1484), .QB (line721), .D(g29238), .CK(clk));
DFFX1 gate722(.Q (g4922), .QB (line722), .D(g34639), .CK(clk));
DFFX1 gate723(.Q (g5080), .QB (line723), .D(g25695), .CK(clk));
DFFX1 gate724(.Q (g5863), .QB (line724), .D(g33057), .CK(clk));
DFFX1 gate725(.Q (g4581), .QB (line725), .D(g26969), .CK(clk));
DFFX1 gate726(.Q (g3021), .QB (line726), .D(g31879), .CK(clk));
DFFX1 gate727(.Q (g2518), .QB (line727), .D(g29253), .CK(clk));
DFFX1 gate728(.Q (g2567), .QB (line728), .D(g34021), .CK(clk));
DFFX1 gate729(.Q (g568), .QB (line729), .D(g26895), .CK(clk));
DFFX1 gate730(.Q (g3263), .QB (line730), .D(g30413), .CK(clk));
DFFX1 gate731(.Q (g6613), .QB (line731), .D(g30549), .CK(clk));
DFFX1 gate732(.Q (g6044), .QB (line732), .D(g24347), .CK(clk));
DFFX1 gate733(.Q (g6444), .QB (line733), .D(g25758), .CK(clk));
DFFX1 gate734(.Q (g2965), .QB (line734), .D(g34808), .CK(clk));
DFFX1 gate735(.Q (g5857), .QB (line735), .D(g30501), .CK(clk));
DFFX1 gate736(.Q (g1616), .QB (line736), .D(g33969), .CK(clk));
DFFX1 gate737(.Q (g890), .QB (line737), .D(g34440), .CK(clk));
DFFX1 gate738(.Q (g5976), .QB (line738), .D(g5969), .CK(clk));
DFFX1 gate739(.Q (g3562), .QB (line739), .D(g30433), .CK(clk));
DFFX1 gate740(.Q (g4294), .QB (line740), .D(g21900), .CK(clk));
DFFX1 gate741(.Q (g1404), .QB (line741), .D(g26921), .CK(clk));
DFFX1 gate742(.Q (g3723), .QB (line742), .D(g31893), .CK(clk));
DFFX1 gate743(.Q (g3817), .QB (line743), .D(g29270), .CK(clk));
DFFX1 gate744(.Q (g93), .QB (line744), .D(g34878), .CK(clk));
DFFX1 gate745(.Q (g4501), .QB (line745), .D(g33038), .CK(clk));
DFFX1 gate746(.Q (g287), .QB (line746), .D(g31865), .CK(clk));
DFFX1 gate747(.Q (g2724), .QB (line747), .D(g26926), .CK(clk));
DFFX1 gate748(.Q (g4704), .QB (line748), .D(g28083), .CK(clk));
DFFX1 gate749(.Q (g22), .QB (line749), .D(g29209), .CK(clk));
DFFX1 gate750(.Q (g2878), .QB (line750), .D(g34797), .CK(clk));
DFFX1 gate751(.Q (g5220), .QB (line751), .D(g30478), .CK(clk));
DFFX1 gate752(.Q (g617), .QB (line752), .D(g34724), .CK(clk));
DFFX1 gate753(.Q (g637), .QB (line753), .D(g24212), .CK(clk));
DFFX1 gate754(.Q (g316), .QB (line754), .D(g26883), .CK(clk));
DFFX1 gate755(.Q (g1277), .QB (line755), .D(g32985), .CK(clk));
DFFX1 gate756(.Q (g6513), .QB (line756), .D(g25761), .CK(clk));
DFFX1 gate757(.Q (g336), .QB (line757), .D(g26886), .CK(clk));
DFFX1 gate758(.Q (g2882), .QB (line758), .D(g34796), .CK(clk));
DFFX1 gate759(.Q (g933), .QB (line759), .D(g32982), .CK(clk));
DFFX1 gate760(.Q (g1906), .QB (line760), .D(g33561), .CK(clk));
DFFX1 gate761(.Q (g305), .QB (line761), .D(g26880), .CK(clk));
DFFX1 gate762(.Q (g8), .QB (line762), .D(g34591), .CK(clk));
DFFX1 gate763(.Q (g3368), .QB (line763), .D(g31884), .CK(clk));
DFFX1 gate764(.Q (g2799), .QB (line764), .D(g26931), .CK(clk));
DFFX1 gate765(.Q (g887), .QB (line765), .D(g884), .CK(clk));
DFFX1 gate766(.Q (g5327), .QB (line766), .D(g5308), .CK(clk));
DFFX1 gate767(.Q (g4912), .QB (line767), .D(g34641), .CK(clk));
DFFX1 gate768(.Q (g4157), .QB (line768), .D(g34629), .CK(clk));
DFFX1 gate769(.Q (g2541), .QB (line769), .D(g33598), .CK(clk));
DFFX1 gate770(.Q (g2153), .QB (line770), .D(g33576), .CK(clk));
DFFX1 gate771(.Q (g550), .QB (line771), .D(g34720), .CK(clk));
DFFX1 gate772(.Q (g255), .QB (line772), .D(g26902), .CK(clk));
DFFX1 gate773(.Q (g1945), .QB (line773), .D(g29244), .CK(clk));
DFFX1 gate774(.Q (g5240), .QB (line774), .D(g30468), .CK(clk));
DFFX1 gate775(.Q (g1478), .QB (line775), .D(g26924), .CK(clk));
DFFX1 gate776(.Q (g3080), .QB (line776), .D(g25645), .CK(clk));
DFFX1 gate777(.Q (g3863), .QB (line777), .D(g33031), .CK(clk));
DFFX1 gate778(.Q (g1959), .QB (line778), .D(g29245), .CK(clk));
DFFX1 gate779(.Q (g3480), .QB (line779), .D(g29266), .CK(clk));
DFFX1 gate780(.Q (g6653), .QB (line780), .D(g30559), .CK(clk));
DFFX1 gate781(.Q (g6719), .QB (line781), .D(g6715), .CK(clk));
DFFX1 gate782(.Q (g2864), .QB (line782), .D(g34794), .CK(clk));
DFFX1 gate783(.Q (g4894), .QB (line783), .D(g28087), .CK(clk));
DFFX1 gate784(.Q (g5681), .QB (line784), .D(g5677), .CK(clk));
DFFX1 gate785(.Q (g3857), .QB (line785), .D(g30435), .CK(clk));
DFFX1 gate786(.Q (g3976), .QB (line786), .D(g3969), .CK(clk));
DFFX1 gate787(.Q (g499), .QB (line787), .D(g25609), .CK(clk));
DFFX1 gate788(.Q (g5413), .QB (line788), .D(g28095), .CK(clk));
DFFX1 gate789(.Q (g1002), .QB (line789), .D(g28057), .CK(clk));
DFFX1 gate790(.Q (g776), .QB (line790), .D(g34439), .CK(clk));
DFFX1 gate791(.Q (g28), .QB (line791), .D(g34595), .CK(clk));
DFFX1 gate792(.Q (g1236), .QB (line792), .D(g1233), .CK(clk));
DFFX1 gate793(.Q (g4646), .QB (line793), .D(g34260), .CK(clk));
DFFX1 gate794(.Q (g2476), .QB (line794), .D(g33012), .CK(clk));
DFFX1 gate795(.Q (g1657), .QB (line795), .D(g32989), .CK(clk));
DFFX1 gate796(.Q (g2375), .QB (line796), .D(g34006), .CK(clk));
DFFX1 gate797(.Q (g63), .QB (line797), .D(g34847), .CK(clk));
DFFX1 gate798(.Q (g6012), .QB (line798), .D(g5983), .CK(clk));
DFFX1 gate799(.Q (g358), .QB (line799), .D(g365), .CK(clk));
DFFX1 gate800(.Q (g896), .QB (line800), .D(g26910), .CK(clk));
DFFX1 gate801(.Q (g967), .QB (line801), .D(g21722), .CK(clk));
DFFX1 gate802(.Q (g3423), .QB (line802), .D(g25658), .CK(clk));
DFFX1 gate803(.Q (g283), .QB (line803), .D(g28043), .CK(clk));
DFFX1 gate804(.Q (g3161), .QB (line804), .D(g33021), .CK(clk));
DFFX1 gate805(.Q (g2384), .QB (line805), .D(g29251), .CK(clk));
DFFX1 gate806(.Q (g3361), .QB (line806), .D(g25665), .CK(clk));
DFFX1 gate807(.Q (g6675), .QB (line807), .D(g6697), .CK(clk));
DFFX1 gate808(.Q (g4616), .QB (line808), .D(g34456), .CK(clk));
DFFX1 gate809(.Q (g4561), .QB (line809), .D(g26968), .CK(clk));
DFFX1 gate810(.Q (g2024), .QB (line810), .D(g33991), .CK(clk));
DFFX1 gate811(.Q (g3451), .QB (line811), .D(g3443), .CK(clk));
DFFX1 gate812(.Q (g2795), .QB (line812), .D(g26930), .CK(clk));
DFFX1 gate813(.Q (g613), .QB (line813), .D(g34599), .CK(clk));
DFFX1 gate814(.Q (g4527), .QB (line814), .D(g28082), .CK(clk));
DFFX1 gate815(.Q (g1844), .QB (line815), .D(g33557), .CK(clk));
DFFX1 gate816(.Q (g5937), .QB (line816), .D(g30511), .CK(clk));
DFFX1 gate817(.Q (g4546), .QB (line817), .D(g33045), .CK(clk));
DFFX1 gate818(.Q (g3103), .QB (line818), .D(g3096), .CK(clk));
DFFX1 gate819(.Q (g2523), .QB (line819), .D(g30379), .CK(clk));
DFFX1 gate820(.Q (g3303), .QB (line820), .D(g24267), .CK(clk));
DFFX1 gate821(.Q (g2643), .QB (line821), .D(g34020), .CK(clk));
DFFX1 gate822(.Q (g6109), .QB (line822), .D(g28100), .CK(clk));
DFFX1 gate823(.Q (g1489), .QB (line823), .D(g24249), .CK(clk));
DFFX1 gate824(.Q (g5390), .QB (line824), .D(g31908), .CK(clk));
DFFX1 gate825(.Q (g194), .QB (line825), .D(g25592), .CK(clk));
DFFX1 gate826(.Q (g2551), .QB (line826), .D(g30382), .CK(clk));
DFFX1 gate827(.Q (g5156), .QB (line827), .D(g29285), .CK(clk));
DFFX1 gate828(.Q (g3072), .QB (line828), .D(g25644), .CK(clk));
DFFX1 gate829(.Q (g1242), .QB (line829), .D(g1227), .CK(clk));
DFFX1 gate830(.Q (g47), .QB (line830), .D(g34992), .CK(clk));
DFFX1 gate831(.Q (g3443), .QB (line831), .D(g25662), .CK(clk));
DFFX1 gate832(.Q (g4277), .QB (line832), .D(g21896), .CK(clk));
DFFX1 gate833(.Q (g1955), .QB (line833), .D(g33563), .CK(clk));
DFFX1 gate834(.Q (g6049), .QB (line834), .D(g33622), .CK(clk));
DFFX1 gate835(.Q (g3034), .QB (line835), .D(g31876), .CK(clk));
DFFX1 gate836(.Q (g2273), .QB (line836), .D(g33582), .CK(clk));
DFFX1 gate837(.Q (g6715), .QB (line837), .D(g6711), .CK(clk));
DFFX1 gate838(.Q (g4771), .QB (line838), .D(g28086), .CK(clk));
DFFX1 gate839(.Q (g6098), .QB (line839), .D(g25744), .CK(clk));
DFFX1 gate840(.Q (g3147), .QB (line840), .D(g29262), .CK(clk));
DFFX1 gate841(.Q (g3347), .QB (line841), .D(g24270), .CK(clk));
DFFX1 gate842(.Q (g2269), .QB (line842), .D(g33581), .CK(clk));
DFFX1 gate843(.Q (g191), .QB (line843), .D(g194), .CK(clk));
DFFX1 gate844(.Q (g2712), .QB (line844), .D(g26937), .CK(clk));
DFFX1 gate845(.Q (g626), .QB (line845), .D(g34849), .CK(clk));
DFFX1 gate846(.Q (g2729), .QB (line846), .D(g28060), .CK(clk));
DFFX1 gate847(.Q (g5357), .QB (line847), .D(g33618), .CK(clk));
DFFX1 gate848(.Q (g4991), .QB (line848), .D(g34038), .CK(clk));
DFFX1 gate849(.Q (g6019), .QB (line849), .D(g6000), .CK(clk));
DFFX1 gate850(.Q (g4709), .QB (line850), .D(g34032), .CK(clk));
DFFX1 gate851(.Q (g6419), .QB (line851), .D(g31927), .CK(clk));
DFFX1 gate852(.Q (g6052), .QB (line852), .D(g31919), .CK(clk));
DFFX1 gate853(.Q (g2927), .QB (line853), .D(g34803), .CK(clk));
DFFX1 gate854(.Q (g4340), .QB (line854), .D(g34459), .CK(clk));
DFFX1 gate855(.Q (g5929), .QB (line855), .D(g30509), .CK(clk));
DFFX1 gate856(.Q (g4907), .QB (line856), .D(g34640), .CK(clk));
DFFX1 gate857(.Q (g3317), .QB (line857), .D(g3298), .CK(clk));
DFFX1 gate858(.Q (g4035), .QB (line858), .D(g28069), .CK(clk));
DFFX1 gate859(.Q (g2946), .QB (line859), .D(g21899), .CK(clk));
DFFX1 gate860(.Q (g918), .QB (line860), .D(g31868), .CK(clk));
DFFX1 gate861(.Q (g4082), .QB (line861), .D(g26938), .CK(clk));
DFFX1 gate862(.Q (g6486), .QB (line862), .D(g25756), .CK(clk));
DFFX1 gate863(.Q (g2036), .QB (line863), .D(g30363), .CK(clk));
DFFX1 gate864(.Q (g577), .QB (line864), .D(g30334), .CK(clk));
DFFX1 gate865(.Q (g1620), .QB (line865), .D(g33970), .CK(clk));
DFFX1 gate866(.Q (g2831), .QB (line866), .D(g30391), .CK(clk));
DFFX1 gate867(.Q (g667), .QB (line867), .D(g25615), .CK(clk));
DFFX1 gate868(.Q (g930), .QB (line868), .D(g33540), .CK(clk));
DFFX1 gate869(.Q (g3937), .QB (line869), .D(g30445), .CK(clk));
DFFX1 gate870(.Q (g5782), .QB (line870), .D(g25725), .CK(clk));
DFFX1 gate871(.Q (g817), .QB (line871), .D(g25617), .CK(clk));
DFFX1 gate872(.Q (g1249), .QB (line872), .D(g24247), .CK(clk));
DFFX1 gate873(.Q (g837), .QB (line873), .D(g24215), .CK(clk));
DFFX1 gate874(.Q (g3668), .QB (line874), .D(g3649), .CK(clk));
DFFX1 gate875(.Q (g599), .QB (line875), .D(g33964), .CK(clk));
DFFX1 gate876(.Q (g5475), .QB (line876), .D(g25719), .CK(clk));
DFFX1 gate877(.Q (g739), .QB (line877), .D(g29228), .CK(clk));
DFFX1 gate878(.Q (g5949), .QB (line878), .D(g30514), .CK(clk));
DFFX1 gate879(.Q (g6682), .QB (line879), .D(g33627), .CK(clk));
DFFX1 gate880(.Q (g6105), .QB (line880), .D(g28101), .CK(clk));
DFFX1 gate881(.Q (g904), .QB (line881), .D(g24231), .CK(clk));
DFFX1 gate882(.Q (g2873), .QB (line882), .D(g34615), .CK(clk));
DFFX1 gate883(.Q (g1854), .QB (line883), .D(g30356), .CK(clk));
DFFX1 gate884(.Q (g5084), .QB (line884), .D(g25696), .CK(clk));
DFFX1 gate885(.Q (g5603), .QB (line885), .D(g30493), .CK(clk));
DFFX1 gate886(.Q (g4222), .QB (line886), .D(g4219), .CK(clk));
DFFX1 gate887(.Q (g2495), .QB (line887), .D(g33594), .CK(clk));
DFFX1 gate888(.Q (g2437), .QB (line888), .D(g34009), .CK(clk));
DFFX1 gate889(.Q (g2102), .QB (line889), .D(g30365), .CK(clk));
DFFX1 gate890(.Q (g2208), .QB (line890), .D(g33004), .CK(clk));
DFFX1 gate891(.Q (g2579), .QB (line891), .D(g34018), .CK(clk));
DFFX1 gate892(.Q (g4064), .QB (line892), .D(g25685), .CK(clk));
DFFX1 gate893(.Q (g4899), .QB (line893), .D(g34040), .CK(clk));
DFFX1 gate894(.Q (g2719), .QB (line894), .D(g25639), .CK(clk));
DFFX1 gate895(.Q (g4785), .QB (line895), .D(g34029), .CK(clk));
DFFX1 gate896(.Q (g5583), .QB (line896), .D(g30488), .CK(clk));
DFFX1 gate897(.Q (g781), .QB (line897), .D(g34600), .CK(clk));
DFFX1 gate898(.Q (g6173), .QB (line898), .D(g29300), .CK(clk));
DFFX1 gate899(.Q (g6373), .QB (line899), .D(g6369), .CK(clk));
DFFX1 gate900(.Q (g2917), .QB (line900), .D(g34802), .CK(clk));
DFFX1 gate901(.Q (g686), .QB (line901), .D(g25614), .CK(clk));
DFFX1 gate902(.Q (g1252), .QB (line902), .D(g28058), .CK(clk));
DFFX1 gate903(.Q (g671), .QB (line903), .D(g29225), .CK(clk));
DFFX1 gate904(.Q (g2265), .QB (line904), .D(g33580), .CK(clk));
DFFX1 gate905(.Q (g6283), .QB (line905), .D(g30532), .CK(clk));
DFFX1 gate906(.Q (g6369), .QB (line906), .D(g6365), .CK(clk));
DFFX1 gate907(.Q (g5276), .QB (line907), .D(g5320), .CK(clk));
DFFX1 gate908(.Q (g6459), .QB (line908), .D(g25760), .CK(clk));
DFFX1 gate909(.Q (g901), .QB (line909), .D(g25620), .CK(clk));
DFFX1 gate910(.Q (g4194), .QB (line910), .D(g4188), .CK(clk));
DFFX1 gate911(.Q (g5527), .QB (line911), .D(g33054), .CK(clk));
DFFX1 gate912(.Q (g4489), .QB (line912), .D(g26962), .CK(clk));
DFFX1 gate913(.Q (g1974), .QB (line913), .D(g33564), .CK(clk));
DFFX1 gate914(.Q (g1270), .QB (line914), .D(g32984), .CK(clk));
DFFX1 gate915(.Q (g4966), .QB (line915), .D(g34039), .CK(clk));
DFFX1 gate916(.Q (g6415), .QB (line916), .D(g31932), .CK(clk));
DFFX1 gate917(.Q (g6227), .QB (line917), .D(g33065), .CK(clk));
DFFX1 gate918(.Q (g3929), .QB (line918), .D(g30443), .CK(clk));
DFFX1 gate919(.Q (g5503), .QB (line919), .D(g29291), .CK(clk));
DFFX1 gate920(.Q (g4242), .QB (line920), .D(g24279), .CK(clk));
DFFX1 gate921(.Q (g5925), .QB (line921), .D(g30508), .CK(clk));
DFFX1 gate922(.Q (g1124), .QB (line922), .D(g29232), .CK(clk));
DFFX1 gate923(.Q (g4955), .QB (line923), .D(g34269), .CK(clk));
DFFX1 gate924(.Q (g5224), .QB (line924), .D(g30464), .CK(clk));
DFFX1 gate925(.Q (g2012), .QB (line925), .D(g33988), .CK(clk));
DFFX1 gate926(.Q (g6203), .QB (line926), .D(g30522), .CK(clk));
DFFX1 gate927(.Q (g5120), .QB (line927), .D(g25708), .CK(clk));
DFFX1 gate928(.Q (g5320), .QB (line928), .D(g5290), .CK(clk));
DFFX1 gate929(.Q (g2389), .QB (line929), .D(g30374), .CK(clk));
DFFX1 gate930(.Q (g4438), .QB (line930), .D(g26953), .CK(clk));
DFFX1 gate931(.Q (g2429), .QB (line931), .D(g34008), .CK(clk));
DFFX1 gate932(.Q (g2787), .QB (line932), .D(g34444), .CK(clk));
DFFX1 gate933(.Q (g1287), .QB (line933), .D(g34731), .CK(clk));
DFFX1 gate934(.Q (g2675), .QB (line934), .D(g33606), .CK(clk));
DFFX1 gate935(.Q (g66), .QB (line935), .D(g24334), .CK(clk));
DFFX1 gate936(.Q (g4836), .QB (line936), .D(g34265), .CK(clk));
DFFX1 gate937(.Q (g1199), .QB (line937), .D(g30340), .CK(clk));
DFFX1 gate938(.Q (g1399), .QB (line938), .D(g24257), .CK(clk));
DFFX1 gate939(.Q (g5547), .QB (line939), .D(g30482), .CK(clk));
DFFX1 gate940(.Q (g3782), .QB (line940), .D(g25673), .CK(clk));
DFFX1 gate941(.Q (g6428), .QB (line941), .D(g31929), .CK(clk));
DFFX1 gate942(.Q (g2138), .QB (line942), .D(g34604), .CK(clk));
DFFX1 gate943(.Q (g3661), .QB (line943), .D(g3632), .CK(clk));
DFFX1 gate944(.Q (g2338), .QB (line944), .D(g33591), .CK(clk));
DFFX1 gate945(.Q (g4229), .QB (line945), .D(g4226), .CK(clk));
DFFX1 gate946(.Q (g6247), .QB (line946), .D(g30525), .CK(clk));
DFFX1 gate947(.Q (g2791), .QB (line947), .D(g26929), .CK(clk));
DFFX1 gate948(.Q (g3949), .QB (line948), .D(g30448), .CK(clk));
DFFX1 gate949(.Q (g1291), .QB (line949), .D(g34602), .CK(clk));
DFFX1 gate950(.Q (g5945), .QB (line950), .D(g30513), .CK(clk));
DFFX1 gate951(.Q (g5244), .QB (line951), .D(g30469), .CK(clk));
DFFX1 gate952(.Q (g2759), .QB (line952), .D(g33608), .CK(clk));
DFFX1 gate953(.Q (g6741), .QB (line953), .D(g33626), .CK(clk));
DFFX1 gate954(.Q (g785), .QB (line954), .D(g34725), .CK(clk));
DFFX1 gate955(.Q (g1259), .QB (line955), .D(g30342), .CK(clk));
DFFX1 gate956(.Q (g3484), .QB (line956), .D(g29267), .CK(clk));
DFFX1 gate957(.Q (g209), .QB (line957), .D(g25593), .CK(clk));
DFFX1 gate958(.Q (g6609), .QB (line958), .D(g30548), .CK(clk));
DFFX1 gate959(.Q (g5517), .QB (line959), .D(g33052), .CK(clk));
DFFX1 gate960(.Q (g2449), .QB (line960), .D(g34012), .CK(clk));
DFFX1 gate961(.Q (g2575), .QB (line961), .D(g34017), .CK(clk));
DFFX1 gate962(.Q (g65), .QB (line962), .D(g34785), .CK(clk));
DFFX1 gate963(.Q (g2715), .QB (line963), .D(g24263), .CK(clk));
DFFX1 gate964(.Q (g936), .QB (line964), .D(g26912), .CK(clk));
DFFX1 gate965(.Q (g2098), .QB (line965), .D(g30364), .CK(clk));
DFFX1 gate966(.Q (g4462), .QB (line966), .D(g34254), .CK(clk));
DFFX1 gate967(.Q (g604), .QB (line967), .D(g34251), .CK(clk));
DFFX1 gate968(.Q (g6589), .QB (line968), .D(g30560), .CK(clk));
DFFX1 gate969(.Q (g1886), .QB (line969), .D(g33983), .CK(clk));
DFFX1 gate970(.Q (g6466), .QB (line970), .D(g25752), .CK(clk));
DFFX1 gate971(.Q (g6365), .QB (line971), .D(g6346), .CK(clk));
DFFX1 gate972(.Q (g6711), .QB (line972), .D(g6692), .CK(clk));
DFFX1 gate973(.Q (g429), .QB (line973), .D(g24204), .CK(clk));
DFFX1 gate974(.Q (g1870), .QB (line974), .D(g33980), .CK(clk));
DFFX1 gate975(.Q (g4249), .QB (line975), .D(g34631), .CK(clk));
DFFX1 gate976(.Q (g6455), .QB (line976), .D(g28103), .CK(clk));
DFFX1 gate977(.Q (g3004), .QB (line977), .D(g31873), .CK(clk));
DFFX1 gate978(.Q (g1825), .QB (line978), .D(g29243), .CK(clk));
DFFX1 gate979(.Q (g6133), .QB (line979), .D(g25740), .CK(clk));
DFFX1 gate980(.Q (g1008), .QB (line980), .D(g25623), .CK(clk));
DFFX1 gate981(.Q (g4392), .QB (line981), .D(g26950), .CK(clk));
DFFX1 gate982(.Q (g5002), .QB (line982), .D(g4999), .CK(clk));
DFFX1 gate983(.Q (g3546), .QB (line983), .D(g30431), .CK(clk));
DFFX1 gate984(.Q (g5236), .QB (line984), .D(g30467), .CK(clk));
DFFX1 gate985(.Q (g1768), .QB (line985), .D(g30353), .CK(clk));
DFFX1 gate986(.Q (g4854), .QB (line986), .D(g34467), .CK(clk));
DFFX1 gate987(.Q (g3925), .QB (line987), .D(g30442), .CK(clk));
DFFX1 gate988(.Q (g6509), .QB (line988), .D(g29305), .CK(clk));
DFFX1 gate989(.Q (g732), .QB (line989), .D(g25616), .CK(clk));
DFFX1 gate990(.Q (g2504), .QB (line990), .D(g29252), .CK(clk));
DFFX1 gate991(.Q (g1322), .QB (line991), .D(g1459), .CK(clk));
DFFX1 gate992(.Q (g4520), .QB (line992), .D(g6972), .CK(clk));
DFFX1 gate993(.Q (g4219), .QB (line993), .D(g4216), .CK(clk));
DFFX1 gate994(.Q (g2185), .QB (line994), .D(g33003), .CK(clk));
DFFX1 gate995(.Q (g37), .QB (line995), .D(g34613), .CK(clk));
DFFX1 gate996(.Q (g4031), .QB (line996), .D(g4027), .CK(clk));
DFFX1 gate997(.Q (g2070), .QB (line997), .D(g33570), .CK(clk));
DFFX1 gate998(.Q (g4812), .QB (line998), .D(g4809), .CK(clk));
DFFX1 gate999(.Q (g6093), .QB (line999), .D(g33061), .CK(clk));
DFFX1 gate1000(.Q (g968), .QB (line1000), .D(g21723), .CK(clk));
DFFX1 gate1001(.Q (g4176), .QB (line1001), .D(g34734), .CK(clk));
DFFX1 gate1002(.Q (g4005), .QB (line1002), .D(g24275), .CK(clk));
DFFX1 gate1003(.Q (g4405), .QB (line1003), .D(g4408), .CK(clk));
DFFX1 gate1004(.Q (g872), .QB (line1004), .D(g887), .CK(clk));
DFFX1 gate1005(.Q (g6181), .QB (line1005), .D(g29302), .CK(clk));
DFFX1 gate1006(.Q (g6381), .QB (line1006), .D(g24349), .CK(clk));
DFFX1 gate1007(.Q (g4765), .QB (line1007), .D(g34264), .CK(clk));
DFFX1 gate1008(.Q (g5563), .QB (line1008), .D(g30484), .CK(clk));
DFFX1 gate1009(.Q (g1395), .QB (line1009), .D(g25634), .CK(clk));
DFFX1 gate1010(.Q (g1913), .QB (line1010), .D(g33567), .CK(clk));
DFFX1 gate1011(.Q (g2331), .QB (line1011), .D(g33585), .CK(clk));
DFFX1 gate1012(.Q (g6263), .QB (line1012), .D(g30527), .CK(clk));
DFFX1 gate1013(.Q (g50), .QB (line1013), .D(g34995), .CK(clk));
DFFX1 gate1014(.Q (g3945), .QB (line1014), .D(g30447), .CK(clk));
DFFX1 gate1015(.Q (g347), .QB (line1015), .D(g344), .CK(clk));
DFFX1 gate1016(.Q (g5731), .QB (line1016), .D(g31914), .CK(clk));
DFFX1 gate1017(.Q (g4473), .QB (line1017), .D(g34256), .CK(clk));
DFFX1 gate1018(.Q (g1266), .QB (line1018), .D(g25630), .CK(clk));
DFFX1 gate1019(.Q (g5489), .QB (line1019), .D(g29290), .CK(clk));
DFFX1 gate1020(.Q (g714), .QB (line1020), .D(g29227), .CK(clk));
DFFX1 gate1021(.Q (g2748), .QB (line1021), .D(g31872), .CK(clk));
DFFX1 gate1022(.Q (g5471), .QB (line1022), .D(g29287), .CK(clk));
DFFX1 gate1023(.Q (g4540), .QB (line1023), .D(g31897), .CK(clk));
DFFX1 gate1024(.Q (g6723), .QB (line1024), .D(g6719), .CK(clk));
DFFX1 gate1025(.Q (g6605), .QB (line1025), .D(g30562), .CK(clk));
DFFX1 gate1026(.Q (g2445), .QB (line1026), .D(g34011), .CK(clk));
DFFX1 gate1027(.Q (g2173), .QB (line1027), .D(g33996), .CK(clk));
DFFX1 gate1028(.Q (g4287), .QB (line1028), .D(g21898), .CK(clk));
DFFX1 gate1029(.Q (g2491), .QB (line1029), .D(g33014), .CK(clk));
DFFX1 gate1030(.Q (g4849), .QB (line1030), .D(g34465), .CK(clk));
DFFX1 gate1031(.Q (g2169), .QB (line1031), .D(g33995), .CK(clk));
DFFX1 gate1032(.Q (g2283), .QB (line1032), .D(g30372), .CK(clk));
DFFX1 gate1033(.Q (g6585), .QB (line1033), .D(g30545), .CK(clk));
DFFX1 gate1034(.Q (g121), .QB (line1034), .D(g30389), .CK(clk));
DFFX1 gate1035(.Q (g2407), .QB (line1035), .D(g33590), .CK(clk));
DFFX1 gate1036(.Q (g2868), .QB (line1036), .D(g34616), .CK(clk));
DFFX1 gate1037(.Q (g2767), .QB (line1037), .D(g26927), .CK(clk));
DFFX1 gate1038(.Q (g1783), .QB (line1038), .D(g32992), .CK(clk));
DFFX1 gate1039(.Q (g3310), .QB (line1039), .D(g3281), .CK(clk));
DFFX1 gate1040(.Q (g1312), .QB (line1040), .D(g25631), .CK(clk));
DFFX1 gate1041(.Q (g5212), .QB (line1041), .D(g30477), .CK(clk));
DFFX1 gate1042(.Q (g4245), .QB (line1042), .D(g34632), .CK(clk));
DFFX1 gate1043(.Q (g645), .QB (line1043), .D(g28046), .CK(clk));
DFFX1 gate1044(.Q (g4291), .QB (line1044), .D(g4287), .CK(clk));
DFFX1 gate1045(.Q (g79), .QB (line1045), .D(g26896), .CK(clk));
DFFX1 gate1046(.Q (g182), .QB (line1046), .D(g25602), .CK(clk));
DFFX1 gate1047(.Q (g1129), .QB (line1047), .D(g26916), .CK(clk));
DFFX1 gate1048(.Q (g2227), .QB (line1048), .D(g33578), .CK(clk));
DFFX1 gate1049(.Q (g6058), .QB (line1049), .D(g25745), .CK(clk));
DFFX1 gate1050(.Q (g4207), .QB (line1050), .D(g4204), .CK(clk));
DFFX1 gate1051(.Q (g2246), .QB (line1051), .D(g33579), .CK(clk));
DFFX1 gate1052(.Q (g1830), .QB (line1052), .D(g30354), .CK(clk));
DFFX1 gate1053(.Q (g3590), .QB (line1053), .D(g30425), .CK(clk));
DFFX1 gate1054(.Q (g392), .QB (line1054), .D(g24200), .CK(clk));
DFFX1 gate1055(.Q (g1592), .QB (line1055), .D(g33544), .CK(clk));
DFFX1 gate1056(.Q (g6505), .QB (line1056), .D(g25764), .CK(clk));
DFFX1 gate1057(.Q (g6411), .QB (line1057), .D(g31930), .CK(clk));
DFFX1 gate1058(.Q (g1221), .QB (line1058), .D(g24246), .CK(clk));
DFFX1 gate1059(.Q (g5921), .QB (line1059), .D(g30507), .CK(clk));
DFFX1 gate1060(.Q (g106), .QB (line1060), .D(g26889), .CK(clk));
DFFX1 gate1061(.Q (g146), .QB (line1061), .D(g30333), .CK(clk));
DFFX1 gate1062(.Q (g218), .QB (line1062), .D(g215), .CK(clk));
DFFX1 gate1063(.Q (g6474), .QB (line1063), .D(g25753), .CK(clk));
DFFX1 gate1064(.Q (g1932), .QB (line1064), .D(g32998), .CK(clk));
DFFX1 gate1065(.Q (g1624), .QB (line1065), .D(g32987), .CK(clk));
DFFX1 gate1066(.Q (g5062), .QB (line1066), .D(g25702), .CK(clk));
DFFX1 gate1067(.Q (g5462), .QB (line1067), .D(g29286), .CK(clk));
DFFX1 gate1068(.Q (g2689), .QB (line1068), .D(g34606), .CK(clk));
DFFX1 gate1069(.Q (g6573), .QB (line1069), .D(g33070), .CK(clk));
DFFX1 gate1070(.Q (g1677), .QB (line1070), .D(g29240), .CK(clk));
DFFX1 gate1071(.Q (g2028), .QB (line1071), .D(g32999), .CK(clk));
DFFX1 gate1072(.Q (g2671), .QB (line1072), .D(g33605), .CK(clk));
DFFX1 gate1073(.Q (g1576), .QB (line1073), .D(g24255), .CK(clk));
DFFX1 gate1074(.Q (g4408), .QB (line1074), .D(g26945), .CK(clk));
DFFX1 gate1075(.Q (g34), .QB (line1075), .D(g34877), .CK(clk));
DFFX1 gate1076(.Q (g1848), .QB (line1076), .D(g33558), .CK(clk));
DFFX1 gate1077(.Q (g3089), .QB (line1077), .D(g25647), .CK(clk));
DFFX1 gate1078(.Q (g3731), .QB (line1078), .D(g31889), .CK(clk));
DFFX1 gate1079(.Q (g86), .QB (line1079), .D(g25699), .CK(clk));
DFFX1 gate1080(.Q (g5485), .QB (line1080), .D(g29289), .CK(clk));
DFFX1 gate1081(.Q (g2741), .QB (line1081), .D(g30388), .CK(clk));
DFFX1 gate1082(.Q (g802), .QB (line1082), .D(g799), .CK(clk));
DFFX1 gate1083(.Q (g2638), .QB (line1083), .D(g29254), .CK(clk));
DFFX1 gate1084(.Q (g4122), .QB (line1084), .D(g28074), .CK(clk));
DFFX1 gate1085(.Q (g4322), .QB (line1085), .D(g34450), .CK(clk));
DFFX1 gate1086(.Q (g5941), .QB (line1086), .D(g30512), .CK(clk));
DFFX1 gate1087(.Q (g2108), .QB (line1087), .D(g33572), .CK(clk));
DFFX1 gate1088(.Q (g6000), .QB (line1088), .D(g5976), .CK(clk));
DFFX1 gate1089(.Q (g25), .QB (line1089), .D(g15048), .CK(clk));
DFFX1 gate1090(.Q (g1644), .QB (line1090), .D(g33551), .CK(clk));
DFFX1 gate1091(.Q (g595), .QB (line1091), .D(g33538), .CK(clk));
DFFX1 gate1092(.Q (g2217), .QB (line1092), .D(g33005), .CK(clk));
DFFX1 gate1093(.Q (g1319), .QB (line1093), .D(g24248), .CK(clk));
DFFX1 gate1094(.Q (g2066), .QB (line1094), .D(g33002), .CK(clk));
DFFX1 gate1095(.Q (g1152), .QB (line1095), .D(g24234), .CK(clk));
DFFX1 gate1096(.Q (g5252), .QB (line1096), .D(g30471), .CK(clk));
DFFX1 gate1097(.Q (g2165), .QB (line1097), .D(g34000), .CK(clk));
DFFX1 gate1098(.Q (g2571), .QB (line1098), .D(g34016), .CK(clk));
DFFX1 gate1099(.Q (g5176), .QB (line1099), .D(g33048), .CK(clk));
DFFX1 gate1100(.Q (g391), .QB (line1100), .D(g26911), .CK(clk));
DFFX1 gate1101(.Q (g5005), .QB (line1101), .D(g5002), .CK(clk));
DFFX1 gate1102(.Q (g2711), .QB (line1102), .D(g18528), .CK(clk));
DFFX1 gate1103(.Q (g6023), .QB (line1103), .D(g6019), .CK(clk));
DFFX1 gate1104(.Q (g1211), .QB (line1104), .D(g25628), .CK(clk));
DFFX1 gate1105(.Q (g2827), .QB (line1105), .D(g26934), .CK(clk));
DFFX1 gate1106(.Q (g6423), .QB (line1106), .D(g31928), .CK(clk));
DFFX1 gate1107(.Q (g875), .QB (line1107), .D(g869), .CK(clk));
DFFX1 gate1108(.Q (g4859), .QB (line1108), .D(g34468), .CK(clk));
DFFX1 gate1109(.Q (g424), .QB (line1109), .D(g24202), .CK(clk));
DFFX1 gate1110(.Q (g1274), .QB (line1110), .D(g33542), .CK(clk));
DFFX1 gate1111(.Q (g1426), .QB (line1111), .D(g1422), .CK(clk));
DFFX1 gate1112(.Q (g85), .QB (line1112), .D(g34717), .CK(clk));
DFFX1 gate1113(.Q (g2803), .QB (line1113), .D(g34445), .CK(clk));
DFFX1 gate1114(.Q (g6451), .QB (line1114), .D(g28104), .CK(clk));
DFFX1 gate1115(.Q (g1821), .QB (line1115), .D(g33555), .CK(clk));
DFFX1 gate1116(.Q (g2509), .QB (line1116), .D(g34013), .CK(clk));
DFFX1 gate1117(.Q (g5073), .QB (line1117), .D(g28091), .CK(clk));
DFFX1 gate1118(.Q (g1280), .QB (line1118), .D(g26919), .CK(clk));
DFFX1 gate1119(.Q (g4815), .QB (line1119), .D(g4812), .CK(clk));
DFFX1 gate1120(.Q (g6346), .QB (line1120), .D(g6322), .CK(clk));
DFFX1 gate1121(.Q (g6633), .QB (line1121), .D(g30554), .CK(clk));
DFFX1 gate1122(.Q (g5124), .QB (line1122), .D(g29281), .CK(clk));
DFFX1 gate1123(.Q (g1083), .QB (line1123), .D(g1079), .CK(clk));
DFFX1 gate1124(.Q (g6303), .QB (line1124), .D(g30537), .CK(clk));
DFFX1 gate1125(.Q (g5069), .QB (line1125), .D(g28092), .CK(clk));
DFFX1 gate1126(.Q (g2994), .QB (line1126), .D(g34732), .CK(clk));
DFFX1 gate1127(.Q (g650), .QB (line1127), .D(g28049), .CK(clk));
DFFX1 gate1128(.Q (g1636), .QB (line1128), .D(g33545), .CK(clk));
DFFX1 gate1129(.Q (g3921), .QB (line1129), .D(g30441), .CK(clk));
DFFX1 gate1130(.Q (g2093), .QB (line1130), .D(g29247), .CK(clk));
DFFX1 gate1131(.Q (g6732), .QB (line1131), .D(g24354), .CK(clk));
DFFX1 gate1132(.Q (g1306), .QB (line1132), .D(g25636), .CK(clk));
DFFX1 gate1133(.Q (g5377), .QB (line1133), .D(g31911), .CK(clk));
DFFX1 gate1134(.Q (g1061), .QB (line1134), .D(g26914), .CK(clk));
DFFX1 gate1135(.Q (g3462), .QB (line1135), .D(g25670), .CK(clk));
DFFX1 gate1136(.Q (g2181), .QB (line1136), .D(g33998), .CK(clk));
DFFX1 gate1137(.Q (g956), .QB (line1137), .D(g25626), .CK(clk));
DFFX1 gate1138(.Q (g1756), .QB (line1138), .D(g33977), .CK(clk));
DFFX1 gate1139(.Q (g5849), .QB (line1139), .D(g29297), .CK(clk));
DFFX1 gate1140(.Q (g4112), .QB (line1140), .D(g28071), .CK(clk));
DFFX1 gate1141(.Q (g2685), .QB (line1141), .D(g30387), .CK(clk));
DFFX1 gate1142(.Q (g2197), .QB (line1142), .D(g33577), .CK(clk));
DFFX1 gate1143(.Q (g6116), .QB (line1143), .D(g25737), .CK(clk));
DFFX1 gate1144(.Q (g2421), .QB (line1144), .D(g33592), .CK(clk));
DFFX1 gate1145(.Q (g1046), .QB (line1145), .D(g26913), .CK(clk));
DFFX1 gate1146(.Q (g482), .QB (line1146), .D(g28044), .CK(clk));
DFFX1 gate1147(.Q (g4401), .QB (line1147), .D(g26948), .CK(clk));
DFFX1 gate1148(.Q (g6434), .QB (line1148), .D(g31931), .CK(clk));
DFFX1 gate1149(.Q (g1514), .QB (line1149), .D(g30344), .CK(clk));
DFFX1 gate1150(.Q (g329), .QB (line1150), .D(g26885), .CK(clk));
DFFX1 gate1151(.Q (g6565), .QB (line1151), .D(g33069), .CK(clk));
DFFX1 gate1152(.Q (g2950), .QB (line1152), .D(g34621), .CK(clk));
DFFX1 gate1153(.Q (g4129), .QB (line1153), .D(g28075), .CK(clk));
DFFX1 gate1154(.Q (g1345), .QB (line1154), .D(g28059), .CK(clk));
DFFX1 gate1155(.Q (g6533), .QB (line1155), .D(g25762), .CK(clk));
DFFX1 gate1156(.Q (g3298), .QB (line1156), .D(g3274), .CK(clk));
DFFX1 gate1157(.Q (g3085), .QB (line1157), .D(g25646), .CK(clk));
DFFX1 gate1158(.Q (g4727), .QB (line1158), .D(g34633), .CK(clk));
DFFX1 gate1159(.Q (g6697), .QB (line1159), .D(g24352), .CK(clk));
DFFX1 gate1160(.Q (g1536), .QB (line1160), .D(g26925), .CK(clk));
DFFX1 gate1161(.Q (g3941), .QB (line1161), .D(g30446), .CK(clk));
DFFX1 gate1162(.Q (g370), .QB (line1162), .D(g25597), .CK(clk));
DFFX1 gate1163(.Q (g5694), .QB (line1163), .D(g24342), .CK(clk));
DFFX1 gate1164(.Q (g1858), .QB (line1164), .D(g30357), .CK(clk));
DFFX1 gate1165(.Q (g446), .QB (line1165), .D(g26908), .CK(clk));
DFFX1 gate1166(.Q (g4932), .QB (line1166), .D(g21905), .CK(clk));
DFFX1 gate1167(.Q (g3219), .QB (line1167), .D(g30399), .CK(clk));
DFFX1 gate1168(.Q (g1811), .QB (line1168), .D(g29242), .CK(clk));
DFFX1 gate1169(.Q (g3431), .QB (line1169), .D(g25659), .CK(clk));
DFFX1 gate1170(.Q (g6601), .QB (line1170), .D(g30547), .CK(clk));
DFFX1 gate1171(.Q (g3376), .QB (line1171), .D(g31881), .CK(clk));
DFFX1 gate1172(.Q (g2441), .QB (line1172), .D(g34010), .CK(clk));
DFFX1 gate1173(.Q (g1874), .QB (line1173), .D(g33986), .CK(clk));
DFFX1 gate1174(.Q (g4349), .QB (line1174), .D(g34257), .CK(clk));
DFFX1 gate1175(.Q (g6581), .QB (line1175), .D(g30544), .CK(clk));
DFFX1 gate1176(.Q (g6597), .QB (line1176), .D(g30561), .CK(clk));
DFFX1 gate1177(.Q (g5008), .QB (line1177), .D(g5005), .CK(clk));
DFFX1 gate1178(.Q (g3610), .QB (line1178), .D(g30430), .CK(clk));
DFFX1 gate1179(.Q (g2890), .QB (line1179), .D(g34799), .CK(clk));
DFFX1 gate1180(.Q (g1978), .QB (line1180), .D(g33565), .CK(clk));
DFFX1 gate1181(.Q (g1612), .QB (line1181), .D(g33968), .CK(clk));
DFFX1 gate1182(.Q (g112), .QB (line1182), .D(g34879), .CK(clk));
DFFX1 gate1183(.Q (g2856), .QB (line1183), .D(g34793), .CK(clk));
DFFX1 gate1184(.Q (g6479), .QB (line1184), .D(g25754), .CK(clk));
DFFX1 gate1185(.Q (g1982), .QB (line1185), .D(g33566), .CK(clk));
DFFX1 gate1186(.Q (g6668), .QB (line1186), .D(g6661), .CK(clk));
DFFX1 gate1187(.Q (g5228), .QB (line1187), .D(g30465), .CK(clk));
DFFX1 gate1188(.Q (g4119), .QB (line1188), .D(g28073), .CK(clk));
DFFX1 gate1189(.Q (g6390), .QB (line1189), .D(g24351), .CK(clk));
DFFX1 gate1190(.Q (g1542), .QB (line1190), .D(g30346), .CK(clk));
DFFX1 gate1191(.Q (g4258), .QB (line1191), .D(g21893), .CK(clk));
DFFX1 gate1192(.Q (g4818), .QB (line1192), .D(g4815), .CK(clk));
DFFX1 gate1193(.Q (g5033), .QB (line1193), .D(g31904), .CK(clk));
DFFX1 gate1194(.Q (g4717), .QB (line1194), .D(g34635), .CK(clk));
DFFX1 gate1195(.Q (g1554), .QB (line1195), .D(g25637), .CK(clk));
DFFX1 gate1196(.Q (g3849), .QB (line1196), .D(g29274), .CK(clk));
DFFX1 gate1197(.Q (g6704), .QB (line1197), .D(g6675), .CK(clk));
DFFX1 gate1198(.Q (g3199), .QB (line1198), .D(g30396), .CK(clk));
DFFX1 gate1199(.Q (g5845), .QB (line1199), .D(g25735), .CK(clk));
DFFX1 gate1200(.Q (g4975), .QB (line1200), .D(g34037), .CK(clk));
DFFX1 gate1201(.Q (g790), .QB (line1201), .D(g34791), .CK(clk));
DFFX1 gate1202(.Q (g5913), .QB (line1202), .D(g30520), .CK(clk));
DFFX1 gate1203(.Q (g1902), .QB (line1203), .D(g30358), .CK(clk));
DFFX1 gate1204(.Q (g6163), .QB (line1204), .D(g29299), .CK(clk));
DFFX1 gate1205(.Q (g4125), .QB (line1205), .D(g28081), .CK(clk));
DFFX1 gate1206(.Q (g4821), .QB (line1206), .D(g28096), .CK(clk));
DFFX1 gate1207(.Q (g4939), .QB (line1207), .D(g28088), .CK(clk));
DFFX1 gate1208(.Q (g1056), .QB (line1208), .D(g24241), .CK(clk));
DFFX1 gate1209(.Q (g3207), .QB (line1209), .D(g30397), .CK(clk));
DFFX1 gate1210(.Q (g4483), .QB (line1210), .D(g4520), .CK(clk));
DFFX1 gate1211(.Q (g3259), .QB (line1211), .D(g30409), .CK(clk));
DFFX1 gate1212(.Q (g5142), .QB (line1212), .D(g29284), .CK(clk));
DFFX1 gate1213(.Q (g5248), .QB (line1213), .D(g30470), .CK(clk));
DFFX1 gate1214(.Q (g2126), .QB (line1214), .D(g30367), .CK(clk));
DFFX1 gate1215(.Q (g3694), .QB (line1215), .D(g24273), .CK(clk));
DFFX1 gate1216(.Q (g5481), .QB (line1216), .D(g29288), .CK(clk));
DFFX1 gate1217(.Q (g1964), .QB (line1217), .D(g30359), .CK(clk));
DFFX1 gate1218(.Q (g5097), .QB (line1218), .D(g25698), .CK(clk));
DFFX1 gate1219(.Q (g3215), .QB (line1219), .D(g30398), .CK(clk));
DFFX1 gate1220(.Q (g4027), .QB (line1220), .D(g4023), .CK(clk));
DFFX1 gate1221(.Q (g111), .QB (line1221), .D(g34718), .CK(clk));
DFFX1 gate1222(.Q (g4427), .QB (line1222), .D(g26952), .CK(clk));
DFFX1 gate1223(.Q (g7), .QB (line1223), .D(g34590), .CK(clk));
DFFX1 gate1224(.Q (g2779), .QB (line1224), .D(g26928), .CK(clk));
DFFX1 gate1225(.Q (g4200), .QB (line1225), .D(g4197), .CK(clk));
DFFX1 gate1226(.Q (g4446), .QB (line1226), .D(g26954), .CK(clk));
DFFX1 gate1227(.Q (g1720), .QB (line1227), .D(g30351), .CK(clk));
DFFX1 gate1228(.Q (g1367), .QB (line1228), .D(g31871), .CK(clk));
DFFX1 gate1229(.Q (g5112), .QB (line1229), .D(g5105), .CK(clk));
DFFX1 gate1230(.Q (g19), .QB (line1230), .D(g34594), .CK(clk));
DFFX1 gate1231(.Q (g4145), .QB (line1231), .D(g26939), .CK(clk));
DFFX1 gate1232(.Q (g2161), .QB (line1232), .D(g33994), .CK(clk));
DFFX1 gate1233(.Q (g376), .QB (line1233), .D(g25596), .CK(clk));
DFFX1 gate1234(.Q (g2361), .QB (line1234), .D(g33586), .CK(clk));
DFFX1 gate1235(.Q (g4191), .QB (line1235), .D(g21901), .CK(clk));
DFFX1 gate1236(.Q (g582), .QB (line1236), .D(g31866), .CK(clk));
DFFX1 gate1237(.Q (g2051), .QB (line1237), .D(g33000), .CK(clk));
DFFX1 gate1238(.Q (g1193), .QB (line1238), .D(g26918), .CK(clk));
DFFX1 gate1239(.Q (g5401), .QB (line1239), .D(g33051), .CK(clk));
DFFX1 gate1240(.Q (g3408), .QB (line1240), .D(g28065), .CK(clk));
DFFX1 gate1241(.Q (g2327), .QB (line1241), .D(g30373), .CK(clk));
DFFX1 gate1242(.Q (g907), .QB (line1242), .D(g28056), .CK(clk));
DFFX1 gate1243(.Q (g947), .QB (line1243), .D(g34601), .CK(clk));
DFFX1 gate1244(.Q (g1834), .QB (line1244), .D(g30355), .CK(clk));
DFFX1 gate1245(.Q (g3594), .QB (line1245), .D(g30426), .CK(clk));
DFFX1 gate1246(.Q (g2999), .QB (line1246), .D(g34805), .CK(clk));
DFFX1 gate1247(.Q (g5727), .QB (line1247), .D(g31913), .CK(clk));
DFFX1 gate1248(.Q (g2303), .QB (line1248), .D(g34002), .CK(clk));
DFFX1 gate1249(.Q (g6661), .QB (line1249), .D(g6704), .CK(clk));
DFFX1 gate1250(.Q (g3065), .QB (line1250), .D(g25652), .CK(clk));
DFFX1 gate1251(.Q (g699), .QB (line1251), .D(g28053), .CK(clk));
DFFX1 gate1252(.Q (g723), .QB (line1252), .D(g29229), .CK(clk));
DFFX1 gate1253(.Q (g5703), .QB (line1253), .D(g33620), .CK(clk));
DFFX1 gate1254(.Q (g546), .QB (line1254), .D(g34722), .CK(clk));
DFFX1 gate1255(.Q (g2472), .QB (line1255), .D(g33599), .CK(clk));
DFFX1 gate1256(.Q (g5953), .QB (line1256), .D(g30515), .CK(clk));
DFFX1 gate1257(.Q (g3096), .QB (line1257), .D(g25649), .CK(clk));
DFFX1 gate1258(.Q (g6439), .QB (line1258), .D(g33066), .CK(clk));
DFFX1 gate1259(.Q (g1740), .QB (line1259), .D(g33979), .CK(clk));
DFFX1 gate1260(.Q (g3550), .QB (line1260), .D(g30417), .CK(clk));
DFFX1 gate1261(.Q (g3845), .QB (line1261), .D(g25683), .CK(clk));
DFFX1 gate1262(.Q (g2116), .QB (line1262), .D(g33574), .CK(clk));
DFFX1 gate1263(.Q (g5677), .QB (line1263), .D(g5673), .CK(clk));
DFFX1 gate1264(.Q (g3195), .QB (line1264), .D(g30410), .CK(clk));
DFFX1 gate1265(.Q (g3913), .QB (line1265), .D(g30454), .CK(clk));
DFFX1 gate1266(.Q (g4537), .QB (line1266), .D(g34024), .CK(clk));
DFFX1 gate1267(.Q (g1687), .QB (line1267), .D(g33547), .CK(clk));
DFFX1 gate1268(.Q (g2681), .QB (line1268), .D(g30386), .CK(clk));
DFFX1 gate1269(.Q (g2533), .QB (line1269), .D(g33596), .CK(clk));
DFFX1 gate1270(.Q (g324), .QB (line1270), .D(g26887), .CK(clk));
DFFX1 gate1271(.Q (g2697), .QB (line1271), .D(g34607), .CK(clk));
DFFX1 gate1272(.Q (g5747), .QB (line1272), .D(g33056), .CK(clk));
DFFX1 gate1273(.Q (g4417), .QB (line1273), .D(g31895), .CK(clk));
DFFX1 gate1274(.Q (g6561), .QB (line1274), .D(g33068), .CK(clk));
DFFX1 gate1275(.Q (g1141), .QB (line1275), .D(g29233), .CK(clk));
DFFX1 gate1276(.Q (g1570), .QB (line1276), .D(g24258), .CK(clk));
DFFX1 gate1277(.Q (g2413), .QB (line1277), .D(g30376), .CK(clk));
DFFX1 gate1278(.Q (g1710), .QB (line1278), .D(g33549), .CK(clk));
DFFX1 gate1279(.Q (g6527), .QB (line1279), .D(g29308), .CK(clk));
DFFX1 gate1280(.Q (g6404), .QB (line1280), .D(g25759), .CK(clk));
DFFX1 gate1281(.Q (g3255), .QB (line1281), .D(g30408), .CK(clk));
DFFX1 gate1282(.Q (g1691), .QB (line1282), .D(g29241), .CK(clk));
DFFX1 gate1283(.Q (g2936), .QB (line1283), .D(g34620), .CK(clk));
DFFX1 gate1284(.Q (g5644), .QB (line1284), .D(g33621), .CK(clk));
DFFX1 gate1285(.Q (g5152), .QB (line1285), .D(g25707), .CK(clk));
DFFX1 gate1286(.Q (g5352), .QB (line1286), .D(g24339), .CK(clk));
DFFX1 gate1287(.Q (g4213), .QB (line1287), .D(g4185), .CK(clk));
DFFX1 gate1288(.Q (g6120), .QB (line1288), .D(g25738), .CK(clk));
DFFX1 gate1289(.Q (g2775), .QB (line1289), .D(g34443), .CK(clk));
DFFX1 gate1290(.Q (g2922), .QB (line1290), .D(g34619), .CK(clk));
DFFX1 gate1291(.Q (g1111), .QB (line1291), .D(g29234), .CK(clk));
DFFX1 gate1292(.Q (g5893), .QB (line1292), .D(g30503), .CK(clk));
DFFX1 gate1293(.Q (g1311), .QB (line1293), .D(g21724), .CK(clk));
DFFX1 gate1294(.Q (g3267), .QB (line1294), .D(g3310), .CK(clk));
DFFX1 gate1295(.Q (g6617), .QB (line1295), .D(g30550), .CK(clk));
DFFX1 gate1296(.Q (g2060), .QB (line1296), .D(g33001), .CK(clk));
DFFX1 gate1297(.Q (g4512), .QB (line1297), .D(g33040), .CK(clk));
DFFX1 gate1298(.Q (g5599), .QB (line1298), .D(g30492), .CK(clk));
DFFX1 gate1299(.Q (g3401), .QB (line1299), .D(g25664), .CK(clk));
DFFX1 gate1300(.Q (g4366), .QB (line1300), .D(g26944), .CK(clk));
DFFX1 gate1301(.Q (g3676), .QB (line1301), .D(g3672), .CK(clk));
DFFX1 gate1302(.Q (g94), .QB (line1302), .D(g34614), .CK(clk));
DFFX1 gate1303(.Q (g3129), .QB (line1303), .D(g29260), .CK(clk));
DFFX1 gate1304(.Q (g3329), .QB (line1304), .D(g3325), .CK(clk));
DFFX1 gate1305(.Q (g5170), .QB (line1305), .D(g33047), .CK(clk));
DFFX1 gate1306(.Q (g4456), .QB (line1306), .D(g25692), .CK(clk));
DFFX1 gate1307(.Q (g5821), .QB (line1307), .D(g25733), .CK(clk));
DFFX1 gate1308(.Q (g6299), .QB (line1308), .D(g30536), .CK(clk));
DFFX1 gate1309(.Q (g1239), .QB (line1309), .D(g1157), .CK(clk));
DFFX1 gate1310(.Q (g3727), .QB (line1310), .D(g31888), .CK(clk));
DFFX1 gate1311(.Q (g2079), .QB (line1311), .D(g29246), .CK(clk));
DFFX1 gate1312(.Q (g4698), .QB (line1312), .D(g34261), .CK(clk));
DFFX1 gate1313(.Q (g3703), .QB (line1313), .D(g33611), .CK(clk));
DFFX1 gate1314(.Q (g1559), .QB (line1314), .D(g25638), .CK(clk));
DFFX1 gate1315(.Q (g943), .QB (line1315), .D(g34728), .CK(clk));
DFFX1 gate1316(.Q (g411), .QB (line1316), .D(g29222), .CK(clk));
DFFX1 gate1317(.Q (g6140), .QB (line1317), .D(g25742), .CK(clk));
DFFX1 gate1318(.Q (g3953), .QB (line1318), .D(g30449), .CK(clk));
DFFX1 gate1319(.Q (g3068), .QB (line1319), .D(g25643), .CK(clk));
DFFX1 gate1320(.Q (g2704), .QB (line1320), .D(g34608), .CK(clk));
DFFX1 gate1321(.Q (g6035), .QB (line1321), .D(g24345), .CK(clk));
DFFX1 gate1322(.Q (g6082), .QB (line1322), .D(g31922), .CK(clk));
DFFX1 gate1323(.Q (g49), .QB (line1323), .D(g34994), .CK(clk));
DFFX1 gate1324(.Q (g1300), .QB (line1324), .D(g25635), .CK(clk));
DFFX1 gate1325(.Q (g4057), .QB (line1325), .D(g25686), .CK(clk));
DFFX1 gate1326(.Q (g5200), .QB (line1326), .D(g30461), .CK(clk));
DFFX1 gate1327(.Q (g4843), .QB (line1327), .D(g34466), .CK(clk));
DFFX1 gate1328(.Q (g5046), .QB (line1328), .D(g31901), .CK(clk));
DFFX1 gate1329(.Q (g2250), .QB (line1329), .D(g29249), .CK(clk));
DFFX1 gate1330(.Q (g319), .QB (line1330), .D(g26882), .CK(clk));
DFFX1 gate1331(.Q (g4549), .QB (line1331), .D(g33041), .CK(clk));
DFFX1 gate1332(.Q (g2453), .QB (line1332), .D(g33011), .CK(clk));
DFFX1 gate1333(.Q (g5841), .QB (line1333), .D(g25734), .CK(clk));
DFFX1 gate1334(.Q (g5763), .QB (line1334), .D(g28097), .CK(clk));
DFFX1 gate1335(.Q (g3747), .QB (line1335), .D(g33030), .CK(clk));
DFFX1 gate1336(.Q (g5637), .QB (line1336), .D(g5659), .CK(clk));
DFFX1 gate1337(.Q (g2912), .QB (line1337), .D(g34618), .CK(clk));
DFFX1 gate1338(.Q (g2357), .QB (line1338), .D(g33010), .CK(clk));
DFFX1 gate1339(.Q (g4232), .QB (line1339), .D(g4229), .CK(clk));
DFFX1 gate1340(.Q (g164), .QB (line1340), .D(g31864), .CK(clk));
DFFX1 gate1341(.Q (g4253), .QB (line1341), .D(g34630), .CK(clk));
DFFX1 gate1342(.Q (g5016), .QB (line1342), .D(g31898), .CK(clk));
DFFX1 gate1343(.Q (g3119), .QB (line1343), .D(g25653), .CK(clk));
DFFX1 gate1344(.Q (g1351), .QB (line1344), .D(g25632), .CK(clk));
DFFX1 gate1345(.Q (g1648), .QB (line1345), .D(g32988), .CK(clk));
DFFX1 gate1346(.Q (g4519), .QB (line1346), .D(g33616), .CK(clk));
DFFX1 gate1347(.Q (g5115), .QB (line1347), .D(g29280), .CK(clk));
DFFX1 gate1348(.Q (g3352), .QB (line1348), .D(g33609), .CK(clk));
DFFX1 gate1349(.Q (g6657), .QB (line1349), .D(g30563), .CK(clk));
DFFX1 gate1350(.Q (g4552), .QB (line1350), .D(g33044), .CK(clk));
DFFX1 gate1351(.Q (g3893), .QB (line1351), .D(g30437), .CK(clk));
DFFX1 gate1352(.Q (g3211), .QB (line1352), .D(g30412), .CK(clk));
DFFX1 gate1353(.Q (g5654), .QB (line1353), .D(g5630), .CK(clk));
DFFX1 gate1354(.Q (g929), .QB (line1354), .D(g21725), .CK(clk));
DFFX1 gate1355(.Q (g3274), .QB (line1355), .D(g3267), .CK(clk));
DFFX1 gate1356(.Q (g5595), .QB (line1356), .D(g30491), .CK(clk));
DFFX1 gate1357(.Q (g3614), .QB (line1357), .D(g30434), .CK(clk));
DFFX1 gate1358(.Q (g2894), .QB (line1358), .D(g34612), .CK(clk));
DFFX1 gate1359(.Q (g3125), .QB (line1359), .D(g29259), .CK(clk));
DFFX1 gate1360(.Q (g3325), .QB (line1360), .D(g3321), .CK(clk));
DFFX1 gate1361(.Q (g3821), .QB (line1361), .D(g25681), .CK(clk));
DFFX1 gate1362(.Q (g4141), .QB (line1362), .D(g25687), .CK(clk));
DFFX1 gate1363(.Q (g4570), .QB (line1363), .D(g33617), .CK(clk));
DFFX1 gate1364(.Q (g5272), .QB (line1364), .D(g30479), .CK(clk));
DFFX1 gate1365(.Q (g2735), .QB (line1365), .D(g29256), .CK(clk));
DFFX1 gate1366(.Q (g728), .QB (line1366), .D(g28054), .CK(clk));
DFFX1 gate1367(.Q (g6295), .QB (line1367), .D(g30535), .CK(clk));
DFFX1 gate1368(.Q (g5417), .QB (line1368), .D(g28094), .CK(clk));
DFFX1 gate1369(.Q (g2661), .QB (line1369), .D(g30385), .CK(clk));
DFFX1 gate1370(.Q (g1988), .QB (line1370), .D(g30361), .CK(clk));
DFFX1 gate1371(.Q (g5128), .QB (line1371), .D(g25705), .CK(clk));
DFFX1 gate1372(.Q (g1548), .QB (line1372), .D(g24260), .CK(clk));
DFFX1 gate1373(.Q (g3106), .QB (line1373), .D(g29257), .CK(clk));
DFFX1 gate1374(.Q (g4659), .QB (line1374), .D(g34461), .CK(clk));
DFFX1 gate1375(.Q (g4358), .QB (line1375), .D(g34258), .CK(clk));
DFFX1 gate1376(.Q (g1792), .QB (line1376), .D(g32993), .CK(clk));
DFFX1 gate1377(.Q (g2084), .QB (line1377), .D(g33992), .CK(clk));
DFFX1 gate1378(.Q (g3061), .QB (line1378), .D(g28061), .CK(clk));
DFFX1 gate1379(.Q (g3187), .QB (line1379), .D(g30394), .CK(clk));
DFFX1 gate1380(.Q (g4311), .QB (line1380), .D(g34449), .CK(clk));
DFFX1 gate1381(.Q (g2583), .QB (line1381), .D(g34019), .CK(clk));
DFFX1 gate1382(.Q (g3003), .QB (line1382), .D(g21726), .CK(clk));
DFFX1 gate1383(.Q (g1094), .QB (line1383), .D(g29231), .CK(clk));
DFFX1 gate1384(.Q (g3841), .QB (line1384), .D(g25682), .CK(clk));
DFFX1 gate1385(.Q (g4284), .QB (line1385), .D(g21897), .CK(clk));
DFFX1 gate1386(.Q (g3763), .QB (line1386), .D(g28067), .CK(clk));
DFFX1 gate1387(.Q (g3191), .QB (line1387), .D(g30395), .CK(clk));
DFFX1 gate1388(.Q (g4239), .QB (line1388), .D(g21892), .CK(clk));
DFFX1 gate1389(.Q (g3391), .QB (line1389), .D(g31885), .CK(clk));
DFFX1 gate1390(.Q (g4180), .QB (line1390), .D(g4210), .CK(clk));
DFFX1 gate1391(.Q (g691), .QB (line1391), .D(g28048), .CK(clk));
DFFX1 gate1392(.Q (g534), .QB (line1392), .D(g34723), .CK(clk));
DFFX1 gate1393(.Q (g5366), .QB (line1393), .D(g25717), .CK(clk));
DFFX1 gate1394(.Q (g385), .QB (line1394), .D(g25598), .CK(clk));
DFFX1 gate1395(.Q (g2004), .QB (line1395), .D(g33987), .CK(clk));
DFFX1 gate1396(.Q (g2527), .QB (line1396), .D(g30380), .CK(clk));
DFFX1 gate1397(.Q (g5456), .QB (line1397), .D(g5448), .CK(clk));
DFFX1 gate1398(.Q (g4420), .QB (line1398), .D(g26965), .CK(clk));
DFFX1 gate1399(.Q (g5148), .QB (line1399), .D(g25706), .CK(clk));
DFFX1 gate1400(.Q (g4507), .QB (line1400), .D(g30458), .CK(clk));
DFFX1 gate1401(.Q (g5348), .QB (line1401), .D(g24338), .CK(clk));
DFFX1 gate1402(.Q (g3223), .QB (line1402), .D(g30400), .CK(clk));
DFFX1 gate1403(.Q (g4931), .QB (line1403), .D(g21904), .CK(clk));
DFFX1 gate1404(.Q (g2970), .QB (line1404), .D(g34623), .CK(clk));
DFFX1 gate1405(.Q (g5698), .QB (line1405), .D(g24343), .CK(clk));
DFFX1 gate1406(.Q (g3416), .QB (line1406), .D(g25666), .CK(clk));
DFFX1 gate1407(.Q (g5260), .QB (line1407), .D(g30473), .CK(clk));
DFFX1 gate1408(.Q (g1521), .QB (line1408), .D(g24252), .CK(clk));
DFFX1 gate1409(.Q (g3522), .QB (line1409), .D(g33028), .CK(clk));
DFFX1 gate1410(.Q (g3115), .QB (line1410), .D(g29258), .CK(clk));
DFFX1 gate1411(.Q (g3251), .QB (line1411), .D(g30407), .CK(clk));
DFFX1 gate1412(.Q (g1), .QB (line1412), .D(g26958), .CK(clk));
DFFX1 gate1413(.Q (g4628), .QB (line1413), .D(g34457), .CK(clk));
DFFX1 gate1414(.Q (g1996), .QB (line1414), .D(g33568), .CK(clk));
DFFX1 gate1415(.Q (g3447), .QB (line1415), .D(g25663), .CK(clk));
DFFX1 gate1416(.Q (g4515), .QB (line1416), .D(g26964), .CK(clk));
DFFX1 gate1417(.Q (g4204), .QB (line1417), .D(g4200), .CK(clk));
DFFX1 gate1418(.Q (g4300), .QB (line1418), .D(g34735), .CK(clk));
DFFX1 gate1419(.Q (g1724), .QB (line1419), .D(g30352), .CK(clk));
DFFX1 gate1420(.Q (g1379), .QB (line1420), .D(g33543), .CK(clk));
DFFX1 gate1421(.Q (g3654), .QB (line1421), .D(g24271), .CK(clk));
DFFX1 gate1422(.Q (g12), .QB (line1422), .D(g30326), .CK(clk));
DFFX1 gate1423(.Q (g1878), .QB (line1423), .D(g33981), .CK(clk));
DFFX1 gate1424(.Q (g5619), .QB (line1424), .D(g30500), .CK(clk));
DFFX1 gate1425(.Q (g71), .QB (line1425), .D(g34786), .CK(clk));
DFFX1 gate1426(.Q (g59), .QB (line1426), .D(g29277), .CK(clk));
INVX1 gate1427(.O (I28349), .I (g28367));
INVX1 gate1428(.O (g19408), .I (g16066));
INVX1 gate1429(.O (I21294), .I (g18274));
INVX1 gate1430(.O (g13297), .I (g10831));
INVX1 gate1431(.O (g19635), .I (g16349));
INVX1 gate1432(.O (g32394), .I (g30601));
INVX1 gate1433(.O (I19778), .I (g17781));
INVX1 gate1434(.O (g9900), .I (g6));
INVX1 gate1435(.O (g11889), .I (g9954));
INVX1 gate1436(.O (g13103), .I (g10905));
INVX1 gate1437(.O (g17470), .I (g14454));
INVX1 gate1438(.O (g23499), .I (g20785));
INVX1 gate1439(.O (g6895), .I (g3288));
INVX1 gate1440(.O (g9797), .I (g5441));
INVX1 gate1441(.O (g31804), .I (g29385));
INVX1 gate1442(.O (g6837), .I (g968));
INVX1 gate1443(.O (I15824), .I (g1116));
INVX1 gate1444(.O (g20066), .I (g17433));
INVX1 gate1445(.O (g33804), .I (g33250));
INVX1 gate1446(.O (g20231), .I (g17821));
INVX1 gate1447(.O (I19786), .I (g17844));
INVX1 gate1448(.O (g24066), .I (g21127));
INVX1 gate1449(.O (g11888), .I (g10160));
INVX1 gate1450(.O (g9510), .I (g5835));
INVX1 gate1451(.O (I22692), .I (g21308));
INVX1 gate1452(.O (g12884), .I (g10392));
INVX1 gate1453(.O (g22494), .I (g19801));
INVX1 gate1454(.O (g9245), .I (I13031));
INVX1 gate1455(.O (g8925), .I (I12910));
INVX1 gate1456(.O (g34248), .I (I32243));
INVX1 gate1457(.O (g10289), .I (g1319));
INVX1 gate1458(.O (g11181), .I (g8134));
INVX1 gate1459(.O (I20116), .I (g15737));
INVX1 gate1460(.O (g7888), .I (g1536));
INVX1 gate1461(.O (g9291), .I (g3021));
INVX1 gate1462(.O (g28559), .I (g27700));
INVX1 gate1463(.O (g21056), .I (g15426));
INVX1 gate1464(.O (I33246), .I (g34970));
INVX1 gate1465(.O (g10288), .I (I13718));
INVX1 gate1466(.O (g8224), .I (g3774));
INVX1 gate1467(.O (g21611), .I (I21210));
INVX1 gate1468(.O (g16718), .I (I17932));
INVX1 gate1469(.O (g21722), .I (I21285));
INVX1 gate1470(.O (I12530), .I (g4815));
INVX1 gate1471(.O (g16521), .I (g13543));
INVX1 gate1472(.O (I22400), .I (g19620));
INVX1 gate1473(.O (g23611), .I (g18833));
INVX1 gate1474(.O (g10571), .I (g10233));
INVX1 gate1475(.O (g17467), .I (g14339));
INVX1 gate1476(.O (g17494), .I (g14339));
INVX1 gate1477(.O (g10308), .I (g4459));
INVX1 gate1478(.O (g27015), .I (g26869));
INVX1 gate1479(.O (g23988), .I (g19277));
INVX1 gate1480(.O (g23924), .I (g18997));
INVX1 gate1481(.O (g12217), .I (I15070));
INVX1 gate1482(.O (g14571), .I (I16688));
INVX1 gate1483(.O (g32318), .I (g31596));
INVX1 gate1484(.O (g32446), .I (g31596));
INVX1 gate1485(.O (g14308), .I (I16471));
INVX1 gate1486(.O (I24041), .I (g22182));
INVX1 gate1487(.O (I14935), .I (g9902));
INVX1 gate1488(.O (g34778), .I (I32976));
INVX1 gate1489(.O (g20511), .I (g17929));
INVX1 gate1490(.O (g26672), .I (g25275));
INVX1 gate1491(.O (g11931), .I (I14749));
INVX1 gate1492(.O (g20763), .I (I20816));
INVX1 gate1493(.O (g23432), .I (g21514));
INVX1 gate1494(.O (I18165), .I (g13177));
INVX1 gate1495(.O (I18523), .I (g14443));
INVX1 gate1496(.O (g21271), .I (I21002));
INVX1 gate1497(.O (I31776), .I (g33204));
INVX1 gate1498(.O (g23271), .I (g20785));
INVX1 gate1499(.O (g22155), .I (g19074));
INVX1 gate1500(.O (I22539), .I (g19606));
INVX1 gate1501(.O (I32231), .I (g34123));
INVX1 gate1502(.O (g34786), .I (I32988));
INVX1 gate1503(.O (g9259), .I (g5176));
INVX1 gate1504(.O (I15190), .I (g6005));
INVX1 gate1505(.O (g17782), .I (I18788));
INVX1 gate1506(.O (g8277), .I (I12483));
INVX1 gate1507(.O (g9819), .I (g92));
INVX1 gate1508(.O (I16969), .I (g13943));
INVX1 gate1509(.O (g32540), .I (g30614));
INVX1 gate1510(.O (g25027), .I (I24191));
INVX1 gate1511(.O (g19711), .I (g17062));
INVX1 gate1512(.O (g22170), .I (g19210));
INVX1 gate1513(.O (g13190), .I (g10939));
INVX1 gate1514(.O (g7297), .I (g6069));
INVX1 gate1515(.O (g17419), .I (g14965));
INVX1 gate1516(.O (g20660), .I (g17873));
INVX1 gate1517(.O (g16861), .I (I18051));
INVX1 gate1518(.O (g21461), .I (g15348));
INVX1 gate1519(.O (g10816), .I (I14054));
INVX1 gate1520(.O (g28713), .I (g27907));
INVX1 gate1521(.O (g15755), .I (g13134));
INVX1 gate1522(.O (g23461), .I (g18833));
INVX1 gate1523(.O (I24237), .I (g23823));
INVX1 gate1524(.O (g34945), .I (g34933));
INVX1 gate1525(.O (g8789), .I (I12779));
INVX1 gate1526(.O (g31833), .I (g29385));
INVX1 gate1527(.O (I18006), .I (g13638));
INVX1 gate1528(.O (I20035), .I (g15706));
INVX1 gate1529(.O (I17207), .I (g13835));
INVX1 gate1530(.O (g30999), .I (g29722));
INVX1 gate1531(.O (g25249), .I (g22228));
INVX1 gate1532(.O (g9488), .I (g1878));
INVX1 gate1533(.O (g19537), .I (g15938));
INVX1 gate1534(.O (g17155), .I (I18205));
INVX1 gate1535(.O (I16855), .I (g10473));
INVX1 gate1536(.O (g15563), .I (I17140));
INVX1 gate1537(.O (g23031), .I (g19801));
INVX1 gate1538(.O (g30090), .I (g29134));
INVX1 gate1539(.O (g30998), .I (g29719));
INVX1 gate1540(.O (g25248), .I (g22228));
INVX1 gate1541(.O (g23650), .I (g20653));
INVX1 gate1542(.O (g7138), .I (g5360));
INVX1 gate1543(.O (g16099), .I (g13437));
INVX1 gate1544(.O (g34998), .I (g34981));
INVX1 gate1545(.O (g23887), .I (g18997));
INVX1 gate1546(.O (g25552), .I (g22594));
INVX1 gate1547(.O (g20916), .I (g18008));
INVX1 gate1548(.O (g27084), .I (g26673));
INVX1 gate1549(.O (g30182), .I (I28419));
INVX1 gate1550(.O (g7963), .I (g4146));
INVX1 gate1551(.O (g10374), .I (g6903));
INVX1 gate1552(.O (I32763), .I (g34511));
INVX1 gate1553(.O (g19606), .I (g17614));
INVX1 gate1554(.O (g19492), .I (g16349));
INVX1 gate1555(.O (g22167), .I (g19074));
INVX1 gate1556(.O (g22194), .I (I21776));
INVX1 gate1557(.O (g7109), .I (g5011));
INVX1 gate1558(.O (g7791), .I (I12199));
INVX1 gate1559(.O (g34672), .I (I32800));
INVX1 gate1560(.O (g16777), .I (I18003));
INVX1 gate1561(.O (g20550), .I (g15864));
INVX1 gate1562(.O (g23529), .I (g20558));
INVX1 gate1563(.O (g6854), .I (g2685));
INVX1 gate1564(.O (g18930), .I (g15789));
INVX1 gate1565(.O (g13024), .I (g11900));
INVX1 gate1566(.O (g32902), .I (g30673));
INVX1 gate1567(.O (g6941), .I (g3990));
INVX1 gate1568(.O (g12110), .I (I14970));
INVX1 gate1569(.O (g32957), .I (g31672));
INVX1 gate1570(.O (g9951), .I (g6133));
INVX1 gate1571(.O (g32377), .I (g30984));
INVX1 gate1572(.O (g12922), .I (g12297));
INVX1 gate1573(.O (g23528), .I (g18833));
INVX1 gate1574(.O (g12321), .I (g9637));
INVX1 gate1575(.O (g28678), .I (g27800));
INVX1 gate1576(.O (g32739), .I (g30735));
INVX1 gate1577(.O (g21393), .I (g17264));
INVX1 gate1578(.O (g23843), .I (g19147));
INVX1 gate1579(.O (g26026), .I (I25105));
INVX1 gate1580(.O (g25081), .I (g22342));
INVX1 gate1581(.O (g20085), .I (g16187));
INVX1 gate1582(.O (g23393), .I (g20739));
INVX1 gate1583(.O (g19750), .I (g16326));
INVX1 gate1584(.O (g30331), .I (I28594));
INVX1 gate1585(.O (g24076), .I (g19984));
INVX1 gate1586(.O (g24085), .I (g20857));
INVX1 gate1587(.O (g17589), .I (g14981));
INVX1 gate1588(.O (g20596), .I (I20690));
INVX1 gate1589(.O (g34932), .I (g34914));
INVX1 gate1590(.O (g23764), .I (g21308));
INVX1 gate1591(.O (g25786), .I (g24518));
INVX1 gate1592(.O (I25869), .I (g25851));
INVX1 gate1593(.O (g32738), .I (g31376));
INVX1 gate1594(.O (g32562), .I (g30673));
INVX1 gate1595(.O (g32645), .I (g30825));
INVX1 gate1596(.O (g14669), .I (g12301));
INVX1 gate1597(.O (g20054), .I (g17328));
INVX1 gate1598(.O (I26337), .I (g26835));
INVX1 gate1599(.O (g24054), .I (g19919));
INVX1 gate1600(.O (I20130), .I (g15748));
INVX1 gate1601(.O (g17588), .I (g14782));
INVX1 gate1602(.O (g17524), .I (g14933));
INVX1 gate1603(.O (I18600), .I (g5335));
INVX1 gate1604(.O (g23869), .I (g19277));
INVX1 gate1605(.O (g32699), .I (g31528));
INVX1 gate1606(.O (g10392), .I (g6989));
INVX1 gate1607(.O (I28576), .I (g28431));
INVX1 gate1608(.O (I28585), .I (g30217));
INVX1 gate1609(.O (I15987), .I (g12381));
INVX1 gate1610(.O (g14668), .I (g12450));
INVX1 gate1611(.O (g25356), .I (g22763));
INVX1 gate1612(.O (g24431), .I (g22722));
INVX1 gate1613(.O (g29725), .I (g28349));
INVX1 gate1614(.O (I15250), .I (g9152));
INVX1 gate1615(.O (g28294), .I (g27295));
INVX1 gate1616(.O (g8945), .I (g608));
INVX1 gate1617(.O (g10489), .I (g9259));
INVX1 gate1618(.O (g11987), .I (I14833));
INVX1 gate1619(.O (g13625), .I (g10971));
INVX1 gate1620(.O (I25161), .I (g24920));
INVX1 gate1621(.O (g17477), .I (g14848));
INVX1 gate1622(.O (g23868), .I (g19277));
INVX1 gate1623(.O (g32698), .I (g30614));
INVX1 gate1624(.O (g31812), .I (g29385));
INVX1 gate1625(.O (g11250), .I (g7502));
INVX1 gate1626(.O (g25380), .I (g23776));
INVX1 gate1627(.O (I32550), .I (g34398));
INVX1 gate1628(.O (g7957), .I (g1252));
INVX1 gate1629(.O (g13250), .I (I15811));
INVX1 gate1630(.O (g20269), .I (g15844));
INVX1 gate1631(.O (g34505), .I (g34409));
INVX1 gate1632(.O (g7049), .I (g5853));
INVX1 gate1633(.O (g20773), .I (I20830));
INVX1 gate1634(.O (g25090), .I (g23630));
INVX1 gate1635(.O (g6958), .I (g4372));
INVX1 gate1636(.O (g20268), .I (g18008));
INVX1 gate1637(.O (g14424), .I (g11136));
INVX1 gate1638(.O (g34717), .I (I32881));
INVX1 gate1639(.O (g12417), .I (g7175));
INVX1 gate1640(.O (g25182), .I (g22763));
INVX1 gate1641(.O (g12936), .I (g12601));
INVX1 gate1642(.O (g20655), .I (I20753));
INVX1 gate1643(.O (g8340), .I (g3050));
INVX1 gate1644(.O (g13943), .I (I16231));
INVX1 gate1645(.O (g21225), .I (g17428));
INVX1 gate1646(.O (g24156), .I (I23312));
INVX1 gate1647(.O (g23259), .I (g21070));
INVX1 gate1648(.O (g24655), .I (g23067));
INVX1 gate1649(.O (I12109), .I (g749));
INVX1 gate1650(.O (I18063), .I (g14357));
INVX1 gate1651(.O (g7715), .I (g1178));
INVX1 gate1652(.O (g29744), .I (g28431));
INVX1 gate1653(.O (g8478), .I (g3103));
INVX1 gate1654(.O (g20180), .I (g17533));
INVX1 gate1655(.O (g17616), .I (g14309));
INVX1 gate1656(.O (g20670), .I (g15426));
INVX1 gate1657(.O (I29447), .I (g30729));
INVX1 gate1658(.O (g10830), .I (g10087));
INVX1 gate1659(.O (I32243), .I (g34134));
INVX1 gate1660(.O (g22305), .I (g19801));
INVX1 gate1661(.O (g24180), .I (I23384));
INVX1 gate1662(.O (g32632), .I (g31070));
INVX1 gate1663(.O (g31795), .I (I29371));
INVX1 gate1664(.O (g9594), .I (g2307));
INVX1 gate1665(.O (g6829), .I (g1319));
INVX1 gate1666(.O (g7498), .I (g6675));
INVX1 gate1667(.O (g23258), .I (g20924));
INVX1 gate1668(.O (g26811), .I (g25206));
INVX1 gate1669(.O (I16590), .I (g11966));
INVX1 gate1670(.O (g10544), .I (I13906));
INVX1 gate1671(.O (g15573), .I (I17154));
INVX1 gate1672(.O (I27492), .I (g27511));
INVX1 gate1673(.O (g9806), .I (g5782));
INVX1 gate1674(.O (g14544), .I (I16663));
INVX1 gate1675(.O (I14653), .I (g9417));
INVX1 gate1676(.O (I33044), .I (g34775));
INVX1 gate1677(.O (I16741), .I (g5677));
INVX1 gate1678(.O (g25513), .I (g23870));
INVX1 gate1679(.O (g32661), .I (g31070));
INVX1 gate1680(.O (g20993), .I (g15615));
INVX1 gate1681(.O (g32547), .I (g30614));
INVX1 gate1682(.O (g32895), .I (g30673));
INVX1 gate1683(.O (g8876), .I (I12855));
INVX1 gate1684(.O (g24839), .I (g23436));
INVX1 gate1685(.O (g23244), .I (I22343));
INVX1 gate1686(.O (g24993), .I (g22384));
INVX1 gate1687(.O (g22177), .I (g19074));
INVX1 gate1688(.O (g16162), .I (g13437));
INVX1 gate1689(.O (g11855), .I (I14671));
INVX1 gate1690(.O (g20667), .I (g15224));
INVX1 gate1691(.O (g17466), .I (g12983));
INVX1 gate1692(.O (g9887), .I (g5802));
INVX1 gate1693(.O (g6974), .I (I11746));
INVX1 gate1694(.O (g24667), .I (g23112));
INVX1 gate1695(.O (g9934), .I (g5849));
INVX1 gate1696(.O (g21069), .I (g15277));
INVX1 gate1697(.O (g25505), .I (g22228));
INVX1 gate1698(.O (g34433), .I (I32470));
INVX1 gate1699(.O (g34387), .I (g34188));
INVX1 gate1700(.O (g10042), .I (g2671));
INVX1 gate1701(.O (g24131), .I (g21209));
INVX1 gate1702(.O (g32481), .I (g31194));
INVX1 gate1703(.O (g14705), .I (I16803));
INVX1 gate1704(.O (I13321), .I (g6486));
INVX1 gate1705(.O (g18975), .I (g15938));
INVX1 gate1706(.O (g19553), .I (g16782));
INVX1 gate1707(.O (g19862), .I (I20233));
INVX1 gate1708(.O (g30097), .I (g29118));
INVX1 gate1709(.O (g8915), .I (I12884));
INVX1 gate1710(.O (g16629), .I (g13990));
INVX1 gate1711(.O (I16150), .I (g10430));
INVX1 gate1712(.O (g21657), .I (g17657));
INVX1 gate1713(.O (g16472), .I (g14098));
INVX1 gate1714(.O (I20781), .I (g17155));
INVX1 gate1715(.O (g21068), .I (g15277));
INVX1 gate1716(.O (g14255), .I (g12381));
INVX1 gate1717(.O (I21477), .I (g18695));
INVX1 gate1718(.O (g14189), .I (I16391));
INVX1 gate1719(.O (g32551), .I (g30735));
INVX1 gate1720(.O (g32572), .I (g30735));
INVX1 gate1721(.O (g23375), .I (g20924));
INVX1 gate1722(.O (I24781), .I (g24264));
INVX1 gate1723(.O (I33146), .I (g34903));
INVX1 gate1724(.O (g7162), .I (g4521));
INVX1 gate1725(.O (g25212), .I (g22763));
INVX1 gate1726(.O (g7268), .I (g1636));
INVX1 gate1727(.O (I11740), .I (g4519));
INVX1 gate1728(.O (g7362), .I (g1906));
INVX1 gate1729(.O (g12909), .I (g10412));
INVX1 gate1730(.O (g9433), .I (g5148));
INVX1 gate1731(.O (g26850), .I (I25576));
INVX1 gate1732(.O (g12543), .I (g9417));
INVX1 gate1733(.O (g17642), .I (g14691));
INVX1 gate1734(.O (g20502), .I (g15373));
INVX1 gate1735(.O (g10678), .I (I13990));
INVX1 gate1736(.O (I22725), .I (g21250));
INVX1 gate1737(.O (I13740), .I (g85));
INVX1 gate1738(.O (g23879), .I (g19210));
INVX1 gate1739(.O (g20557), .I (I20647));
INVX1 gate1740(.O (g23970), .I (g19277));
INVX1 gate1741(.O (g34343), .I (g34089));
INVX1 gate1742(.O (g20210), .I (g16897));
INVX1 gate1743(.O (I22114), .I (g19935));
INVX1 gate1744(.O (g12908), .I (g10414));
INVX1 gate1745(.O (g20618), .I (g15277));
INVX1 gate1746(.O (g11867), .I (I14679));
INVX1 gate1747(.O (g11894), .I (I14702));
INVX1 gate1748(.O (I11685), .I (g117));
INVX1 gate1749(.O (g8310), .I (g2051));
INVX1 gate1750(.O (g23878), .I (g19147));
INVX1 gate1751(.O (g21337), .I (g15758));
INVX1 gate1752(.O (g20443), .I (g15171));
INVX1 gate1753(.O (g10383), .I (g6978));
INVX1 gate1754(.O (g23337), .I (g20924));
INVX1 gate1755(.O (g19757), .I (g17224));
INVX1 gate1756(.O (g9496), .I (g3303));
INVX1 gate1757(.O (g14383), .I (I16535));
INVX1 gate1758(.O (g17733), .I (g14238));
INVX1 gate1759(.O (I16526), .I (g10430));
INVX1 gate1760(.O (g8663), .I (g3343));
INVX1 gate1761(.O (g10030), .I (g116));
INVX1 gate1762(.O (g23886), .I (g21468));
INVX1 gate1763(.O (I18614), .I (g6315));
INVX1 gate1764(.O (g32490), .I (g30673));
INVX1 gate1765(.O (g10093), .I (g5703));
INVX1 gate1766(.O (g18884), .I (g15938));
INVX1 gate1767(.O (g27242), .I (g26183));
INVX1 gate1768(.O (I14576), .I (g8791));
INVX1 gate1769(.O (g11714), .I (g8107));
INVX1 gate1770(.O (g22166), .I (g18997));
INVX1 gate1771(.O (g11450), .I (I14455));
INVX1 gate1772(.O (I17114), .I (g14358));
INVX1 gate1773(.O (I27192), .I (g27662));
INVX1 gate1774(.O (g23792), .I (g19074));
INVX1 gate1775(.O (g23967), .I (g19210));
INVX1 gate1776(.O (g23994), .I (g19277));
INVX1 gate1777(.O (g32784), .I (g31672));
INVX1 gate1778(.O (g9891), .I (g6173));
INVX1 gate1779(.O (I18320), .I (g13605));
INVX1 gate1780(.O (g28037), .I (g26365));
INVX1 gate1781(.O (g8002), .I (g1389));
INVX1 gate1782(.O (g9337), .I (g1608));
INVX1 gate1783(.O (g9913), .I (g2403));
INVX1 gate1784(.O (g32956), .I (g30825));
INVX1 gate1785(.O (I21285), .I (g18215));
INVX1 gate1786(.O (g11819), .I (g7717));
INVX1 gate1787(.O (g11910), .I (g10185));
INVX1 gate1788(.O (g14065), .I (g11048));
INVX1 gate1789(.O (g7086), .I (g4826));
INVX1 gate1790(.O (g13707), .I (g11360));
INVX1 gate1791(.O (g31829), .I (g29385));
INVX1 gate1792(.O (g32889), .I (g31376));
INVX1 gate1793(.O (g11202), .I (I14267));
INVX1 gate1794(.O (g8236), .I (g4812));
INVX1 gate1795(.O (g33920), .I (I31786));
INVX1 gate1796(.O (I21254), .I (g16540));
INVX1 gate1797(.O (g24039), .I (g21256));
INVX1 gate1798(.O (g25620), .I (I24759));
INVX1 gate1799(.O (g21425), .I (g15509));
INVX1 gate1800(.O (g29221), .I (I27579));
INVX1 gate1801(.O (I17744), .I (g14912));
INVX1 gate1802(.O (g23459), .I (g21611));
INVX1 gate1803(.O (I16917), .I (g10582));
INVX1 gate1804(.O (g20038), .I (g17328));
INVX1 gate1805(.O (g23425), .I (g20751));
INVX1 gate1806(.O (g31828), .I (g29385));
INVX1 gate1807(.O (g32888), .I (g30673));
INVX1 gate1808(.O (I15070), .I (g10108));
INVX1 gate1809(.O (g25097), .I (g22342));
INVX1 gate1810(.O (g32824), .I (g31376));
INVX1 gate1811(.O (g10219), .I (g2697));
INVX1 gate1812(.O (g13055), .I (I15682));
INVX1 gate1813(.O (g9807), .I (g5712));
INVX1 gate1814(.O (I30901), .I (g32407));
INVX1 gate1815(.O (g19673), .I (g16931));
INVX1 gate1816(.O (g24038), .I (g21193));
INVX1 gate1817(.O (g14219), .I (g12381));
INVX1 gate1818(.O (g19397), .I (g16449));
INVX1 gate1819(.O (g21458), .I (g15758));
INVX1 gate1820(.O (g6849), .I (g2551));
INVX1 gate1821(.O (I15590), .I (g11988));
INVX1 gate1822(.O (g28155), .I (I26664));
INVX1 gate1823(.O (I13762), .I (g6755));
INVX1 gate1824(.O (g13070), .I (g11984));
INVX1 gate1825(.O (g23458), .I (I22583));
INVX1 gate1826(.O (g32671), .I (g31528));
INVX1 gate1827(.O (I21036), .I (g17221));
INVX1 gate1828(.O (g34229), .I (g33936));
INVX1 gate1829(.O (g10218), .I (g2527));
INVX1 gate1830(.O (I18034), .I (g13680));
INVX1 gate1831(.O (g16172), .I (g13584));
INVX1 gate1832(.O (g20601), .I (g17433));
INVX1 gate1833(.O (g21010), .I (g15634));
INVX1 gate1834(.O (g11986), .I (I14830));
INVX1 gate1835(.O (g7470), .I (g5623));
INVX1 gate1836(.O (I12483), .I (g3096));
INVX1 gate1837(.O (g17476), .I (g14665));
INVX1 gate1838(.O (g17485), .I (I18408));
INVX1 gate1839(.O (I16077), .I (g10430));
INVX1 gate1840(.O (I14745), .I (g10029));
INVX1 gate1841(.O (g11741), .I (g10033));
INVX1 gate1842(.O (g22907), .I (g20453));
INVX1 gate1843(.O (g23545), .I (g21562));
INVX1 gate1844(.O (g23444), .I (I22561));
INVX1 gate1845(.O (g25369), .I (g22228));
INVX1 gate1846(.O (g32931), .I (g30937));
INVX1 gate1847(.O (g33682), .I (I31515));
INVX1 gate1848(.O (g6900), .I (g3440));
INVX1 gate1849(.O (g19634), .I (g16349));
INVX1 gate1850(.O (g19872), .I (g17015));
INVX1 gate1851(.O (g34716), .I (I32878));
INVX1 gate1852(.O (I20542), .I (g16508));
INVX1 gate1853(.O (I25598), .I (g25424));
INVX1 gate1854(.O (g8928), .I (g4340));
INVX1 gate1855(.O (g29812), .I (g28381));
INVX1 gate1856(.O (I28241), .I (g28709));
INVX1 gate1857(.O (g12841), .I (g10357));
INVX1 gate1858(.O (g22594), .I (I21934));
INVX1 gate1859(.O (I16688), .I (g10981));
INVX1 gate1860(.O (g9815), .I (g6098));
INVX1 gate1861(.O (g8064), .I (g3376));
INVX1 gate1862(.O (I18408), .I (g13017));
INVX1 gate1863(.O (I20913), .I (g16964));
INVX1 gate1864(.O (g23086), .I (g20283));
INVX1 gate1865(.O (I32815), .I (g34470));
INVX1 gate1866(.O (g30310), .I (g28830));
INVX1 gate1867(.O (g8899), .I (g807));
INVX1 gate1868(.O (g11735), .I (g8534));
INVX1 gate1869(.O (g29371), .I (I27735));
INVX1 gate1870(.O (I11908), .I (g4449));
INVX1 gate1871(.O (g9692), .I (g1756));
INVX1 gate1872(.O (g13877), .I (g11350));
INVX1 gate1873(.O (I32601), .I (g34319));
INVX1 gate1874(.O (g8785), .I (I12767));
INVX1 gate1875(.O (g24169), .I (I23351));
INVX1 gate1876(.O (g24791), .I (g23850));
INVX1 gate1877(.O (g9497), .I (I13166));
INVX1 gate1878(.O (I16102), .I (g10430));
INVX1 gate1879(.O (g26681), .I (g25396));
INVX1 gate1880(.O (g20168), .I (g17533));
INVX1 gate1881(.O (g9154), .I (I12994));
INVX1 gate1882(.O (g25133), .I (g23733));
INVX1 gate1883(.O (g34925), .I (I33167));
INVX1 gate1884(.O (I26309), .I (g26825));
INVX1 gate1885(.O (g9354), .I (g2719));
INVX1 gate1886(.O (g27014), .I (g25888));
INVX1 gate1887(.O (I27564), .I (g28166));
INVX1 gate1888(.O (g24168), .I (I23348));
INVX1 gate1889(.O (g23322), .I (I22425));
INVX1 gate1890(.O (g32546), .I (g31170));
INVX1 gate1891(.O (g9960), .I (g6474));
INVX1 gate1892(.O (g22519), .I (g19801));
INVX1 gate1893(.O (g22176), .I (g18997));
INVX1 gate1894(.O (g14201), .I (I16401));
INVX1 gate1895(.O (g26802), .I (I25514));
INVX1 gate1896(.O (g28119), .I (g27008));
INVX1 gate1897(.O (g12835), .I (g10352));
INVX1 gate1898(.O (g7635), .I (g1002));
INVX1 gate1899(.O (g14277), .I (I16455));
INVX1 gate1900(.O (g20666), .I (g15224));
INVX1 gate1901(.O (g13018), .I (I15636));
INVX1 gate1902(.O (I16231), .I (g10520));
INVX1 gate1903(.O (g32024), .I (I29582));
INVX1 gate1904(.O (g25228), .I (g23828));
INVX1 gate1905(.O (I19802), .I (g15727));
INVX1 gate1906(.O (g19574), .I (g16826));
INVX1 gate1907(.O (g7766), .I (I12189));
INVX1 gate1908(.O (g19452), .I (g16326));
INVX1 gate1909(.O (g6819), .I (g1046));
INVX1 gate1910(.O (g16540), .I (I17744));
INVX1 gate1911(.O (I19857), .I (g16640));
INVX1 gate1912(.O (g22154), .I (g19074));
INVX1 gate1913(.O (g7087), .I (g6336));
INVX1 gate1914(.O (I33297), .I (g35000));
INVX1 gate1915(.O (g25011), .I (g22763));
INVX1 gate1916(.O (g32860), .I (g30673));
INVX1 gate1917(.O (I18891), .I (g16676));
INVX1 gate1918(.O (g7487), .I (g1259));
INVX1 gate1919(.O (I33103), .I (g34846));
INVX1 gate1920(.O (g8237), .I (g255));
INVX1 gate1921(.O (g18953), .I (g16077));
INVX1 gate1922(.O (I14761), .I (g7753));
INVX1 gate1923(.O (g19912), .I (g17328));
INVX1 gate1924(.O (g17519), .I (I18460));
INVX1 gate1925(.O (g21561), .I (g15595));
INVX1 gate1926(.O (I12183), .I (g2719));
INVX1 gate1927(.O (g21656), .I (g17700));
INVX1 gate1928(.O (g6923), .I (g3791));
INVX1 gate1929(.O (g26765), .I (g25309));
INVX1 gate1930(.O (I25680), .I (g25641));
INVX1 gate1931(.O (g22935), .I (g20283));
INVX1 gate1932(.O (g17092), .I (g14011));
INVX1 gate1933(.O (g34944), .I (g34932));
INVX1 gate1934(.O (g10037), .I (g1848));
INVX1 gate1935(.O (I32791), .I (g34578));
INVX1 gate1936(.O (g32497), .I (g30673));
INVX1 gate1937(.O (g21295), .I (g17533));
INVX1 gate1938(.O (g23353), .I (g20924));
INVX1 gate1939(.O (g29507), .I (g28353));
INVX1 gate1940(.O (I32884), .I (g34690));
INVX1 gate1941(.O (g8844), .I (I12826));
INVX1 gate1942(.O (g11402), .I (g7594));
INVX1 gate1943(.O (g17518), .I (g14918));
INVX1 gate1944(.O (g26549), .I (I25391));
INVX1 gate1945(.O (g17154), .I (g14348));
INVX1 gate1946(.O (g22883), .I (g20391));
INVX1 gate1947(.O (g20556), .I (g15483));
INVX1 gate1948(.O (g23823), .I (I22989));
INVX1 gate1949(.O (g17637), .I (g12933));
INVX1 gate1950(.O (g20580), .I (g17328));
INVX1 gate1951(.O (g26548), .I (g25255));
INVX1 gate1952(.O (g10419), .I (g8821));
INVX1 gate1953(.O (g11866), .I (g9883));
INVX1 gate1954(.O (g11917), .I (I14727));
INVX1 gate1955(.O (g32700), .I (g31579));
INVX1 gate1956(.O (I26687), .I (g27880));
INVX1 gate1957(.O (g32659), .I (g30735));
INVX1 gate1958(.O (g21336), .I (g17367));
INVX1 gate1959(.O (g32625), .I (g31070));
INVX1 gate1960(.O (g10352), .I (g6804));
INVX1 gate1961(.O (g23336), .I (g20924));
INVX1 gate1962(.O (I32479), .I (g34302));
INVX1 gate1963(.O (g19592), .I (I20035));
INVX1 gate1964(.O (g34429), .I (I32458));
INVX1 gate1965(.O (g10155), .I (g2643));
INVX1 gate1966(.O (g10418), .I (g8818));
INVX1 gate1967(.O (g12041), .I (I14905));
INVX1 gate1968(.O (g32658), .I (g31579));
INVX1 gate1969(.O (g19780), .I (g16449));
INVX1 gate1970(.O (g16739), .I (g13223));
INVX1 gate1971(.O (g12430), .I (I15250));
INVX1 gate1972(.O (I16660), .I (g10981));
INVX1 gate1973(.O (g34428), .I (I32455));
INVX1 gate1974(.O (I21074), .I (g17766));
INVX1 gate1975(.O (g23966), .I (g19210));
INVX1 gate1976(.O (g22215), .I (g19277));
INVX1 gate1977(.O (g28036), .I (g26365));
INVX1 gate1978(.O (g27237), .I (g26162));
INVX1 gate1979(.O (g32943), .I (g31710));
INVX1 gate1980(.O (g20110), .I (g16897));
INVX1 gate1981(.O (g11706), .I (I14579));
INVX1 gate1982(.O (g24084), .I (g20720));
INVX1 gate1983(.O (g16738), .I (I17956));
INVX1 gate1984(.O (g9761), .I (g2445));
INVX1 gate1985(.O (g13706), .I (g11280));
INVX1 gate1986(.O (g16645), .I (g13756));
INVX1 gate1987(.O (g12465), .I (g7192));
INVX1 gate1988(.O (I11992), .I (g763));
INVX1 gate1989(.O (g24110), .I (g21209));
INVX1 gate1990(.O (g20922), .I (I20891));
INVX1 gate1991(.O (g27983), .I (g26725));
INVX1 gate1992(.O (g20321), .I (g17821));
INVX1 gate1993(.O (g23017), .I (g20453));
INVX1 gate1994(.O (g32644), .I (g30735));
INVX1 gate1995(.O (g33648), .I (I31482));
INVX1 gate1996(.O (I21238), .I (g16540));
INVX1 gate1997(.O (g34690), .I (I32840));
INVX1 gate1998(.O (g6870), .I (g3089));
INVX1 gate1999(.O (g9828), .I (g2024));
INVX1 gate2000(.O (g20179), .I (g17249));
INVX1 gate2001(.O (g34549), .I (I32617));
INVX1 gate2002(.O (g8948), .I (g785));
INVX1 gate2003(.O (g20531), .I (g15907));
INVX1 gate2004(.O (g12983), .I (I15600));
INVX1 gate2005(.O (g24179), .I (I23381));
INVX1 gate2006(.O (g16290), .I (g13260));
INVX1 gate2007(.O (g32969), .I (g30735));
INVX1 gate2008(.O (g13280), .I (I15846));
INVX1 gate2009(.O (g6825), .I (g979));
INVX1 gate2010(.O (g33755), .I (I31610));
INVX1 gate2011(.O (g17501), .I (I18434));
INVX1 gate2012(.O (g7369), .I (g1996));
INVX1 gate2013(.O (g27142), .I (g26105));
INVX1 gate2014(.O (g8955), .I (g1418));
INVX1 gate2015(.O (g20178), .I (g16971));
INVX1 gate2016(.O (g10194), .I (g6741));
INVX1 gate2017(.O (g19396), .I (g16431));
INVX1 gate2018(.O (g17577), .I (I18504));
INVX1 gate2019(.O (g13624), .I (g10951));
INVX1 gate2020(.O (I14241), .I (g8356));
INVX1 gate2021(.O (I21941), .I (g18918));
INVX1 gate2022(.O (g24178), .I (I23378));
INVX1 gate2023(.O (g14167), .I (I16371));
INVX1 gate2024(.O (g32968), .I (g31376));
INVX1 gate2025(.O (g19731), .I (g17093));
INVX1 gate2026(.O (g29920), .I (g28824));
INVX1 gate2027(.O (g34504), .I (g34408));
INVX1 gate2028(.O (g29358), .I (I27718));
INVX1 gate2029(.O (g7868), .I (g1099));
INVX1 gate2030(.O (I15102), .I (g5313));
INVX1 gate2031(.O (I26195), .I (g26260));
INVX1 gate2032(.O (I11835), .I (g101));
INVX1 gate2033(.O (I20891), .I (g17700));
INVX1 gate2034(.O (g9746), .I (I13326));
INVX1 gate2035(.O (g20373), .I (g17929));
INVX1 gate2036(.O (g32855), .I (g30825));
INVX1 gate2037(.O (g23289), .I (g20924));
INVX1 gate2038(.O (g24685), .I (g23139));
INVX1 gate2039(.O (g24373), .I (g22908));
INVX1 gate2040(.O (I33024), .I (g34783));
INVX1 gate2041(.O (g8150), .I (g2185));
INVX1 gate2042(.O (g10401), .I (g7041));
INVX1 gate2043(.O (g22906), .I (g20453));
INVX1 gate2044(.O (g20654), .I (I20750));
INVX1 gate2045(.O (I16596), .I (g12640));
INVX1 gate2046(.O (g34317), .I (g34115));
INVX1 gate2047(.O (g8350), .I (g4646));
INVX1 gate2048(.O (g18908), .I (g16100));
INVX1 gate2049(.O (g32870), .I (g31021));
INVX1 gate2050(.O (g7535), .I (g1500));
INVX1 gate2051(.O (g32527), .I (g30673));
INVX1 gate2052(.O (I13007), .I (g65));
INVX1 gate2053(.O (g8038), .I (I12360));
INVX1 gate2054(.O (g10119), .I (g2841));
INVX1 gate2055(.O (I24474), .I (g22546));
INVX1 gate2056(.O (g16632), .I (g14454));
INVX1 gate2057(.O (g21308), .I (g17485));
INVX1 gate2058(.O (g8438), .I (g3100));
INVX1 gate2059(.O (g23571), .I (g18833));
INVX1 gate2060(.O (g28693), .I (g27837));
INVX1 gate2061(.O (g23308), .I (g21024));
INVX1 gate2062(.O (g31794), .I (I29368));
INVX1 gate2063(.O (g6972), .I (I11740));
INVX1 gate2064(.O (g31845), .I (g29385));
INVX1 gate2065(.O (g8009), .I (g3106));
INVX1 gate2066(.O (I31497), .I (g33187));
INVX1 gate2067(.O (g7261), .I (g4449));
INVX1 gate2068(.O (g24417), .I (g22171));
INVX1 gate2069(.O (g33845), .I (I31694));
INVX1 gate2070(.O (g10118), .I (g2541));
INVX1 gate2071(.O (I19775), .I (g17780));
INVX1 gate2072(.O (g9932), .I (g5805));
INVX1 gate2073(.O (g28166), .I (I26687));
INVX1 gate2074(.O (g28009), .I (I26516));
INVX1 gate2075(.O (g16661), .I (g14454));
INVX1 gate2076(.O (I17507), .I (g13416));
INVX1 gate2077(.O (g25549), .I (g22763));
INVX1 gate2078(.O (g13876), .I (g11432));
INVX1 gate2079(.O (g13885), .I (g10862));
INVX1 gate2080(.O (g32503), .I (g31194));
INVX1 gate2081(.O (g23495), .I (I22622));
INVX1 gate2082(.O (I31659), .I (g33219));
INVX1 gate2083(.O (g14749), .I (I16829));
INVX1 gate2084(.O (g32867), .I (g30673));
INVX1 gate2085(.O (g32894), .I (g30614));
INVX1 gate2086(.O (I31625), .I (g33197));
INVX1 gate2087(.O (g14616), .I (I16733));
INVX1 gate2088(.O (g34245), .I (I32234));
INVX1 gate2089(.O (I32953), .I (g34656));
INVX1 gate2090(.O (g8836), .I (g736));
INVX1 gate2091(.O (g30299), .I (g28765));
INVX1 gate2092(.O (g6887), .I (g3333));
INVX1 gate2093(.O (g23816), .I (g21308));
INVX1 gate2094(.O (g25548), .I (g22550));
INVX1 gate2095(.O (g34323), .I (g34105));
INVX1 gate2096(.O (g34299), .I (g34080));
INVX1 gate2097(.O (I32654), .I (g34378));
INVX1 gate2098(.O (g22139), .I (I21722));
INVX1 gate2099(.O (g8918), .I (I12893));
INVX1 gate2100(.O (g24964), .I (I24128));
INVX1 gate2101(.O (g7246), .I (g4446));
INVX1 gate2102(.O (I11746), .I (g4570));
INVX1 gate2103(.O (g26856), .I (I25586));
INVX1 gate2104(.O (g13763), .I (g10971));
INVX1 gate2105(.O (g14276), .I (I16452));
INVX1 gate2106(.O (g31521), .I (I29182));
INVX1 gate2107(.O (I32800), .I (g34582));
INVX1 gate2108(.O (g32581), .I (g31070));
INVX1 gate2109(.O (g32714), .I (g31528));
INVX1 gate2110(.O (g32450), .I (g31591));
INVX1 gate2111(.O (g10053), .I (g6381));
INVX1 gate2112(.O (g23985), .I (g19210));
INVX1 gate2113(.O (g22138), .I (g21370));
INVX1 gate2114(.O (g15739), .I (g13284));
INVX1 gate2115(.O (I26705), .I (g27967));
INVX1 gate2116(.O (g34775), .I (I32967));
INVX1 gate2117(.O (I20750), .I (g16677));
INVX1 gate2118(.O (g20587), .I (g15373));
INVX1 gate2119(.O (g32707), .I (g31579));
INVX1 gate2120(.O (g32819), .I (g30825));
INVX1 gate2121(.O (g9576), .I (g6565));
INVX1 gate2122(.O (g31832), .I (g29385));
INVX1 gate2123(.O (I20982), .I (g16300));
INVX1 gate2124(.O (g23954), .I (I23099));
INVX1 gate2125(.O (g24587), .I (g23112));
INVX1 gate2126(.O (g8229), .I (g3881));
INVX1 gate2127(.O (g9716), .I (g5057));
INVX1 gate2128(.O (I22788), .I (g18940));
INVX1 gate2129(.O (I26679), .I (g27773));
INVX1 gate2130(.O (g12863), .I (g10371));
INVX1 gate2131(.O (g8993), .I (g385));
INVX1 gate2132(.O (g15562), .I (g14943));
INVX1 gate2133(.O (g32818), .I (g30735));
INVX1 gate2134(.O (g10036), .I (g1816));
INVX1 gate2135(.O (g32496), .I (g30614));
INVX1 gate2136(.O (g19787), .I (g17096));
INVX1 gate2137(.O (g16127), .I (g13437));
INVX1 gate2138(.O (g8822), .I (g4975));
INVX1 gate2139(.O (g10177), .I (g1834));
INVX1 gate2140(.O (g20909), .I (g17955));
INVX1 gate2141(.O (g20543), .I (g17955));
INVX1 gate2142(.O (I13684), .I (g128));
INVX1 gate2143(.O (g31861), .I (I29441));
INVX1 gate2144(.O (g9848), .I (g4462));
INVX1 gate2145(.O (g21669), .I (I21230));
INVX1 gate2146(.O (g19357), .I (I19837));
INVX1 gate2147(.O (g17415), .I (g14797));
INVX1 gate2148(.O (g6845), .I (g2126));
INVX1 gate2149(.O (g7502), .I (I11992));
INVX1 gate2150(.O (I15550), .I (g10430));
INVX1 gate2151(.O (g32590), .I (g31154));
INVX1 gate2152(.O (g9699), .I (g2311));
INVX1 gate2153(.O (g9747), .I (I13329));
INVX1 gate2154(.O (g24117), .I (g21209));
INVX1 gate2155(.O (g24000), .I (g19277));
INVX1 gate2156(.O (I33197), .I (g34930));
INVX1 gate2157(.O (g23260), .I (g21070));
INVX1 gate2158(.O (g19743), .I (g17125));
INVX1 gate2159(.O (I14584), .I (g9766));
INVX1 gate2160(.O (g33926), .I (I31796));
INVX1 gate2161(.O (g25245), .I (g22763));
INVX1 gate2162(.O (g34697), .I (g34545));
INVX1 gate2163(.O (g26831), .I (g24836));
INVX1 gate2164(.O (g20569), .I (g15277));
INVX1 gate2165(.O (I20840), .I (g17727));
INVX1 gate2166(.O (g34995), .I (I33285));
INVX1 gate2167(.O (g23842), .I (g19147));
INVX1 gate2168(.O (g32741), .I (g31710));
INVX1 gate2169(.O (g13314), .I (g10893));
INVX1 gate2170(.O (I23348), .I (g23384));
INVX1 gate2171(.O (g25299), .I (g22763));
INVX1 gate2172(.O (g32384), .I (g31666));
INVX1 gate2173(.O (I19831), .I (g16533));
INVX1 gate2174(.O (g33388), .I (g32382));
INVX1 gate2175(.O (I18252), .I (g13177));
INVX1 gate2176(.O (I16502), .I (g10430));
INVX1 gate2177(.O (g20568), .I (g15509));
INVX1 gate2178(.O (g23489), .I (g21468));
INVX1 gate2179(.O (g25533), .I (g22550));
INVX1 gate2180(.O (g13085), .I (I15717));
INVX1 gate2181(.O (g19769), .I (g16987));
INVX1 gate2182(.O (g24568), .I (g22942));
INVX1 gate2183(.O (g20242), .I (g16308));
INVX1 gate2184(.O (g25298), .I (g23760));
INVX1 gate2185(.O (g11721), .I (g10074));
INVX1 gate2186(.O (g7689), .I (I12159));
INVX1 gate2187(.O (g29927), .I (g28861));
INVX1 gate2188(.O (I17121), .I (g14366));
INVX1 gate2189(.O (g34512), .I (g34420));
INVX1 gate2190(.O (g21424), .I (g15426));
INVX1 gate2191(.O (g23559), .I (g21070));
INVX1 gate2192(.O (g13596), .I (g10971));
INVX1 gate2193(.O (g23525), .I (g21562));
INVX1 gate2194(.O (g23488), .I (g21468));
INVX1 gate2195(.O (g28675), .I (g27779));
INVX1 gate2196(.O (g23016), .I (g20453));
INVX1 gate2197(.O (I32909), .I (g34712));
INVX1 gate2198(.O (g7216), .I (g822));
INVX1 gate2199(.O (g11431), .I (g7618));
INVX1 gate2200(.O (g12952), .I (I15572));
INVX1 gate2201(.O (g23558), .I (g20924));
INVX1 gate2202(.O (g13431), .I (I15932));
INVX1 gate2203(.O (g32801), .I (g30937));
INVX1 gate2204(.O (g14630), .I (g12402));
INVX1 gate2205(.O (g32735), .I (g31021));
INVX1 gate2206(.O (g24123), .I (g21143));
INVX1 gate2207(.O (g32877), .I (g30825));
INVX1 gate2208(.O (g7028), .I (I11785));
INVX1 gate2209(.O (I30686), .I (g32381));
INVX1 gate2210(.O (g8895), .I (g599));
INVX1 gate2211(.O (g10166), .I (g6040));
INVX1 gate2212(.O (g17576), .I (g14953));
INVX1 gate2213(.O (g17585), .I (g14974));
INVX1 gate2214(.O (g20772), .I (g15171));
INVX1 gate2215(.O (g9644), .I (g2016));
INVX1 gate2216(.O (g22200), .I (g19277));
INVX1 gate2217(.O (g23893), .I (g19074));
INVX1 gate2218(.O (I15773), .I (g10430));
INVX1 gate2219(.O (g11269), .I (g7516));
INVX1 gate2220(.O (I15942), .I (g12381));
INVX1 gate2221(.O (g14166), .I (g11048));
INVX1 gate2222(.O (g8620), .I (g3065));
INVX1 gate2223(.O (g19881), .I (g15915));
INVX1 gate2224(.O (g8462), .I (g1183));
INVX1 gate2225(.O (g25232), .I (g22228));
INVX1 gate2226(.O (g29491), .I (I27777));
INVX1 gate2227(.O (g7247), .I (g5377));
INVX1 gate2228(.O (g20639), .I (g15224));
INVX1 gate2229(.O (I17173), .I (g13716));
INVX1 gate2230(.O (g16931), .I (I18101));
INVX1 gate2231(.O (I16468), .I (g12760));
INVX1 gate2232(.O (g23544), .I (g21562));
INVX1 gate2233(.O (g23865), .I (g21308));
INVX1 gate2234(.O (I12046), .I (g613));
INVX1 gate2235(.O (g32695), .I (g30735));
INVX1 gate2236(.O (I31581), .I (g33164));
INVX1 gate2237(.O (g11268), .I (g7515));
INVX1 gate2238(.O (g20230), .I (I20499));
INVX1 gate2239(.O (g12790), .I (g7097));
INVX1 gate2240(.O (g17609), .I (g14817));
INVX1 gate2241(.O (g29755), .I (I28002));
INVX1 gate2242(.O (g7564), .I (g336));
INVX1 gate2243(.O (g9152), .I (g2834));
INVX1 gate2244(.O (g20638), .I (g15224));
INVX1 gate2245(.O (I18509), .I (g5623));
INVX1 gate2246(.O (g9818), .I (g6490));
INVX1 gate2247(.O (g13655), .I (g10573));
INVX1 gate2248(.O (g34316), .I (g34093));
INVX1 gate2249(.O (g17200), .I (I18238));
INVX1 gate2250(.O (g32526), .I (g30614));
INVX1 gate2251(.O (g20265), .I (g17821));
INVX1 gate2252(.O (g29981), .I (g28942));
INVX1 gate2253(.O (g6815), .I (g929));
INVX1 gate2254(.O (I12787), .I (g4311));
INVX1 gate2255(.O (g12873), .I (g10380));
INVX1 gate2256(.O (I22028), .I (g20204));
INVX1 gate2257(.O (I29211), .I (g30298));
INVX1 gate2258(.O (g8788), .I (I12776));
INVX1 gate2259(.O (I18872), .I (g13745));
INVX1 gate2260(.O (I23333), .I (g22683));
INVX1 gate2261(.O (g30989), .I (g29672));
INVX1 gate2262(.O (g33766), .I (I31619));
INVX1 gate2263(.O (g19662), .I (g17432));
INVX1 gate2264(.O (g21610), .I (g15615));
INVX1 gate2265(.O (g14454), .I (I16613));
INVX1 gate2266(.O (g23610), .I (g18833));
INVX1 gate2267(.O (g10570), .I (g9021));
INVX1 gate2268(.O (g34989), .I (I33267));
INVX1 gate2269(.O (g8249), .I (g1917));
INVX1 gate2270(.O (g20391), .I (I20562));
INVX1 gate2271(.O (g32457), .I (g30735));
INVX1 gate2272(.O (g21189), .I (g15634));
INVX1 gate2273(.O (g24992), .I (g22417));
INVX1 gate2274(.O (I33070), .I (g34810));
INVX1 gate2275(.O (g20510), .I (g17226));
INVX1 gate2276(.O (g23189), .I (g20060));
INVX1 gate2277(.O (g11930), .I (g9281));
INVX1 gate2278(.O (g12422), .I (I15238));
INVX1 gate2279(.O (g26736), .I (g25349));
INVX1 gate2280(.O (g9186), .I (I13010));
INVX1 gate2281(.O (g17745), .I (g14978));
INVX1 gate2282(.O (g34988), .I (I33264));
INVX1 gate2283(.O (g22973), .I (g20330));
INVX1 gate2284(.O (g34924), .I (I33164));
INVX1 gate2285(.O (g6960), .I (g1));
INVX1 gate2286(.O (g9386), .I (g5727));
INVX1 gate2287(.O (I15667), .I (g12143));
INVX1 gate2288(.O (I32639), .I (g34345));
INVX1 gate2289(.O (g21270), .I (I20999));
INVX1 gate2290(.O (g32866), .I (g30614));
INVX1 gate2291(.O (g32917), .I (g30937));
INVX1 gate2292(.O (g23270), .I (g20785));
INVX1 gate2293(.O (g19482), .I (g16349));
INVX1 gate2294(.O (g21678), .I (g16540));
INVX1 gate2295(.O (g17813), .I (I18813));
INVX1 gate2296(.O (g12834), .I (g10349));
INVX1 gate2297(.O (g20579), .I (g17249));
INVX1 gate2298(.O (g34432), .I (I32467));
INVX1 gate2299(.O (g7308), .I (g1668));
INVX1 gate2300(.O (g11965), .I (I14797));
INVX1 gate2301(.O (g8085), .I (I12382));
INVX1 gate2302(.O (g9599), .I (g3310));
INVX1 gate2303(.O (g10074), .I (g718));
INVX1 gate2304(.O (g19710), .I (g17059));
INVX1 gate2305(.O (g18983), .I (g16077));
INVX1 gate2306(.O (g24579), .I (g23067));
INVX1 gate2307(.O (g34271), .I (g34160));
INVX1 gate2308(.O (g19552), .I (g16856));
INVX1 gate2309(.O (g21460), .I (g15628));
INVX1 gate2310(.O (g21686), .I (g16540));
INVX1 gate2311(.O (g9274), .I (g5857));
INVX1 gate2312(.O (g20578), .I (g15563));
INVX1 gate2313(.O (g26843), .I (I25567));
INVX1 gate2314(.O (g23460), .I (g21611));
INVX1 gate2315(.O (g23939), .I (g19074));
INVX1 gate2316(.O (g21383), .I (g17367));
INVX1 gate2317(.O (g19779), .I (g16431));
INVX1 gate2318(.O (I19843), .I (g16594));
INVX1 gate2319(.O (g9614), .I (g5128));
INVX1 gate2320(.O (I33067), .I (g34812));
INVX1 gate2321(.O (g17674), .I (I18647));
INVX1 gate2322(.O (g12021), .I (g9543));
INVX1 gate2323(.O (g14238), .I (g10823));
INVX1 gate2324(.O (g20586), .I (g15171));
INVX1 gate2325(.O (g23030), .I (g20453));
INVX1 gate2326(.O (g32706), .I (g30673));
INVX1 gate2327(.O (g23938), .I (g18997));
INVX1 gate2328(.O (g32597), .I (g31154));
INVX1 gate2329(.O (I18574), .I (g13075));
INVX1 gate2330(.O (g25316), .I (g22763));
INVX1 gate2331(.O (g8854), .I (g613));
INVX1 gate2332(.O (g21267), .I (g15680));
INVX1 gate2333(.O (g24586), .I (g23067));
INVX1 gate2334(.O (I32391), .I (g34153));
INVX1 gate2335(.O (g23267), .I (g20097));
INVX1 gate2336(.O (g9821), .I (g115));
INVX1 gate2337(.O (I13236), .I (g5452));
INVX1 gate2338(.O (I18205), .I (g14563));
INVX1 gate2339(.O (g34145), .I (I32096));
INVX1 gate2340(.O (I16168), .I (g3321));
INVX1 gate2341(.O (g26869), .I (g24842));
INVX1 gate2342(.O (g32689), .I (g30825));
INVX1 gate2343(.O (g15824), .I (I17324));
INVX1 gate2344(.O (g20442), .I (g15171));
INVX1 gate2345(.O (g10382), .I (g6958));
INVX1 gate2346(.O (I18912), .I (g15050));
INVX1 gate2347(.O (I22240), .I (g20086));
INVX1 gate2348(.O (g32923), .I (g31021));
INVX1 gate2349(.O (g33451), .I (g32132));
INVX1 gate2350(.O (g19786), .I (g17062));
INVX1 gate2351(.O (I14833), .I (g10142));
INVX1 gate2352(.O (g16659), .I (I17857));
INVX1 gate2353(.O (g12614), .I (g9935));
INVX1 gate2354(.O (g22761), .I (g21024));
INVX1 gate2355(.O (g9280), .I (I13054));
INVX1 gate2356(.O (g10519), .I (g9326));
INVX1 gate2357(.O (g34736), .I (I32904));
INVX1 gate2358(.O (g10176), .I (g44));
INVX1 gate2359(.O (I16479), .I (g10430));
INVX1 gate2360(.O (g27320), .I (I26004));
INVX1 gate2361(.O (g16987), .I (I18135));
INVX1 gate2362(.O (g32688), .I (g30735));
INVX1 gate2363(.O (g32624), .I (g30825));
INVX1 gate2364(.O (I23312), .I (g21681));
INVX1 gate2365(.O (g13279), .I (I15843));
INVX1 gate2366(.O (I16217), .I (g3632));
INVX1 gate2367(.O (I21115), .I (g15714));
INVX1 gate2368(.O (g16658), .I (g14157));
INVX1 gate2369(.O (I22604), .I (g21143));
INVX1 gate2370(.O (g10518), .I (g9311));
INVX1 gate2371(.O (g10154), .I (g2547));
INVX1 gate2372(.O (g12905), .I (g10408));
INVX1 gate2373(.O (g20615), .I (g15509));
INVX1 gate2374(.O (g33246), .I (g32212));
INVX1 gate2375(.O (g9083), .I (g626));
INVX1 gate2376(.O (g23875), .I (g18997));
INVX1 gate2377(.O (g25080), .I (g23742));
INVX1 gate2378(.O (g24116), .I (g21143));
INVX1 gate2379(.O (g14518), .I (I16639));
INVX1 gate2380(.O (g23219), .I (I22316));
INVX1 gate2381(.O (I18051), .I (g13680));
INVX1 gate2382(.O (g30330), .I (I28591));
INVX1 gate2383(.O (g13278), .I (g10738));
INVX1 gate2384(.O (g26709), .I (g25435));
INVX1 gate2385(.O (I29969), .I (g30991));
INVX1 gate2386(.O (g8219), .I (g3731));
INVX1 gate2387(.O (g27565), .I (g26645));
INVX1 gate2388(.O (I17491), .I (g13416));
INVX1 gate2389(.O (I16486), .I (g11204));
INVX1 gate2390(.O (g20041), .I (g15569));
INVX1 gate2391(.O (g9636), .I (g72));
INVX1 gate2392(.O (g22214), .I (g19210));
INVX1 gate2393(.O (g7827), .I (g4688));
INVX1 gate2394(.O (g12122), .I (g9705));
INVX1 gate2395(.O (g20275), .I (g17929));
INVX1 gate2396(.O (g24041), .I (g19968));
INVX1 gate2397(.O (g19998), .I (g15915));
INVX1 gate2398(.O (g8431), .I (g3085));
INVX1 gate2399(.O (g11468), .I (g7624));
INVX1 gate2400(.O (g16644), .I (I17842));
INVX1 gate2401(.O (g13039), .I (I15663));
INVX1 gate2402(.O (g8812), .I (I12805));
INVX1 gate2403(.O (g15426), .I (I17121));
INVX1 gate2404(.O (g22207), .I (I21787));
INVX1 gate2405(.O (g6828), .I (g1300));
INVX1 gate2406(.O (g19672), .I (g16931));
INVX1 gate2407(.O (g34132), .I (g33831));
INVX1 gate2408(.O (g17400), .I (I18333));
INVX1 gate2409(.O (I12890), .I (g4219));
INVX1 gate2410(.O (g29045), .I (g27779));
INVX1 gate2411(.O (g34960), .I (I33218));
INVX1 gate2412(.O (g11038), .I (g8632));
INVX1 gate2413(.O (g16969), .I (g14262));
INVX1 gate2414(.O (g6830), .I (g1389));
INVX1 gate2415(.O (g17013), .I (g14262));
INVX1 gate2416(.O (I18350), .I (g13716));
INVX1 gate2417(.O (g8005), .I (g3025));
INVX1 gate2418(.O (g20237), .I (g17213));
INVX1 gate2419(.O (g21160), .I (g17508));
INVX1 gate2420(.O (g7196), .I (I11860));
INVX1 gate2421(.O (g11815), .I (g7582));
INVX1 gate2422(.O (g8405), .I (I12572));
INVX1 gate2423(.O (g9187), .I (g518));
INVX1 gate2424(.O (g16968), .I (g14238));
INVX1 gate2425(.O (I27552), .I (g28162));
INVX1 gate2426(.O (I15677), .I (g5654));
INVX1 gate2427(.O (g31859), .I (g29385));
INVX1 gate2428(.O (I32116), .I (g33937));
INVX1 gate2429(.O (g20035), .I (g16430));
INVX1 gate2430(.O (g31825), .I (g29385));
INVX1 gate2431(.O (g32876), .I (g30735));
INVX1 gate2432(.O (g32885), .I (g31021));
INVX1 gate2433(.O (g34161), .I (g33851));
INVX1 gate2434(.O (g16197), .I (g13861));
INVX1 gate2435(.O (g24035), .I (g20841));
INVX1 gate2436(.O (g11677), .I (g7689));
INVX1 gate2437(.O (g21455), .I (g15426));
INVX1 gate2438(.O (I12003), .I (g767));
INVX1 gate2439(.O (g8286), .I (g53));
INVX1 gate2440(.O (g8765), .I (g3333));
INVX1 gate2441(.O (g17328), .I (I18313));
INVX1 gate2442(.O (g31858), .I (g29385));
INVX1 gate2443(.O (g13975), .I (g11048));
INVX1 gate2444(.O (g32854), .I (g30735));
INVX1 gate2445(.O (g7780), .I (g2878));
INVX1 gate2446(.O (I12779), .I (g4210));
INVX1 gate2447(.O (g16527), .I (g14048));
INVX1 gate2448(.O (g25198), .I (g22228));
INVX1 gate2449(.O (g30259), .I (g28463));
INVX1 gate2450(.O (g25529), .I (g22763));
INVX1 gate2451(.O (g14215), .I (g12198));
INVX1 gate2452(.O (g32511), .I (g30614));
INVX1 gate2453(.O (g23915), .I (g19277));
INVX1 gate2454(.O (g32763), .I (g31710));
INVX1 gate2455(.O (I15937), .I (g11676));
INVX1 gate2456(.O (I17395), .I (g12952));
INVX1 gate2457(.O (I28434), .I (g28114));
INVX1 gate2458(.O (g30087), .I (g29121));
INVX1 gate2459(.O (g11143), .I (g8032));
INVX1 gate2460(.O (g19961), .I (g17328));
INVX1 gate2461(.O (g26810), .I (g25220));
INVX1 gate2462(.O (I29894), .I (g31771));
INVX1 gate2463(.O (I14033), .I (g8912));
INVX1 gate2464(.O (g34471), .I (g34423));
INVX1 gate2465(.O (g9200), .I (g1548));
INVX1 gate2466(.O (g25528), .I (g22594));
INVX1 gate2467(.O (I21934), .I (g21273));
INVX1 gate2468(.O (g31844), .I (g29385));
INVX1 gate2469(.O (I31597), .I (g33187));
INVX1 gate2470(.O (g8733), .I (g3698));
INVX1 gate2471(.O (g19505), .I (g16349));
INVX1 gate2472(.O (g23277), .I (I22380));
INVX1 gate2473(.O (g7018), .I (g5297));
INVX1 gate2474(.O (g8974), .I (I12930));
INVX1 gate2475(.O (I11726), .I (g4273));
INVX1 gate2476(.O (I32237), .I (g34130));
INVX1 gate2477(.O (I17633), .I (g13258));
INVX1 gate2478(.O (g32660), .I (g30825));
INVX1 gate2479(.O (g7418), .I (g2361));
INVX1 gate2480(.O (I13726), .I (g4537));
INVX1 gate2481(.O (g9003), .I (g790));
INVX1 gate2482(.O (g6953), .I (g4157));
INVX1 gate2483(.O (g7994), .I (I12336));
INVX1 gate2484(.O (g29997), .I (g29060));
INVX1 gate2485(.O (g11884), .I (g8125));
INVX1 gate2486(.O (g21467), .I (g15758));
INVX1 gate2487(.O (I16676), .I (g10588));
INVX1 gate2488(.O (g25869), .I (g25250));
INVX1 gate2489(.O (g10349), .I (g6956));
INVX1 gate2490(.O (g23494), .I (I22619));
INVX1 gate2491(.O (g26337), .I (g24818));
INVX1 gate2492(.O (I32806), .I (g34585));
INVX1 gate2493(.O (g8796), .I (g4785));
INVX1 gate2494(.O (I32684), .I (g34430));
INVX1 gate2495(.O (g32456), .I (g31376));
INVX1 gate2496(.O (g34244), .I (I32231));
INVX1 gate2497(.O (I33300), .I (g35001));
INVX1 gate2498(.O (g20130), .I (g17328));
INVX1 gate2499(.O (g22683), .I (I22000));
INVX1 gate2500(.O (g13410), .I (I15921));
INVX1 gate2501(.O (I12826), .I (g4349));
INVX1 gate2502(.O (g21037), .I (I20913));
INVX1 gate2503(.O (g24130), .I (g20998));
INVX1 gate2504(.O (g32480), .I (g31070));
INVX1 gate2505(.O (g10083), .I (g2407));
INVX1 gate2506(.O (g10348), .I (I13762));
INVX1 gate2507(.O (g32916), .I (g31021));
INVX1 gate2508(.O (g14348), .I (g10887));
INVX1 gate2509(.O (g12891), .I (g10399));
INVX1 gate2510(.O (g8324), .I (g2476));
INVX1 gate2511(.O (g26792), .I (g25439));
INVX1 gate2512(.O (g20523), .I (g17821));
INVX1 gate2513(.O (I16417), .I (g875));
INVX1 gate2514(.O (I21013), .I (g15806));
INVX1 gate2515(.O (g32550), .I (g31376));
INVX1 gate2516(.O (g9637), .I (I13252));
INVX1 gate2517(.O (g23984), .I (g19210));
INVX1 gate2518(.O (g18952), .I (g16053));
INVX1 gate2519(.O (g24165), .I (I23339));
INVX1 gate2520(.O (g30068), .I (g29157));
INVX1 gate2521(.O (g34810), .I (I33020));
INVX1 gate2522(.O (g31227), .I (g29744));
INVX1 gate2523(.O (g17683), .I (g15027));
INVX1 gate2524(.O (g23419), .I (g21468));
INVX1 gate2525(.O (g34068), .I (g33728));
INVX1 gate2526(.O (g21352), .I (g16322));
INVX1 gate2527(.O (g13015), .I (g11875));
INVX1 gate2528(.O (g8540), .I (g3408));
INVX1 gate2529(.O (g23352), .I (g20924));
INVX1 gate2530(.O (g25259), .I (I24445));
INVX1 gate2531(.O (g25225), .I (g23802));
INVX1 gate2532(.O (g21155), .I (g15656));
INVX1 gate2533(.O (g34879), .I (I33109));
INVX1 gate2534(.O (g21418), .I (g17821));
INVX1 gate2535(.O (g22882), .I (g20391));
INVX1 gate2536(.O (g28608), .I (g27670));
INVX1 gate2537(.O (g23418), .I (g21468));
INVX1 gate2538(.O (g32721), .I (g31021));
INVX1 gate2539(.O (g20006), .I (g17328));
INVX1 gate2540(.O (I26466), .I (g26870));
INVX1 gate2541(.O (I15556), .I (g11928));
INVX1 gate2542(.O (g32596), .I (g31070));
INVX1 gate2543(.O (g9223), .I (g1216));
INVX1 gate2544(.O (g12109), .I (I14967));
INVX1 gate2545(.O (g19433), .I (g15915));
INVX1 gate2546(.O (g23170), .I (g20046));
INVX1 gate2547(.O (g7197), .I (g812));
INVX1 gate2548(.O (g22407), .I (g19455));
INVX1 gate2549(.O (g34878), .I (I33106));
INVX1 gate2550(.O (g19387), .I (g16431));
INVX1 gate2551(.O (I16762), .I (g5290));
INVX1 gate2552(.O (g6848), .I (g2417));
INVX1 gate2553(.O (g7397), .I (g890));
INVX1 gate2554(.O (I27449), .I (g27737));
INVX1 gate2555(.O (g15969), .I (I17416));
INVX1 gate2556(.O (I20846), .I (g16923));
INVX1 gate2557(.O (g19620), .I (g17296));
INVX1 gate2558(.O (g12108), .I (I14964));
INVX1 gate2559(.O (g10139), .I (g136));
INVX1 gate2560(.O (I15223), .I (g10119));
INVX1 gate2561(.O (I17612), .I (g13250));
INVX1 gate2562(.O (I24396), .I (g23453));
INVX1 gate2563(.O (g6855), .I (g2711));
INVX1 gate2564(.O (g17414), .I (g14627));
INVX1 gate2565(.O (g27492), .I (g26598));
INVX1 gate2566(.O (g8287), .I (g160));
INVX1 gate2567(.O (I17324), .I (g14119));
INVX1 gate2568(.O (g9416), .I (g2429));
INVX1 gate2569(.O (g13223), .I (I15800));
INVX1 gate2570(.O (g24437), .I (g22654));
INVX1 gate2571(.O (g25244), .I (g23802));
INVX1 gate2572(.O (g19343), .I (g16136));
INVX1 gate2573(.O (g34994), .I (I33282));
INVX1 gate2574(.O (I17098), .I (g14336));
INVX1 gate2575(.O (g32773), .I (g31376));
INVX1 gate2576(.O (g32942), .I (g30825));
INVX1 gate2577(.O (g9251), .I (I13037));
INVX1 gate2578(.O (g20703), .I (g15373));
INVX1 gate2579(.O (g29220), .I (I27576));
INVX1 gate2580(.O (I11635), .I (g9));
INVX1 gate2581(.O (g23589), .I (g21468));
INVX1 gate2582(.O (g10415), .I (g7109));
INVX1 gate2583(.O (g18422), .I (I19238));
INVX1 gate2584(.O (g32655), .I (g30614));
INVX1 gate2585(.O (g8399), .I (g3798));
INVX1 gate2586(.O (g11110), .I (g8728));
INVX1 gate2587(.O (g29911), .I (g28780));
INVX1 gate2588(.O (g19369), .I (g15995));
INVX1 gate2589(.O (g33377), .I (I30901));
INVX1 gate2590(.O (g34425), .I (I32446));
INVX1 gate2591(.O (g12381), .I (I15223));
INVX1 gate2592(.O (g23524), .I (g21562));
INVX1 gate2593(.O (g27091), .I (g26725));
INVX1 gate2594(.O (g28184), .I (I26705));
INVX1 gate2595(.O (g32670), .I (g30673));
INVX1 gate2596(.O (g33120), .I (I30686));
INVX1 gate2597(.O (I12026), .I (g344));
INVX1 gate2598(.O (I21100), .I (g16284));
INVX1 gate2599(.O (g8898), .I (g676));
INVX1 gate2600(.O (g20600), .I (g15348));
INVX1 gate2601(.O (I16117), .I (g10430));
INVX1 gate2602(.O (g34919), .I (I33149));
INVX1 gate2603(.O (g19368), .I (g16326));
INVX1 gate2604(.O (I32222), .I (g34118));
INVX1 gate2605(.O (g20781), .I (I20840));
INVX1 gate2606(.O (g16877), .I (I18071));
INVX1 gate2607(.O (g23477), .I (g21468));
INVX1 gate2608(.O (g32734), .I (g31710));
INVX1 gate2609(.O (g33645), .I (I31477));
INVX1 gate2610(.O (g22759), .I (g19857));
INVX1 gate2611(.O (I17140), .I (g13835));
INVX1 gate2612(.O (g26817), .I (g25242));
INVX1 gate2613(.O (g7631), .I (g74));
INVX1 gate2614(.O (g34918), .I (I33146));
INVX1 gate2615(.O (g17584), .I (g14773));
INVX1 gate2616(.O (I26693), .I (g27930));
INVX1 gate2617(.O (g10664), .I (g8928));
INVX1 gate2618(.O (I20929), .I (g17663));
INVX1 gate2619(.O (g32839), .I (g30735));
INVX1 gate2620(.O (g32930), .I (g31021));
INVX1 gate2621(.O (g20372), .I (g17847));
INVX1 gate2622(.O (g30079), .I (g29097));
INVX1 gate2623(.O (g19412), .I (g16489));
INVX1 gate2624(.O (g7257), .I (I11903));
INVX1 gate2625(.O (g22758), .I (g20330));
INVX1 gate2626(.O (g24372), .I (g22885));
INVX1 gate2627(.O (g16695), .I (g14454));
INVX1 gate2628(.O (g25171), .I (g22228));
INVX1 gate2629(.O (g20175), .I (I20433));
INVX1 gate2630(.O (g7301), .I (g925));
INVX1 gate2631(.O (I16747), .I (g12729));
INVX1 gate2632(.O (g8291), .I (I12503));
INVX1 gate2633(.O (g11373), .I (g7566));
INVX1 gate2634(.O (g23864), .I (g19210));
INVX1 gate2635(.O (g25886), .I (g24537));
INVX1 gate2636(.O (g23022), .I (g20283));
INVX1 gate2637(.O (g32667), .I (g30825));
INVX1 gate2638(.O (g32694), .I (g31376));
INVX1 gate2639(.O (g32838), .I (g31376));
INVX1 gate2640(.O (I31550), .I (g33204));
INVX1 gate2641(.O (g33698), .I (I31539));
INVX1 gate2642(.O (g24175), .I (I23369));
INVX1 gate2643(.O (g29147), .I (I27449));
INVX1 gate2644(.O (g32965), .I (g31710));
INVX1 gate2645(.O (g12840), .I (g10356));
INVX1 gate2646(.O (g6818), .I (g976));
INVX1 gate2647(.O (g17759), .I (g14864));
INVX1 gate2648(.O (g6867), .I (I11685));
INVX1 gate2649(.O (g16526), .I (g13898));
INVX1 gate2650(.O (g23749), .I (g18997));
INVX1 gate2651(.O (I15800), .I (g11607));
INVX1 gate2652(.O (g15714), .I (I17228));
INVX1 gate2653(.O (g9880), .I (g5787));
INVX1 gate2654(.O (g23313), .I (g21070));
INVX1 gate2655(.O (g25994), .I (g24575));
INVX1 gate2656(.O (g8344), .I (I12523));
INVX1 gate2657(.O (g9537), .I (g1748));
INVX1 gate2658(.O (g29950), .I (g28896));
INVX1 gate2659(.O (g24063), .I (g20014));
INVX1 gate2660(.O (g17758), .I (g14861));
INVX1 gate2661(.O (g26656), .I (g25495));
INVX1 gate2662(.O (g20516), .I (I20609));
INVX1 gate2663(.O (g10554), .I (g8974));
INVX1 gate2664(.O (g18905), .I (g16077));
INVX1 gate2665(.O (g24137), .I (g20998));
INVX1 gate2666(.O (g32487), .I (g30825));
INVX1 gate2667(.O (g24516), .I (g22670));
INVX1 gate2668(.O (g7751), .I (g1521));
INVX1 gate2669(.O (g23285), .I (g20887));
INVX1 gate2670(.O (g26680), .I (g25300));
INVX1 gate2671(.O (g32619), .I (g30614));
INVX1 gate2672(.O (g8259), .I (g2217));
INVX1 gate2673(.O (g21305), .I (g15758));
INVX1 gate2674(.O (g21053), .I (g15373));
INVX1 gate2675(.O (g32502), .I (g31070));
INVX1 gate2676(.O (g14609), .I (I16724));
INVX1 gate2677(.O (g15979), .I (I17420));
INVX1 gate2678(.O (g10200), .I (g2138));
INVX1 gate2679(.O (g23305), .I (g20391));
INVX1 gate2680(.O (g32557), .I (g31376));
INVX1 gate2681(.O (g13334), .I (g11048));
INVX1 gate2682(.O (g29151), .I (g27858));
INVX1 gate2683(.O (g29172), .I (g27020));
INVX1 gate2684(.O (I24787), .I (g24266));
INVX1 gate2685(.O (g9978), .I (g2756));
INVX1 gate2686(.O (g30322), .I (g28431));
INVX1 gate2687(.O (g10608), .I (g9155));
INVX1 gate2688(.O (g29996), .I (g28962));
INVX1 gate2689(.O (I12811), .I (g4340));
INVX1 gate2690(.O (g10115), .I (g2283));
INVX1 gate2691(.O (I16639), .I (g4000));
INVX1 gate2692(.O (g21466), .I (g15509));
INVX1 gate2693(.O (g32618), .I (g31154));
INVX1 gate2694(.O (I18662), .I (g6322));
INVX1 gate2695(.O (g8088), .I (g1554));
INVX1 gate2696(.O (g6975), .I (g4507));
INVX1 gate2697(.O (g9417), .I (I13124));
INVX1 gate2698(.O (g34159), .I (I32116));
INVX1 gate2699(.O (g11762), .I (g7964));
INVX1 gate2700(.O (g7041), .I (g5644));
INVX1 gate2701(.O (g9935), .I (I13483));
INVX1 gate2702(.O (I13606), .I (g74));
INVX1 gate2703(.O (g11964), .I (g9154));
INVX1 gate2704(.O (g21036), .I (I20910));
INVX1 gate2705(.O (g7441), .I (g862));
INVX1 gate2706(.O (g20209), .I (g17821));
INVX1 gate2707(.O (g33661), .I (I31497));
INVX1 gate2708(.O (g33895), .I (I31751));
INVX1 gate2709(.O (g9982), .I (g3976));
INVX1 gate2710(.O (g21177), .I (I20957));
INVX1 gate2711(.O (g21560), .I (g17873));
INVX1 gate2712(.O (g16077), .I (I17456));
INVX1 gate2713(.O (g9234), .I (g5170));
INVX1 gate2714(.O (I15587), .I (g11985));
INVX1 gate2715(.O (g32469), .I (g30673));
INVX1 gate2716(.O (I27368), .I (g27881));
INVX1 gate2717(.O (I18482), .I (g13350));
INVX1 gate2718(.O (g20208), .I (g17533));
INVX1 gate2719(.O (g14745), .I (g12423));
INVX1 gate2720(.O (g13216), .I (g10939));
INVX1 gate2721(.O (g17141), .I (I18191));
INVX1 gate2722(.O (I11750), .I (g4474));
INVX1 gate2723(.O (I18248), .I (g12938));
INVX1 gate2724(.O (g19379), .I (g17327));
INVX1 gate2725(.O (g26631), .I (g25467));
INVX1 gate2726(.O (g12862), .I (g10370));
INVX1 gate2727(.O (g17652), .I (g15033));
INVX1 gate2728(.O (g34656), .I (I32770));
INVX1 gate2729(.O (g8215), .I (I12451));
INVX1 gate2730(.O (g30295), .I (I28540));
INVX1 gate2731(.O (g22332), .I (I21838));
INVX1 gate2732(.O (g9542), .I (g2173));
INVX1 gate2733(.O (I16391), .I (g859));
INVX1 gate2734(.O (g26364), .I (I25327));
INVX1 gate2735(.O (g32468), .I (g30614));
INVX1 gate2736(.O (g6821), .I (I11655));
INVX1 gate2737(.O (I18003), .I (g13638));
INVX1 gate2738(.O (g19050), .I (I19759));
INVX1 gate2739(.O (g34680), .I (I32820));
INVX1 gate2740(.O (g8951), .I (g554));
INVX1 gate2741(.O (g16689), .I (g13923));
INVX1 gate2742(.O (g34144), .I (I32093));
INVX1 gate2743(.O (g34823), .I (I33037));
INVX1 gate2744(.O (g20542), .I (g17873));
INVX1 gate2745(.O (g16923), .I (I18089));
INVX1 gate2746(.O (g20453), .I (I20584));
INVX1 gate2747(.O (g16280), .I (g13330));
INVX1 gate2748(.O (g6984), .I (g4709));
INVX1 gate2749(.O (g32038), .I (g30934));
INVX1 gate2750(.O (g24021), .I (g20841));
INVX1 gate2751(.O (g28241), .I (g27064));
INVX1 gate2752(.O (g29318), .I (g29029));
INVX1 gate2753(.O (g16688), .I (g14045));
INVX1 gate2754(.O (g16624), .I (I17814));
INVX1 gate2755(.O (g22406), .I (g19506));
INVX1 gate2756(.O (g8114), .I (g3522));
INVX1 gate2757(.O (g10184), .I (g4486));
INVX1 gate2758(.O (g12040), .I (I14902));
INVX1 gate2759(.O (I16579), .I (g10981));
INVX1 gate2760(.O (g16300), .I (I17626));
INVX1 gate2761(.O (g19386), .I (g16431));
INVX1 gate2762(.O (g10805), .I (I14046));
INVX1 gate2763(.O (I22785), .I (g18940));
INVX1 gate2764(.O (g20913), .I (g15373));
INVX1 gate2765(.O (I18778), .I (g6704));
INVX1 gate2766(.O (g34336), .I (g34112));
INVX1 gate2767(.O (g32815), .I (g30937));
INVX1 gate2768(.O (g14184), .I (g12381));
INVX1 gate2769(.O (g19603), .I (g16349));
INVX1 gate2770(.O (g19742), .I (g17096));
INVX1 gate2771(.O (g13117), .I (g10981));
INVX1 gate2772(.O (g17135), .I (g14297));
INVX1 gate2773(.O (g12904), .I (g10410));
INVX1 gate2774(.O (g20614), .I (g15426));
INVX1 gate2775(.O (g32601), .I (g31376));
INVX1 gate2776(.O (I15569), .I (g11965));
INVX1 gate2777(.O (g9554), .I (g5105));
INVX1 gate2778(.O (g20436), .I (I20569));
INVX1 gate2779(.O (g23874), .I (g18997));
INVX1 gate2780(.O (g8870), .I (I12837));
INVX1 gate2781(.O (g32677), .I (g30673));
INVX1 gate2782(.O (g33127), .I (g31950));
INVX1 gate2783(.O (g25322), .I (I24497));
INVX1 gate2784(.O (I31694), .I (g33176));
INVX1 gate2785(.O (I32834), .I (g34472));
INVX1 gate2786(.O (g32975), .I (I30537));
INVX1 gate2787(.O (g21693), .I (I21254));
INVX1 gate2788(.O (g20607), .I (g17955));
INVX1 gate2789(.O (g13569), .I (g10951));
INVX1 gate2790(.O (g8650), .I (g4664));
INVX1 gate2791(.O (I12896), .I (g4229));
INVX1 gate2792(.O (g20320), .I (g17015));
INVX1 gate2793(.O (I18647), .I (g5320));
INVX1 gate2794(.O (g20073), .I (g16540));
INVX1 gate2795(.O (I28832), .I (g30301));
INVX1 gate2796(.O (I33131), .I (g34906));
INVX1 gate2797(.O (g30017), .I (g29085));
INVX1 gate2798(.O (g20274), .I (g17847));
INVX1 gate2799(.O (g9213), .I (I13020));
INVX1 gate2800(.O (g24073), .I (g21127));
INVX1 gate2801(.O (g20530), .I (g15509));
INVX1 gate2802(.O (g21665), .I (I21226));
INVX1 gate2803(.O (g25158), .I (g22228));
INVX1 gate2804(.O (I21744), .I (g19338));
INVX1 gate2805(.O (g20593), .I (g15277));
INVX1 gate2806(.O (I17754), .I (g13494));
INVX1 gate2807(.O (g23665), .I (g21562));
INVX1 gate2808(.O (g25783), .I (g25250));
INVX1 gate2809(.O (I17355), .I (g14591));
INVX1 gate2810(.O (g32937), .I (g31021));
INVX1 gate2811(.O (g19429), .I (g16489));
INVX1 gate2812(.O (I23345), .I (g23320));
INVX1 gate2813(.O (g33385), .I (g32038));
INVX1 gate2814(.O (I21849), .I (g19620));
INVX1 gate2815(.O (g29044), .I (g27742));
INVX1 gate2816(.O (g10761), .I (g8411));
INVX1 gate2817(.O (g7411), .I (g2040));
INVX1 gate2818(.O (g25561), .I (g22550));
INVX1 gate2819(.O (g18891), .I (g16053));
INVX1 gate2820(.O (g20565), .I (g18008));
INVX1 gate2821(.O (I31619), .I (g33212));
INVX1 gate2822(.O (I15814), .I (g11129));
INVX1 gate2823(.O (g24122), .I (g20857));
INVX1 gate2824(.O (I23399), .I (g23450));
INVX1 gate2825(.O (g8136), .I (g269));
INVX1 gate2826(.O (g19730), .I (g17062));
INVX1 gate2827(.O (g19428), .I (g16090));
INVX1 gate2828(.O (g12183), .I (I15033));
INVX1 gate2829(.O (g9902), .I (g100));
INVX1 gate2830(.O (I18233), .I (g14639));
INVX1 gate2831(.O (g33354), .I (g32329));
INVX1 gate2832(.O (I33210), .I (g34943));
INVX1 gate2833(.O (g32791), .I (g31672));
INVX1 gate2834(.O (g23476), .I (g21468));
INVX1 gate2835(.O (g23485), .I (g20785));
INVX1 gate2836(.O (I25555), .I (g25241));
INVX1 gate2837(.O (g31824), .I (g29385));
INVX1 gate2838(.O (g32884), .I (g30825));
INVX1 gate2839(.O (g33888), .I (g33346));
INVX1 gate2840(.O (g8594), .I (g3849));
INVX1 gate2841(.O (g19765), .I (g16897));
INVX1 gate2842(.O (g6756), .I (I11623));
INVX1 gate2843(.O (g24034), .I (g19968));
INVX1 gate2844(.O (g7074), .I (I11801));
INVX1 gate2845(.O (g11772), .I (I14623));
INVX1 gate2846(.O (g10400), .I (g7002));
INVX1 gate2847(.O (g20641), .I (g15509));
INVX1 gate2848(.O (g26816), .I (g25260));
INVX1 gate2849(.O (g21454), .I (g15373));
INVX1 gate2850(.O (I33279), .I (g34986));
INVX1 gate2851(.O (g23555), .I (I22692));
INVX1 gate2852(.O (I32607), .I (g34358));
INVX1 gate2853(.O (g7474), .I (I11980));
INVX1 gate2854(.O (g17221), .I (I18245));
INVX1 gate2855(.O (g19690), .I (g16826));
INVX1 gate2856(.O (g30309), .I (g28959));
INVX1 gate2857(.O (g7992), .I (g5008));
INVX1 gate2858(.O (g9490), .I (g2563));
INVX1 gate2859(.O (I14563), .I (g802));
INVX1 gate2860(.O (g16511), .I (g14130));
INVX1 gate2861(.O (g9166), .I (g837));
INVX1 gate2862(.O (g20153), .I (g16782));
INVX1 gate2863(.O (g23570), .I (g18833));
INVX1 gate2864(.O (I32274), .I (g34195));
INVX1 gate2865(.O (g23914), .I (g19210));
INVX1 gate2866(.O (g32479), .I (g30735));
INVX1 gate2867(.O (g32666), .I (g31376));
INVX1 gate2868(.O (I13483), .I (g6035));
INVX1 gate2869(.O (g11293), .I (g7527));
INVX1 gate2870(.O (g24153), .I (I23303));
INVX1 gate2871(.O (I31469), .I (g33388));
INVX1 gate2872(.O (g6904), .I (g3494));
INVX1 gate2873(.O (g32363), .I (I29891));
INVX1 gate2874(.O (I12112), .I (g794));
INVX1 gate2875(.O (g12872), .I (g10379));
INVX1 gate2876(.O (g13638), .I (I16057));
INVX1 gate2877(.O (g34308), .I (g34088));
INVX1 gate2878(.O (g9056), .I (g3017));
INVX1 gate2879(.O (g23907), .I (g19074));
INVX1 gate2880(.O (g32478), .I (g31376));
INVX1 gate2881(.O (g32015), .I (I29571));
INVX1 gate2882(.O (g19504), .I (g16349));
INVX1 gate2883(.O (g9456), .I (g6073));
INVX1 gate2884(.O (g33931), .I (I31807));
INVX1 gate2885(.O (I32464), .I (g34245));
INVX1 gate2886(.O (g8228), .I (g3835));
INVX1 gate2887(.O (g9529), .I (g6561));
INVX1 gate2888(.O (g7863), .I (g1249));
INVX1 gate2889(.O (g20136), .I (I20399));
INVX1 gate2890(.O (g20635), .I (g18008));
INVX1 gate2891(.O (I27742), .I (g28819));
INVX1 gate2892(.O (g13416), .I (I15929));
INVX1 gate2893(.O (g25017), .I (g23699));
INVX1 gate2894(.O (I25567), .I (g25272));
INVX1 gate2895(.O (I25594), .I (g25531));
INVX1 gate2896(.O (I18897), .I (g16738));
INVX1 gate2897(.O (g24136), .I (g20857));
INVX1 gate2898(.O (g32486), .I (g30735));
INVX1 gate2899(.O (I13326), .I (g66));
INVX1 gate2900(.O (g23239), .I (g21308));
INVX1 gate2901(.O (g33426), .I (g32017));
INVX1 gate2902(.O (g11841), .I (g9800));
INVX1 gate2903(.O (g9155), .I (I12997));
INVX1 gate2904(.O (I14395), .I (g3654));
INVX1 gate2905(.O (g6841), .I (g2145));
INVX1 gate2906(.O (I17420), .I (g13394));
INVX1 gate2907(.O (g23567), .I (g21562));
INVX1 gate2908(.O (g32556), .I (g31554));
INVX1 gate2909(.O (I32797), .I (g34581));
INVX1 gate2910(.O (I14899), .I (g10198));
INVX1 gate2911(.O (g8033), .I (g157));
INVX1 gate2912(.O (g23238), .I (g20924));
INVX1 gate2913(.O (g11510), .I (g7633));
INVX1 gate2914(.O (g13510), .I (I15981));
INVX1 gate2915(.O (g17812), .I (I18810));
INVX1 gate2916(.O (g34816), .I (I33030));
INVX1 gate2917(.O (I20647), .I (g17010));
INVX1 gate2918(.O (g32580), .I (g30825));
INVX1 gate2919(.O (g9698), .I (g2181));
INVX1 gate2920(.O (g28441), .I (g27629));
INVX1 gate2921(.O (g26260), .I (g24759));
INVX1 gate2922(.O (I14633), .I (g9340));
INVX1 gate2923(.O (g9964), .I (g126));
INVX1 gate2924(.O (I13252), .I (g6751));
INVX1 gate2925(.O (g20164), .I (g16826));
INVX1 gate2926(.O (g34985), .I (I33255));
INVX1 gate2927(.O (I20999), .I (g16709));
INVX1 gate2928(.O (g23941), .I (g19074));
INVX1 gate2929(.O (g18091), .I (I18879));
INVX1 gate2930(.O (g19128), .I (I19778));
INVX1 gate2931(.O (g23382), .I (g20682));
INVX1 gate2932(.O (g24164), .I (I23336));
INVX1 gate2933(.O (g25289), .I (g22228));
INVX1 gate2934(.O (g21176), .I (I20954));
INVX1 gate2935(.O (g21185), .I (g15277));
INVX1 gate2936(.O (g23519), .I (g21468));
INVX1 gate2937(.O (I27730), .I (g28752));
INVX1 gate2938(.O (g12047), .I (g9591));
INVX1 gate2939(.O (g16307), .I (I17633));
INVX1 gate2940(.O (g13835), .I (I16150));
INVX1 gate2941(.O (g34954), .I (I33210));
INVX1 gate2942(.O (g13014), .I (g11872));
INVX1 gate2943(.O (g25023), .I (g22457));
INVX1 gate2944(.O (g24891), .I (g23231));
INVX1 gate2945(.O (I33143), .I (g34903));
INVX1 gate2946(.O (g19626), .I (g17409));
INVX1 gate2947(.O (g25288), .I (g22228));
INVX1 gate2948(.O (g25224), .I (g22763));
INVX1 gate2949(.O (I20233), .I (g17487));
INVX1 gate2950(.O (g16721), .I (g14072));
INVX1 gate2951(.O (I12793), .I (g4578));
INVX1 gate2952(.O (g23518), .I (g21070));
INVX1 gate2953(.O (g23154), .I (I22264));
INVX1 gate2954(.O (g26488), .I (I25366));
INVX1 gate2955(.O (g26424), .I (I25356));
INVX1 gate2956(.O (g20575), .I (g17929));
INVX1 gate2957(.O (g31860), .I (I29438));
INVX1 gate2958(.O (g13007), .I (g11852));
INVX1 gate2959(.O (g25308), .I (g22763));
INVX1 gate2960(.O (g8195), .I (g1783));
INVX1 gate2961(.O (g8137), .I (g411));
INVX1 gate2962(.O (g32922), .I (g31710));
INVX1 gate2963(.O (g8891), .I (g582));
INVX1 gate2964(.O (g19533), .I (g16261));
INVX1 gate2965(.O (g24474), .I (g23620));
INVX1 gate2966(.O (g20711), .I (g15509));
INVX1 gate2967(.O (I16193), .I (g3281));
INVX1 gate2968(.O (g16431), .I (I17675));
INVX1 gate2969(.O (I27549), .I (g28161));
INVX1 gate2970(.O (g27051), .I (I25779));
INVX1 gate2971(.O (g32531), .I (g31070));
INVX1 gate2972(.O (I13847), .I (g7266));
INVX1 gate2973(.O (I31791), .I (g33354));
INVX1 gate2974(.O (g20327), .I (g15224));
INVX1 gate2975(.O (g23935), .I (g19210));
INVX1 gate2976(.O (g24711), .I (g23139));
INVX1 gate2977(.O (g34669), .I (I32791));
INVX1 gate2978(.O (g26830), .I (g24411));
INVX1 gate2979(.O (g27592), .I (g26715));
INVX1 gate2980(.O (g12051), .I (g9595));
INVX1 gate2981(.O (g20537), .I (g15345));
INVX1 gate2982(.O (g24109), .I (g21143));
INVX1 gate2983(.O (g32740), .I (g31672));
INVX1 gate2984(.O (g15885), .I (I17374));
INVX1 gate2985(.O (g8807), .I (g79));
INVX1 gate2986(.O (g11615), .I (g6875));
INVX1 gate2987(.O (g9619), .I (g5845));
INVX1 gate2988(.O (g17507), .I (g15030));
INVX1 gate2989(.O (I24331), .I (g22976));
INVX1 gate2990(.O (g34668), .I (I32788));
INVX1 gate2991(.O (g13116), .I (g10935));
INVX1 gate2992(.O (g16773), .I (g14021));
INVX1 gate2993(.O (I18148), .I (g13526));
INVX1 gate2994(.O (g24108), .I (g20998));
INVX1 gate2995(.O (I28162), .I (g28803));
INVX1 gate2996(.O (g32186), .I (I29720));
INVX1 gate2997(.O (g34392), .I (g34202));
INVX1 gate2998(.O (g32676), .I (g30614));
INVX1 gate2999(.O (g32685), .I (g31528));
INVX1 gate3000(.O (g33659), .I (I31491));
INVX1 gate3001(.O (g28399), .I (g27074));
INVX1 gate3002(.O (g30195), .I (I28434));
INVX1 gate3003(.O (g7400), .I (g911));
INVX1 gate3004(.O (g8859), .I (g772));
INVX1 gate3005(.O (g32953), .I (g31327));
INVX1 gate3006(.O (g19737), .I (g17015));
INVX1 gate3007(.O (g11720), .I (I14589));
INVX1 gate3008(.O (g20283), .I (I20529));
INVX1 gate3009(.O (g6811), .I (g714));
INVX1 gate3010(.O (g34195), .I (I32150));
INVX1 gate3011(.O (g20606), .I (g17955));
INVX1 gate3012(.O (g33250), .I (g32186));
INVX1 gate3013(.O (g16655), .I (g14151));
INVX1 gate3014(.O (g10882), .I (g7601));
INVX1 gate3015(.O (I18104), .I (g13177));
INVX1 gate3016(.O (g10414), .I (g7092));
INVX1 gate3017(.O (I13634), .I (g79));
INVX1 gate3018(.O (g31658), .I (I29242));
INVX1 gate3019(.O (I13872), .I (g7474));
INVX1 gate3020(.O (g13041), .I (I15667));
INVX1 gate3021(.O (g32654), .I (g31070));
INVX1 gate3022(.O (g9843), .I (g4311));
INVX1 gate3023(.O (g33658), .I (g33080));
INVX1 gate3024(.O (g16180), .I (g13437));
INVX1 gate3025(.O (g30016), .I (g29049));
INVX1 gate3026(.O (g9989), .I (g5077));
INVX1 gate3027(.O (I24448), .I (g22923));
INVX1 gate3028(.O (g11430), .I (g7617));
INVX1 gate3029(.O (g22541), .I (I21911));
INVX1 gate3030(.O (g34559), .I (g34384));
INVX1 gate3031(.O (g12350), .I (I15190));
INVX1 gate3032(.O (g10407), .I (g7063));
INVX1 gate3033(.O (g32800), .I (g31021));
INVX1 gate3034(.O (g32936), .I (g31710));
INVX1 gate3035(.O (g19697), .I (g16886));
INVX1 gate3036(.O (I31486), .I (g33197));
INVX1 gate3037(.O (g23215), .I (g20785));
INVX1 gate3038(.O (g12820), .I (g10233));
INVX1 gate3039(.O (I17699), .I (g13416));
INVX1 gate3040(.O (g23501), .I (g20924));
INVX1 gate3041(.O (g6874), .I (g3143));
INVX1 gate3042(.O (I29965), .I (g31189));
INVX1 gate3043(.O (I32109), .I (g33631));
INVX1 gate3044(.O (I21033), .I (g17221));
INVX1 gate3045(.O (g20381), .I (g17955));
INVX1 gate3046(.O (g8342), .I (I12519));
INVX1 gate3047(.O (g11237), .I (I14305));
INVX1 gate3048(.O (g9834), .I (g2579));
INVX1 gate3049(.O (g9971), .I (g2093));
INVX1 gate3050(.O (I21234), .I (g16540));
INVX1 gate3051(.O (g24982), .I (g22763));
INVX1 gate3052(.O (g26679), .I (g25385));
INVX1 gate3053(.O (g34830), .I (I33044));
INVX1 gate3054(.O (g34893), .I (I33119));
INVX1 gate3055(.O (g9686), .I (g73));
INVX1 gate3056(.O (g22359), .I (g19495));
INVX1 gate3057(.O (g8255), .I (g2028));
INVX1 gate3058(.O (g17473), .I (g14841));
INVX1 gate3059(.O (g20091), .I (g17328));
INVX1 gate3060(.O (I22366), .I (g19757));
INVX1 gate3061(.O (g24091), .I (g20720));
INVX1 gate3062(.O (g7183), .I (g4608));
INVX1 gate3063(.O (g8481), .I (I12618));
INVX1 gate3064(.O (I12128), .I (g4253));
INVX1 gate3065(.O (g17789), .I (g14321));
INVX1 gate3066(.O (g29956), .I (I28185));
INVX1 gate3067(.O (g29385), .I (g28180));
INVX1 gate3068(.O (g34544), .I (I32613));
INVX1 gate3069(.O (g15480), .I (I17125));
INVX1 gate3070(.O (I26664), .I (g27708));
INVX1 gate3071(.O (g22358), .I (g19801));
INVX1 gate3072(.O (g32762), .I (g31672));
INVX1 gate3073(.O (g9598), .I (g2571));
INVX1 gate3074(.O (g24174), .I (I23366));
INVX1 gate3075(.O (g8097), .I (g3029));
INVX1 gate3076(.O (g25260), .I (I24448));
INVX1 gate3077(.O (g32964), .I (g31672));
INVX1 gate3078(.O (g29980), .I (g28935));
INVX1 gate3079(.O (g7779), .I (g1413));
INVX1 gate3080(.O (g34713), .I (I32871));
INVX1 gate3081(.O (g8497), .I (g3436));
INVX1 gate3082(.O (g13142), .I (g10632));
INVX1 gate3083(.O (g21349), .I (g15758));
INVX1 gate3084(.O (g8154), .I (g3139));
INVX1 gate3085(.O (I28591), .I (g29371));
INVX1 gate3086(.O (g17325), .I (I18304));
INVX1 gate3087(.O (g8354), .I (g4815));
INVX1 gate3088(.O (g18948), .I (g15800));
INVX1 gate3089(.O (g7023), .I (g5445));
INVX1 gate3090(.O (g31855), .I (g29385));
INVX1 gate3091(.O (g10206), .I (g4489));
INVX1 gate3092(.O (g14441), .I (I16590));
INVX1 gate3093(.O (g14584), .I (g11048));
INVX1 gate3094(.O (g9321), .I (g5863));
INVX1 gate3095(.O (g7423), .I (g2433));
INVX1 gate3096(.O (g9670), .I (g5022));
INVX1 gate3097(.O (I22547), .I (g20720));
INVX1 gate3098(.O (g25195), .I (g22763));
INVX1 gate3099(.O (g16487), .I (I17695));
INVX1 gate3100(.O (g23906), .I (g19074));
INVX1 gate3101(.O (g26093), .I (g24814));
INVX1 gate3102(.O (g30610), .I (I28872));
INVX1 gate3103(.O (g18904), .I (g16053));
INVX1 gate3104(.O (g32587), .I (g30735));
INVX1 gate3105(.O (g15085), .I (I17008));
INVX1 gate3106(.O (I32982), .I (g34749));
INVX1 gate3107(.O (g23284), .I (g20785));
INVX1 gate3108(.O (g19445), .I (g15915));
INVX1 gate3109(.O (g10725), .I (g7846));
INVX1 gate3110(.O (g21304), .I (g17367));
INVX1 gate3111(.O (g25525), .I (g22550));
INVX1 gate3112(.O (g34042), .I (g33674));
INVX1 gate3113(.O (g25424), .I (g23800));
INVX1 gate3114(.O (I20433), .I (g16234));
INVX1 gate3115(.O (g23304), .I (g20785));
INVX1 gate3116(.O (g25016), .I (g23666));
INVX1 gate3117(.O (g6978), .I (g4616));
INVX1 gate3118(.O (I33179), .I (g34893));
INVX1 gate3119(.O (g7161), .I (I11843));
INVX1 gate3120(.O (g19499), .I (g16782));
INVX1 gate3121(.O (g17121), .I (g14321));
INVX1 gate3122(.O (g7361), .I (g1874));
INVX1 gate3123(.O (g22682), .I (g19379));
INVX1 gate3124(.O (g10114), .I (g2116));
INVX1 gate3125(.O (g20192), .I (g17268));
INVX1 gate3126(.O (g9253), .I (g5037));
INVX1 gate3127(.O (I16821), .I (g5983));
INVX1 gate3128(.O (I17661), .I (g13329));
INVX1 gate3129(.O (g27929), .I (I26448));
INVX1 gate3130(.O (g25558), .I (g22594));
INVX1 gate3131(.O (g23566), .I (g21562));
INVX1 gate3132(.O (g32909), .I (g30614));
INVX1 gate3133(.O (g10082), .I (g2375));
INVX1 gate3134(.O (g32543), .I (g31376));
INVX1 gate3135(.O (g34270), .I (g34159));
INVX1 gate3136(.O (I27232), .I (g27993));
INVX1 gate3137(.O (g19498), .I (g16752));
INVX1 gate3138(.O (g34188), .I (g33875));
INVX1 gate3139(.O (g7051), .I (I11793));
INVX1 gate3140(.O (g10107), .I (I13606));
INVX1 gate3141(.O (g22173), .I (I21757));
INVX1 gate3142(.O (g34124), .I (g33819));
INVX1 gate3143(.O (g9909), .I (g1978));
INVX1 gate3144(.O (g12929), .I (g12550));
INVX1 gate3145(.O (g25830), .I (g24485));
INVX1 gate3146(.O (g27583), .I (g26686));
INVX1 gate3147(.O (g20663), .I (g15373));
INVX1 gate3148(.O (g27928), .I (g26810));
INVX1 gate3149(.O (g25893), .I (g24541));
INVX1 gate3150(.O (g8783), .I (I12761));
INVX1 gate3151(.O (g7451), .I (g2070));
INVX1 gate3152(.O (g32908), .I (g31327));
INVX1 gate3153(.O (g6982), .I (g4531));
INVX1 gate3154(.O (g7327), .I (g2165));
INVX1 gate3155(.O (g24522), .I (g22689));
INVX1 gate3156(.O (g33894), .I (I31748));
INVX1 gate3157(.O (g11165), .I (I14222));
INVX1 gate3158(.O (g8112), .I (g3419));
INVX1 gate3159(.O (g8218), .I (g3490));
INVX1 gate3160(.O (g34939), .I (g34922));
INVX1 gate3161(.O (g9740), .I (g5821));
INVX1 gate3162(.O (g8267), .I (g2342));
INVX1 gate3163(.O (g25544), .I (g22594));
INVX1 gate3164(.O (g32569), .I (g30673));
INVX1 gate3165(.O (g34383), .I (I32388));
INVX1 gate3166(.O (g29190), .I (g27046));
INVX1 gate3167(.O (I32840), .I (g34480));
INVX1 gate3168(.O (g17291), .I (I18276));
INVX1 gate3169(.O (g14744), .I (g12578));
INVX1 gate3170(.O (g16286), .I (I17615));
INVX1 gate3171(.O (g21139), .I (g15634));
INVX1 gate3172(.O (g21653), .I (g17663));
INVX1 gate3173(.O (g26837), .I (g24869));
INVX1 gate3174(.O (g7633), .I (I12120));
INVX1 gate3175(.O (g34938), .I (g34920));
INVX1 gate3176(.O (g23653), .I (I22788));
INVX1 gate3177(.O (g9552), .I (g3654));
INVX1 gate3178(.O (g15655), .I (g13202));
INVX1 gate3179(.O (I31800), .I (g33164));
INVX1 gate3180(.O (g10399), .I (g7017));
INVX1 gate3181(.O (g32568), .I (g31170));
INVX1 gate3182(.O (g32747), .I (g30825));
INVX1 gate3183(.O (I18310), .I (g12978));
INVX1 gate3184(.O (I20369), .I (g17690));
INVX1 gate3185(.O (g18062), .I (I18872));
INVX1 gate3186(.O (g21138), .I (g15634));
INVX1 gate3187(.O (g24483), .I (I23688));
INVX1 gate3188(.O (g19432), .I (g15885));
INVX1 gate3189(.O (I19837), .I (g1399));
INVX1 gate3190(.O (g30065), .I (g29049));
INVX1 gate3191(.O (I11820), .I (g3869));
INVX1 gate3192(.O (g23138), .I (g20453));
INVX1 gate3193(.O (I26799), .I (g27660));
INVX1 gate3194(.O (g20553), .I (g17929));
INVX1 gate3195(.O (g31819), .I (g29385));
INVX1 gate3196(.O (g8676), .I (g4821));
INVX1 gate3197(.O (I15727), .I (g10981));
INVX1 gate3198(.O (I32192), .I (g33628));
INVX1 gate3199(.O (g10398), .I (g6999));
INVX1 gate3200(.O (I18379), .I (g13012));
INVX1 gate3201(.O (g14398), .I (I16555));
INVX1 gate3202(.O (g10141), .I (I13634));
INVX1 gate3203(.O (g29211), .I (I27549));
INVX1 gate3204(.O (g10652), .I (g7601));
INVX1 gate3205(.O (g10804), .I (g9772));
INVX1 gate3206(.O (g6800), .I (g203));
INVX1 gate3207(.O (I13152), .I (g6746));
INVX1 gate3208(.O (g9687), .I (I13287));
INVX1 gate3209(.O (g31818), .I (g29385));
INVX1 gate3210(.O (g32814), .I (g31021));
INVX1 gate3211(.O (g20326), .I (g18008));
INVX1 gate3212(.O (g23333), .I (g20785));
INVX1 gate3213(.O (g13222), .I (g10590));
INVX1 gate3214(.O (g19753), .I (g16987));
INVX1 gate3215(.O (g16601), .I (I17783));
INVX1 gate3216(.O (g17760), .I (I18752));
INVX1 gate3217(.O (g16677), .I (I17879));
INVX1 gate3218(.O (I22889), .I (g18926));
INVX1 gate3219(.O (g20536), .I (g18065));
INVX1 gate3220(.O (g20040), .I (g17271));
INVX1 gate3221(.O (g13437), .I (I15937));
INVX1 gate3222(.O (I20412), .I (g16213));
INVX1 gate3223(.O (g32751), .I (g31327));
INVX1 gate3224(.O (g32807), .I (g31021));
INVX1 gate3225(.O (g32772), .I (g31327));
INVX1 gate3226(.O (g28463), .I (I26952));
INVX1 gate3227(.O (g32974), .I (g30937));
INVX1 gate3228(.O (g8830), .I (g767));
INVX1 gate3229(.O (g24040), .I (g19919));
INVX1 gate3230(.O (g7753), .I (I12183));
INVX1 gate3231(.O (g20702), .I (g17955));
INVX1 gate3232(.O (g30218), .I (g28918));
INVX1 gate3233(.O (g25188), .I (g23909));
INVX1 gate3234(.O (g32639), .I (g31070));
INVX1 gate3235(.O (g20904), .I (g17433));
INVX1 gate3236(.O (I17956), .I (g14562));
INVX1 gate3237(.O (g23963), .I (g19147));
INVX1 gate3238(.O (g19650), .I (g16971));
INVX1 gate3239(.O (g28033), .I (g26365));
INVX1 gate3240(.O (g8592), .I (g3805));
INVX1 gate3241(.O (g7072), .I (g6199));
INVX1 gate3242(.O (g14332), .I (I16492));
INVX1 gate3243(.O (I11691), .I (g36));
INVX1 gate3244(.O (I28540), .I (g28954));
INVX1 gate3245(.O (g32638), .I (g30825));
INVX1 gate3246(.O (g7472), .I (g6329));
INVX1 gate3247(.O (g19529), .I (g16349));
INVX1 gate3248(.O (g12640), .I (I15382));
INVX1 gate3249(.O (I15600), .I (g10430));
INVX1 gate3250(.O (g22927), .I (I22128));
INVX1 gate3251(.O (g9860), .I (g5417));
INVX1 gate3252(.O (g10406), .I (g7046));
INVX1 gate3253(.O (I24228), .I (g22409));
INVX1 gate3254(.O (g20564), .I (g15373));
INVX1 gate3255(.O (g10361), .I (g6841));
INVX1 gate3256(.O (I25576), .I (g25296));
INVX1 gate3257(.O (g7443), .I (g914));
INVX1 gate3258(.O (g8703), .I (I12709));
INVX1 gate3259(.O (g14406), .I (g12249));
INVX1 gate3260(.O (g19528), .I (g16349));
INVX1 gate3261(.O (g19696), .I (g17015));
INVX1 gate3262(.O (g34160), .I (I32119));
INVX1 gate3263(.O (g25267), .I (g22228));
INVX1 gate3264(.O (g19330), .I (g17326));
INVX1 gate3265(.O (I17181), .I (g13745));
INVX1 gate3266(.O (I17671), .I (g13280));
INVX1 gate3267(.O (I29363), .I (g30218));
INVX1 gate3268(.O (g23585), .I (g21070));
INVX1 gate3269(.O (g32841), .I (g31672));
INVX1 gate3270(.O (g11236), .I (g8357));
INVX1 gate3271(.O (I21291), .I (g18273));
INVX1 gate3272(.O (g7116), .I (g22));
INVX1 gate3273(.O (g22649), .I (g19063));
INVX1 gate3274(.O (g10500), .I (I13875));
INVX1 gate3275(.O (g27881), .I (I26430));
INVX1 gate3276(.O (g19365), .I (g16249));
INVX1 gate3277(.O (g20673), .I (g15277));
INVX1 gate3278(.O (g32510), .I (g31194));
INVX1 gate3279(.O (g9691), .I (g1706));
INVX1 gate3280(.O (g31801), .I (g29385));
INVX1 gate3281(.O (I15821), .I (g11143));
INVX1 gate3282(.O (I12056), .I (g2748));
INVX1 gate3283(.O (g24183), .I (I23393));
INVX1 gate3284(.O (I32904), .I (g34708));
INVX1 gate3285(.O (g14833), .I (g11405));
INVX1 gate3286(.O (g19869), .I (g16540));
INVX1 gate3287(.O (g21609), .I (g18008));
INVX1 gate3288(.O (g19960), .I (g17433));
INVX1 gate3289(.O (g23609), .I (g21611));
INVX1 gate3290(.O (g24397), .I (g22908));
INVX1 gate3291(.O (g29339), .I (g28274));
INVX1 gate3292(.O (g12881), .I (g10388));
INVX1 gate3293(.O (g7565), .I (I12046));
INVX1 gate3294(.O (g22903), .I (g20330));
INVX1 gate3295(.O (g13175), .I (g10909));
INVX1 gate3296(.O (g34915), .I (I33137));
INVX1 gate3297(.O (I16593), .I (g10498));
INVX1 gate3298(.O (I25115), .I (g25322));
INVX1 gate3299(.O (g32579), .I (g30735));
INVX1 gate3300(.O (g8068), .I (g3457));
INVX1 gate3301(.O (I13020), .I (g6750));
INVX1 gate3302(.O (I32621), .I (g34335));
INVX1 gate3303(.O (g23312), .I (g21070));
INVX1 gate3304(.O (I31569), .I (g33197));
INVX1 gate3305(.O (I28301), .I (g29042));
INVX1 gate3306(.O (g25219), .I (I24393));
INVX1 gate3307(.O (I27271), .I (g27998));
INVX1 gate3308(.O (g21608), .I (g17955));
INVX1 gate3309(.O (g24062), .I (g19968));
INVX1 gate3310(.O (g17649), .I (I18614));
INVX1 gate3311(.O (g20509), .I (g15277));
INVX1 gate3312(.O (g23608), .I (g21611));
INVX1 gate3313(.O (g34201), .I (I32158));
INVX1 gate3314(.O (g9607), .I (g5046));
INVX1 gate3315(.O (g24509), .I (g22689));
INVX1 gate3316(.O (g32578), .I (g31376));
INVX1 gate3317(.O (g32835), .I (g31710));
INVX1 gate3318(.O (g33695), .I (g33187));
INVX1 gate3319(.O (g34277), .I (I32274));
INVX1 gate3320(.O (g25218), .I (g23949));
INVX1 gate3321(.O (g9962), .I (g6519));
INVX1 gate3322(.O (g11790), .I (I14630));
INVX1 gate3323(.O (g14004), .I (g11149));
INVX1 gate3324(.O (g17648), .I (g15024));
INVX1 gate3325(.O (g20508), .I (g15277));
INVX1 gate3326(.O (g9158), .I (g513));
INVX1 gate3327(.O (g27662), .I (I26296));
INVX1 gate3328(.O (g17491), .I (g12983));
INVX1 gate3329(.O (g22981), .I (g20283));
INVX1 gate3330(.O (g20634), .I (g15373));
INVX1 gate3331(.O (I21029), .I (g15816));
INVX1 gate3332(.O (g21052), .I (g15373));
INVX1 gate3333(.O (g28163), .I (I26682));
INVX1 gate3334(.O (g8677), .I (g4854));
INVX1 gate3335(.O (g25837), .I (g25064));
INVX1 gate3336(.O (g7533), .I (g1306));
INVX1 gate3337(.O (g19709), .I (g16987));
INVX1 gate3338(.O (g32586), .I (g31376));
INVX1 gate3339(.O (I22211), .I (g21463));
INVX1 gate3340(.O (g9506), .I (g5774));
INVX1 gate3341(.O (g17604), .I (I18555));
INVX1 gate3342(.O (g34595), .I (I32693));
INVX1 gate3343(.O (g7697), .I (g4087));
INVX1 gate3344(.O (g10613), .I (g10233));
INVX1 gate3345(.O (g23745), .I (g20900));
INVX1 gate3346(.O (I18504), .I (g5283));
INVX1 gate3347(.O (I22024), .I (g19350));
INVX1 gate3348(.O (g32442), .I (g31213));
INVX1 gate3349(.O (I31814), .I (g33149));
INVX1 gate3350(.O (g19471), .I (g16449));
INVX1 gate3351(.O (g30037), .I (g29121));
INVX1 gate3352(.O (g12890), .I (g10397));
INVX1 gate3353(.O (g16580), .I (I17754));
INVX1 gate3354(.O (g23813), .I (g18997));
INVX1 gate3355(.O (g7596), .I (I12070));
INVX1 gate3356(.O (I31751), .I (g33228));
INVX1 gate3357(.O (I31807), .I (g33149));
INVX1 gate3358(.O (g16223), .I (g13437));
INVX1 gate3359(.O (g10273), .I (I13708));
INVX1 gate3360(.O (g33457), .I (I30989));
INVX1 gate3361(.O (I32062), .I (g33653));
INVX1 gate3362(.O (I12199), .I (g6215));
INVX1 gate3363(.O (g10106), .I (g16));
INVX1 gate3364(.O (g9311), .I (g5523));
INVX1 gate3365(.O (I11743), .I (g4564));
INVX1 gate3366(.O (g22845), .I (g20682));
INVX1 gate3367(.O (I12887), .I (g4216));
INVX1 gate3368(.O (g34984), .I (I33252));
INVX1 gate3369(.O (g32615), .I (g31376));
INVX1 gate3370(.O (I15834), .I (g11164));
INVX1 gate3371(.O (g13209), .I (g10632));
INVX1 gate3372(.O (g8848), .I (g358));
INVX1 gate3373(.O (g20213), .I (g17062));
INVX1 gate3374(.O (I15208), .I (g637));
INVX1 gate3375(.O (g33917), .I (I31779));
INVX1 gate3376(.O (g21184), .I (g15509));
INVX1 gate3377(.O (g34419), .I (g34151));
INVX1 gate3378(.O (g9615), .I (I13236));
INVX1 gate3379(.O (g21674), .I (g16540));
INVX1 gate3380(.O (g10812), .I (I14050));
INVX1 gate3381(.O (g32720), .I (g31710));
INVX1 gate3382(.O (g30155), .I (I28390));
INVX1 gate3383(.O (g8398), .I (I12563));
INVX1 gate3384(.O (g28325), .I (g27463));
INVX1 gate3385(.O (g12779), .I (g9444));
INVX1 gate3386(.O (g22898), .I (g20283));
INVX1 gate3387(.O (g9174), .I (g1205));
INVX1 gate3388(.O (g34418), .I (g34150));
INVX1 gate3389(.O (g17794), .I (g13350));
INVX1 gate3390(.O (g26836), .I (g24866));
INVX1 gate3391(.O (g17845), .I (I18835));
INVX1 gate3392(.O (g9374), .I (g5188));
INVX1 gate3393(.O (g20574), .I (g17847));
INVX1 gate3394(.O (g20452), .I (g17200));
INVX1 gate3395(.O (I15542), .I (g1570));
INVX1 gate3396(.O (g32430), .I (g30984));
INVX1 gate3397(.O (g10033), .I (g655));
INVX1 gate3398(.O (g10371), .I (g6918));
INVX1 gate3399(.O (g32746), .I (g30735));
INVX1 gate3400(.O (g32493), .I (g30735));
INVX1 gate3401(.O (g22719), .I (I22024));
INVX1 gate3402(.O (g24452), .I (g22722));
INVX1 gate3403(.O (I26100), .I (g26365));
INVX1 gate3404(.O (g7936), .I (g1061));
INVX1 gate3405(.O (g9985), .I (g4332));
INVX1 gate3406(.O (g24047), .I (g19919));
INVX1 gate3407(.O (g12778), .I (g9856));
INVX1 gate3408(.O (I18245), .I (g14676));
INVX1 gate3409(.O (I12764), .I (g4194));
INVX1 gate3410(.O (g23732), .I (g18833));
INVX1 gate3411(.O (g8241), .I (g1792));
INVX1 gate3412(.O (I20793), .I (g17694));
INVX1 gate3413(.O (g20912), .I (g15171));
INVX1 gate3414(.O (g19602), .I (g16349));
INVX1 gate3415(.O (g32465), .I (g30825));
INVX1 gate3416(.O (g7117), .I (I11816));
INVX1 gate3417(.O (I18323), .I (g13680));
INVX1 gate3418(.O (g19657), .I (g16349));
INVX1 gate3419(.O (g22718), .I (g20887));
INVX1 gate3420(.O (g16740), .I (g13980));
INVX1 gate3421(.O (I12132), .I (g577));
INVX1 gate3422(.O (g19068), .I (g16031));
INVX1 gate3423(.O (g15169), .I (I17094));
INVX1 gate3424(.O (g28121), .I (g27093));
INVX1 gate3425(.O (g9284), .I (g2161));
INVX1 gate3426(.O (g19375), .I (I19863));
INVX1 gate3427(.O (g10795), .I (g7202));
INVX1 gate3428(.O (I25692), .I (g25689));
INVX1 gate3429(.O (g9239), .I (g5511));
INVX1 gate3430(.O (g33923), .I (I31791));
INVX1 gate3431(.O (g9180), .I (g3719));
INVX1 gate3432(.O (g16186), .I (g13555));
INVX1 gate3433(.O (g16676), .I (I17876));
INVX1 gate3434(.O (g16685), .I (g14038));
INVX1 gate3435(.O (I20690), .I (g15733));
INVX1 gate3436(.O (I29936), .I (g30606));
INVX1 gate3437(.O (I17658), .I (g13394));
INVX1 gate3438(.O (g9380), .I (g5471));
INVX1 gate3439(.O (g12945), .I (g12467));
INVX1 gate3440(.O (g31624), .I (I29218));
INVX1 gate3441(.O (g32806), .I (g31710));
INVX1 gate3442(.O (g20072), .I (g17384));
INVX1 gate3443(.O (g32684), .I (g30673));
INVX1 gate3444(.O (g33688), .I (I31523));
INVX1 gate3445(.O (g29707), .I (g28504));
INVX1 gate3446(.O (g9832), .I (g2399));
INVX1 gate3447(.O (I15073), .I (g10109));
INVX1 gate3448(.O (g19878), .I (g17271));
INVX1 gate3449(.O (g24051), .I (g21127));
INVX1 gate3450(.O (g24072), .I (g20982));
INVX1 gate3451(.O (g34589), .I (I32675));
INVX1 gate3452(.O (g17718), .I (g14776));
INVX1 gate3453(.O (g17521), .I (g14727));
INVX1 gate3454(.O (g16654), .I (g14136));
INVX1 gate3455(.O (g20592), .I (g15277));
INVX1 gate3456(.O (g27998), .I (I26512));
INVX1 gate3457(.O (I16575), .I (g3298));
INVX1 gate3458(.O (g15479), .I (g14895));
INVX1 gate3459(.O (g9853), .I (g5297));
INVX1 gate3460(.O (I15593), .I (g11989));
INVX1 gate3461(.O (g8644), .I (g3352));
INVX1 gate3462(.O (g6989), .I (g4575));
INVX1 gate3463(.O (g9020), .I (g4287));
INVX1 gate3464(.O (g24756), .I (g22763));
INVX1 gate3465(.O (I32452), .I (g34241));
INVX1 gate3466(.O (I12709), .I (g4284));
INVX1 gate3467(.O (g21400), .I (g17847));
INVX1 gate3468(.O (g20780), .I (g15509));
INVX1 gate3469(.O (g7922), .I (g1312));
INVX1 gate3470(.O (g8119), .I (g3727));
INVX1 gate3471(.O (g13530), .I (g12641));
INVX1 gate3472(.O (g23400), .I (g20676));
INVX1 gate3473(.O (g12998), .I (g11829));
INVX1 gate3474(.O (g34836), .I (I33050));
INVX1 gate3475(.O (g13593), .I (g10556));
INVX1 gate3476(.O (g28173), .I (I26693));
INVX1 gate3477(.O (g18929), .I (g16100));
INVX1 gate3478(.O (g32517), .I (g31194));
INVX1 gate3479(.O (g23013), .I (g20330));
INVX1 gate3480(.O (I28572), .I (g28274));
INVX1 gate3481(.O (g12233), .I (g10338));
INVX1 gate3482(.O (I31586), .I (g33149));
INVX1 gate3483(.O (g23214), .I (g20785));
INVX1 gate3484(.O (g11122), .I (g8751));
INVX1 gate3485(.O (I14902), .I (g9821));
INVX1 gate3486(.O (I14301), .I (g8571));
INVX1 gate3487(.O (g12182), .I (I15030));
INVX1 gate3488(.O (g29978), .I (g28927));
INVX1 gate3489(.O (g12672), .I (g10003));
INVX1 gate3490(.O (g7581), .I (g1379));
INVX1 gate3491(.O (g21329), .I (g16577));
INVX1 gate3492(.O (g22926), .I (g20391));
INVX1 gate3493(.O (g25155), .I (g22472));
INVX1 gate3494(.O (g9559), .I (g6077));
INVX1 gate3495(.O (g13565), .I (g11006));
INVX1 gate3496(.O (g6971), .I (I11737));
INVX1 gate3497(.O (g8818), .I (I12808));
INVX1 gate3498(.O (I25005), .I (g24417));
INVX1 gate3499(.O (g14421), .I (I16575));
INVX1 gate3500(.O (I19704), .I (g17653));
INVX1 gate3501(.O (g25266), .I (g22228));
INVX1 gate3502(.O (g25170), .I (g22498));
INVX1 gate3503(.O (g9931), .I (g5763));
INVX1 gate3504(.O (g23539), .I (g21070));
INVX1 gate3505(.O (g17573), .I (g12911));
INVX1 gate3506(.O (g7597), .I (g952));
INVX1 gate3507(.O (g11034), .I (g7611));
INVX1 gate3508(.O (g23005), .I (g20283));
INVX1 gate3509(.O (g13034), .I (g11920));
INVX1 gate3510(.O (g17247), .I (I18259));
INVX1 gate3511(.O (I32051), .I (g33631));
INVX1 gate3512(.O (g30022), .I (g29001));
INVX1 gate3513(.O (g34118), .I (I32051));
INVX1 gate3514(.O (I16606), .I (g3649));
INVX1 gate3515(.O (g15580), .I (g13242));
INVX1 gate3516(.O (g12932), .I (I15550));
INVX1 gate3517(.O (g23538), .I (g20924));
INVX1 gate3518(.O (g34864), .I (g34840));
INVX1 gate3519(.O (I16492), .I (g12430));
INVX1 gate3520(.O (g17389), .I (g14915));
INVX1 gate3521(.O (g17926), .I (I18852));
INVX1 gate3522(.O (g16964), .I (I18120));
INVX1 gate3523(.O (g24152), .I (I23300));
INVX1 gate3524(.O (g19458), .I (I19927));
INVX1 gate3525(.O (g30313), .I (g28843));
INVX1 gate3526(.O (g34749), .I (I32921));
INVX1 gate3527(.O (g17612), .I (g15014));
INVX1 gate3528(.O (g24396), .I (g22885));
INVX1 gate3529(.O (g8211), .I (g2319));
INVX1 gate3530(.O (g29067), .I (I27401));
INVX1 gate3531(.O (g9905), .I (g802));
INVX1 gate3532(.O (g10541), .I (g9407));
INVX1 gate3533(.O (g16423), .I (g14066));
INVX1 gate3534(.O (g27961), .I (g26816));
INVX1 gate3535(.O (g8186), .I (g990));
INVX1 gate3536(.O (g34313), .I (g34086));
INVX1 gate3537(.O (I13552), .I (g121));
INVX1 gate3538(.O (g10473), .I (I13857));
INVX1 gate3539(.O (g17324), .I (I18301));
INVX1 gate3540(.O (g32523), .I (g30825));
INVX1 gate3541(.O (I24128), .I (g23009));
INVX1 gate3542(.O (g31854), .I (g29385));
INVX1 gate3543(.O (g14541), .I (g11405));
INVX1 gate3544(.O (g16216), .I (I17557));
INVX1 gate3545(.O (I29909), .I (g31791));
INVX1 gate3546(.O (I33041), .I (g34772));
INVX1 gate3547(.O (g12897), .I (g10400));
INVX1 gate3548(.O (g13409), .I (I15918));
INVX1 gate3549(.O (g16587), .I (I17763));
INVX1 gate3550(.O (g17777), .I (g14908));
INVX1 gate3551(.O (g25167), .I (I24331));
INVX1 gate3552(.O (g25194), .I (g22763));
INVX1 gate3553(.O (I13779), .I (g6868));
INVX1 gate3554(.O (I26584), .I (g26943));
INVX1 gate3555(.O (g9630), .I (g6527));
INVX1 gate3556(.O (g29150), .I (g27886));
INVX1 gate3557(.O (g34276), .I (g34058));
INVX1 gate3558(.O (g34285), .I (I32284));
INVX1 gate3559(.O (g7995), .I (g153));
INVX1 gate3560(.O (g30305), .I (g28939));
INVX1 gate3561(.O (g11136), .I (I14192));
INVX1 gate3562(.O (g30053), .I (g29121));
INVX1 gate3563(.O (g8026), .I (g3857));
INVX1 gate3564(.O (g25524), .I (g22228));
INVX1 gate3565(.O (I27970), .I (g28803));
INVX1 gate3566(.O (g18827), .I (g16000));
INVX1 gate3567(.O (g34053), .I (g33683));
INVX1 gate3568(.O (g7479), .I (g1008));
INVX1 gate3569(.O (g9300), .I (g5180));
INVX1 gate3570(.O (g10359), .I (g6830));
INVX1 gate3571(.O (I32820), .I (g34474));
INVX1 gate3572(.O (g8426), .I (g3045));
INVX1 gate3573(.O (g32475), .I (g30614));
INVX1 gate3574(.O (g14359), .I (I16515));
INVX1 gate3575(.O (g8170), .I (g3770));
INVX1 gate3576(.O (g7840), .I (g4878));
INVX1 gate3577(.O (g22997), .I (g20391));
INVX1 gate3578(.O (g32727), .I (g31710));
INVX1 gate3579(.O (g10358), .I (g6827));
INVX1 gate3580(.O (g33660), .I (I31494));
INVX1 gate3581(.O (g32863), .I (g31021));
INVX1 gate3582(.O (g29196), .I (g27059));
INVX1 gate3583(.O (I32846), .I (g34502));
INVX1 gate3584(.O (g14535), .I (g12318));
INVX1 gate3585(.O (g24405), .I (g22722));
INVX1 gate3586(.O (g8125), .I (g3869));
INVX1 gate3587(.O (g30036), .I (g29085));
INVX1 gate3588(.O (g14358), .I (I16512));
INVX1 gate3589(.O (g25119), .I (g22384));
INVX1 gate3590(.O (I22819), .I (g19862));
INVX1 gate3591(.O (g8821), .I (I12811));
INVX1 gate3592(.O (g16000), .I (I17425));
INVX1 gate3593(.O (g15740), .I (g13342));
INVX1 gate3594(.O (I25683), .I (g25642));
INVX1 gate3595(.O (I29242), .I (g29313));
INVX1 gate3596(.O (g32437), .I (I29965));
INVX1 gate3597(.O (g14828), .I (I16875));
INVX1 gate3598(.O (g23235), .I (g20785));
INVX1 gate3599(.O (g33456), .I (I30986));
INVX1 gate3600(.O (g10121), .I (g2327));
INVX1 gate3601(.O (g11164), .I (g8085));
INVX1 gate3602(.O (g25118), .I (g22417));
INVX1 gate3603(.O (g26693), .I (g25300));
INVX1 gate3604(.O (g8280), .I (g3443));
INVX1 gate3605(.O (g23683), .I (I22816));
INVX1 gate3606(.O (g15373), .I (I17118));
INVX1 gate3607(.O (g9973), .I (g2112));
INVX1 gate3608(.O (g33916), .I (I31776));
INVX1 gate3609(.O (I22111), .I (g19919));
INVX1 gate3610(.O (g7356), .I (g1802));
INVX1 gate3611(.O (I17819), .I (g3618));
INVX1 gate3612(.O (g16747), .I (g14113));
INVX1 gate3613(.O (g20583), .I (g17873));
INVX1 gate3614(.O (g32703), .I (g30825));
INVX1 gate3615(.O (I12994), .I (g6748));
INVX1 gate3616(.O (I15474), .I (g10364));
INVX1 gate3617(.O (g24020), .I (g20014));
INVX1 gate3618(.O (g19532), .I (g16821));
INVX1 gate3619(.O (g22360), .I (I21849));
INVX1 gate3620(.O (g9040), .I (g499));
INVX1 gate3621(.O (g28648), .I (g27693));
INVX1 gate3622(.O (g18881), .I (I19671));
INVX1 gate3623(.O (I13672), .I (g106));
INVX1 gate3624(.O (g13474), .I (g11048));
INVX1 gate3625(.O (I25882), .I (g25776));
INVX1 gate3626(.O (g20046), .I (g16540));
INVX1 gate3627(.O (g9969), .I (g1682));
INVX1 gate3628(.O (g19783), .I (g16931));
INVX1 gate3629(.O (I17111), .I (g13809));
INVX1 gate3630(.O (g16123), .I (g13530));
INVX1 gate3631(.O (g24046), .I (g21256));
INVX1 gate3632(.O (g17871), .I (I18845));
INVX1 gate3633(.O (g16814), .I (g14058));
INVX1 gate3634(.O (g21414), .I (g17929));
INVX1 gate3635(.O (g32600), .I (g31542));
INVX1 gate3636(.O (g7704), .I (I12167));
INVX1 gate3637(.O (I16663), .I (g10981));
INVX1 gate3638(.O (g23515), .I (g20785));
INVX1 gate3639(.O (g28604), .I (g27759));
INVX1 gate3640(.O (g23882), .I (g19277));
INVX1 gate3641(.O (g23414), .I (I22525));
INVX1 gate3642(.O (g32781), .I (g31376));
INVX1 gate3643(.O (I23099), .I (g20682));
INVX1 gate3644(.O (g31596), .I (I29204));
INVX1 gate3645(.O (g8106), .I (g3133));
INVX1 gate3646(.O (g14173), .I (g12076));
INVX1 gate3647(.O (I23324), .I (g21697));
INVX1 gate3648(.O (g20113), .I (g16826));
INVX1 gate3649(.O (g21407), .I (g15171));
INVX1 gate3650(.O (g31243), .I (g29933));
INVX1 gate3651(.O (I17590), .I (g14591));
INVX1 gate3652(.O (g19353), .I (I19831));
INVX1 gate3653(.O (g24113), .I (g19984));
INVX1 gate3654(.O (I32929), .I (g34649));
INVX1 gate3655(.O (g32952), .I (g30937));
INVX1 gate3656(.O (g19144), .I (g16031));
INVX1 gate3657(.O (g12811), .I (g10319));
INVX1 gate3658(.O (g27971), .I (g26673));
INVX1 gate3659(.O (g8187), .I (g1657));
INVX1 gate3660(.O (g32821), .I (g31021));
INVX1 gate3661(.O (g8387), .I (g3080));
INVX1 gate3662(.O (g25036), .I (g23733));
INVX1 gate3663(.O (I31523), .I (g33187));
INVX1 gate3664(.O (g7163), .I (g4593));
INVX1 gate3665(.O (g29597), .I (g28444));
INVX1 gate3666(.O (g25101), .I (g22384));
INVX1 gate3667(.O (g20105), .I (g17433));
INVX1 gate3668(.O (g24357), .I (g22325));
INVX1 gate3669(.O (g25560), .I (g22550));
INVX1 gate3670(.O (g10029), .I (I13548));
INVX1 gate3671(.O (g8756), .I (g4049));
INVX1 gate3672(.O (g22220), .I (I21802));
INVX1 gate3673(.O (g13303), .I (I15869));
INVX1 gate3674(.O (g24105), .I (g19935));
INVX1 gate3675(.O (I17094), .I (g14331));
INVX1 gate3676(.O (I18031), .I (g13680));
INVX1 gate3677(.O (g29689), .I (I27954));
INVX1 gate3678(.O (g14029), .I (g11283));
INVX1 gate3679(.O (g29923), .I (g28874));
INVX1 gate3680(.O (g25642), .I (I24787));
INVX1 gate3681(.O (g32790), .I (g30825));
INVX1 gate3682(.O (g9648), .I (g2177));
INVX1 gate3683(.O (g32137), .I (g31134));
INVX1 gate3684(.O (g10028), .I (g8));
INVX1 gate3685(.O (g9875), .I (g5747));
INVX1 gate3686(.O (g32516), .I (g31070));
INVX1 gate3687(.O (g31655), .I (I29233));
INVX1 gate3688(.O (I29579), .I (g30565));
INVX1 gate3689(.O (g28262), .I (I26785));
INVX1 gate3690(.O (I24445), .I (g22923));
INVX1 gate3691(.O (g20640), .I (g15426));
INVX1 gate3692(.O (I17801), .I (g14936));
INVX1 gate3693(.O (g20769), .I (g17955));
INVX1 gate3694(.O (g17472), .I (g14656));
INVX1 gate3695(.O (I26406), .I (g26187));
INVX1 gate3696(.O (g12368), .I (I15208));
INVX1 gate3697(.O (I16040), .I (g10430));
INVX1 gate3698(.O (I20499), .I (g16224));
INVX1 gate3699(.O (I12086), .I (g622));
INVX1 gate3700(.O (g33670), .I (I31504));
INVX1 gate3701(.O (I31727), .I (g33076));
INVX1 gate3702(.O (g32873), .I (g30614));
INVX1 gate3703(.O (g8046), .I (g528));
INVX1 gate3704(.O (g25064), .I (I24228));
INVX1 gate3705(.O (g16510), .I (g14008));
INVX1 gate3706(.O (g19364), .I (g15825));
INVX1 gate3707(.O (g20768), .I (g17955));
INVX1 gate3708(.O (g28633), .I (g27687));
INVX1 gate3709(.O (g8514), .I (g4258));
INVX1 gate3710(.O (I19238), .I (g15079));
INVX1 gate3711(.O (g34570), .I (g34392));
INVX1 gate3712(.O (g34712), .I (I32868));
INVX1 gate3713(.O (g21725), .I (I21294));
INVX1 gate3714(.O (g11796), .I (g7985));
INVX1 gate3715(.O (g16579), .I (g13267));
INVX1 gate3716(.O (g33335), .I (I30861));
INVX1 gate3717(.O (g8403), .I (I12568));
INVX1 gate3718(.O (g23759), .I (I22886));
INVX1 gate3719(.O (g13174), .I (g10741));
INVX1 gate3720(.O (I21766), .I (g19620));
INVX1 gate3721(.O (I17695), .I (g14330));
INVX1 gate3722(.O (g26941), .I (I25689));
INVX1 gate3723(.O (g34914), .I (I33134));
INVX1 gate3724(.O (g31839), .I (g29385));
INVX1 gate3725(.O (g33839), .I (I31686));
INVX1 gate3726(.O (I32827), .I (g34477));
INVX1 gate3727(.O (g8345), .I (g3794));
INVX1 gate3728(.O (g8841), .I (I12823));
INVX1 gate3729(.O (I14671), .I (g7717));
INVX1 gate3730(.O (g7157), .I (g5706));
INVX1 gate3731(.O (I12159), .I (g608));
INVX1 gate3732(.O (g22147), .I (g18997));
INVX1 gate3733(.O (g26519), .I (I25380));
INVX1 gate3734(.O (g16578), .I (I17750));
INVX1 gate3735(.O (g15569), .I (I17148));
INVX1 gate3736(.O (g8763), .I (I12749));
INVX1 gate3737(.O (I16564), .I (g10429));
INVX1 gate3738(.O (g23435), .I (g18833));
INVX1 gate3739(.O (g31667), .I (g30142));
INVX1 gate3740(.O (g31838), .I (g29385));
INVX1 gate3741(.O (g23082), .I (g21024));
INVX1 gate3742(.O (g32834), .I (g31672));
INVX1 gate3743(.O (g9839), .I (g2724));
INVX1 gate3744(.O (g30074), .I (g29046));
INVX1 gate3745(.O (g26518), .I (g25233));
INVX1 gate3746(.O (g17591), .I (I18526));
INVX1 gate3747(.O (g12896), .I (g10402));
INVX1 gate3748(.O (g17776), .I (g14905));
INVX1 gate3749(.O (g27011), .I (g25917));
INVX1 gate3750(.O (I27561), .I (g28163));
INVX1 gate3751(.O (g15568), .I (g14984));
INVX1 gate3752(.O (g15747), .I (g13307));
INVX1 gate3753(.O (g25009), .I (g22472));
INVX1 gate3754(.O (I13723), .I (g3167));
INVX1 gate3755(.O (I26004), .I (g26818));
INVX1 gate3756(.O (I18868), .I (g14315));
INVX1 gate3757(.O (I23360), .I (g23360));
INVX1 gate3758(.O (g18945), .I (g16100));
INVX1 gate3759(.O (g30567), .I (g29930));
INVX1 gate3760(.O (I30962), .I (g32021));
INVX1 gate3761(.O (g17147), .I (g14321));
INVX1 gate3762(.O (g22858), .I (g20751));
INVX1 gate3763(.O (g34594), .I (I32690));
INVX1 gate3764(.O (I13149), .I (g6745));
INVX1 gate3765(.O (g17754), .I (g14262));
INVX1 gate3766(.O (I16847), .I (g6329));
INVX1 gate3767(.O (g26935), .I (I25677));
INVX1 gate3768(.O (g25008), .I (g22432));
INVX1 gate3769(.O (g32542), .I (g31554));
INVX1 gate3770(.O (g8107), .I (g3179));
INVX1 gate3771(.O (I32803), .I (g34584));
INVX1 gate3772(.O (I25399), .I (g24489));
INVX1 gate3773(.O (g31487), .I (I29149));
INVX1 gate3774(.O (g32021), .I (I29579));
INVX1 gate3775(.O (g32453), .I (I29981));
INVX1 gate3776(.O (I29720), .I (g30931));
INVX1 gate3777(.O (g11192), .I (g8038));
INVX1 gate3778(.O (g22151), .I (I21734));
INVX1 gate3779(.O (I11620), .I (g1));
INVX1 gate3780(.O (I21162), .I (g17292));
INVX1 gate3781(.O (I12144), .I (g554));
INVX1 gate3782(.O (I12823), .I (g4311));
INVX1 gate3783(.O (I18709), .I (g6668));
INVX1 gate3784(.O (g20662), .I (g15171));
INVX1 gate3785(.O (g21399), .I (g15224));
INVX1 gate3786(.O (g23849), .I (g19277));
INVX1 gate3787(.O (g22996), .I (g20330));
INVX1 gate3788(.O (g23940), .I (g19074));
INVX1 gate3789(.O (g25892), .I (g24528));
INVX1 gate3790(.O (I20753), .I (g16677));
INVX1 gate3791(.O (I15663), .I (g5308));
INVX1 gate3792(.O (g23399), .I (g21514));
INVX1 gate3793(.O (g32726), .I (g31672));
INVX1 gate3794(.O (g32913), .I (g30825));
INVX1 gate3795(.O (g24027), .I (g20014));
INVX1 gate3796(.O (I18259), .I (g12946));
INVX1 gate3797(.O (g9618), .I (g5794));
INVX1 gate3798(.O (g11663), .I (g6905));
INVX1 gate3799(.O (g16615), .I (I17801));
INVX1 gate3800(.O (g22844), .I (g21163));
INVX1 gate3801(.O (g13522), .I (g10981));
INVX1 gate3802(.O (g34941), .I (g34926));
INVX1 gate3803(.O (g13663), .I (g10971));
INVX1 gate3804(.O (g21398), .I (g18008));
INVX1 gate3805(.O (g23848), .I (g19210));
INVX1 gate3806(.O (g25555), .I (g22550));
INVX1 gate3807(.O (g32614), .I (g31542));
INVX1 gate3808(.O (g7626), .I (I12112));
INVX1 gate3809(.O (I12336), .I (g52));
INVX1 gate3810(.O (g23398), .I (g21468));
INVX1 gate3811(.O (I32881), .I (g34688));
INVX1 gate3812(.O (g8858), .I (g671));
INVX1 gate3813(.O (g33443), .I (I30971));
INVX1 gate3814(.O (g16720), .I (g14234));
INVX1 gate3815(.O (g9282), .I (g723));
INVX1 gate3816(.O (g34675), .I (I32809));
INVX1 gate3817(.O (I20650), .I (g17010));
INVX1 gate3818(.O (g23652), .I (I22785));
INVX1 gate3819(.O (g32607), .I (g31542));
INVX1 gate3820(.O (g8016), .I (g3391));
INVX1 gate3821(.O (g10981), .I (I14119));
INVX1 gate3822(.O (g8757), .I (I12746));
INVX1 gate3823(.O (g32905), .I (g30825));
INVX1 gate3824(.O (g14563), .I (I16676));
INVX1 gate3825(.O (g8416), .I (I12580));
INVX1 gate3826(.O (g27112), .I (g26793));
INVX1 gate3827(.O (g20710), .I (g15509));
INVX1 gate3828(.O (g16746), .I (g14258));
INVX1 gate3829(.O (I20529), .I (g16309));
INVX1 gate3830(.O (I21911), .I (g21278));
INVX1 gate3831(.O (g17844), .I (I18832));
INVX1 gate3832(.O (g20552), .I (g17847));
INVX1 gate3833(.O (g32530), .I (g30825));
INVX1 gate3834(.O (g9693), .I (g1886));
INVX1 gate3835(.O (g13483), .I (g11270));
INVX1 gate3836(.O (I33264), .I (g34978));
INVX1 gate3837(.O (I15862), .I (g11215));
INVX1 gate3838(.O (g17367), .I (I18320));
INVX1 gate3839(.O (g32593), .I (g31542));
INVX1 gate3840(.O (g18932), .I (g16136));
INVX1 gate3841(.O (g6985), .I (g4669));
INVX1 gate3842(.O (I33137), .I (g34884));
INVX1 gate3843(.O (g20204), .I (g16578));
INVX1 gate3844(.O (g19687), .I (g17096));
INVX1 gate3845(.O (I21246), .I (g16540));
INVX1 gate3846(.O (g24003), .I (g21514));
INVX1 gate3847(.O (g23263), .I (I22366));
INVX1 gate3848(.O (I12631), .I (g1242));
INVX1 gate3849(.O (g8522), .I (g298));
INVX1 gate3850(.O (g20779), .I (g15509));
INVX1 gate3851(.O (g22319), .I (I21831));
INVX1 gate3852(.O (g12378), .I (g9417));
INVX1 gate3853(.O (g34935), .I (I33189));
INVX1 gate3854(.O (g23332), .I (g20785));
INVX1 gate3855(.O (g32565), .I (g30735));
INVX1 gate3856(.O (g32464), .I (g30735));
INVX1 gate3857(.O (g25239), .I (g23972));
INVX1 gate3858(.O (g19954), .I (g16540));
INVX1 gate3859(.O (g11949), .I (I14773));
INVX1 gate3860(.O (I24393), .I (g23453));
INVX1 gate3861(.O (g19374), .I (g16047));
INVX1 gate3862(.O (g20778), .I (g15224));
INVX1 gate3863(.O (g34883), .I (g34852));
INVX1 gate3864(.O (g10794), .I (g8470));
INVX1 gate3865(.O (g9555), .I (I13206));
INVX1 gate3866(.O (g18897), .I (g15509));
INVX1 gate3867(.O (I15536), .I (g1227));
INVX1 gate3868(.O (g10395), .I (g6995));
INVX1 gate3869(.O (g22227), .I (g19801));
INVX1 gate3870(.O (g24778), .I (g23286));
INVX1 gate3871(.O (g9804), .I (g5456));
INVX1 gate3872(.O (g10262), .I (g586));
INVX1 gate3873(.O (g24081), .I (g21209));
INVX1 gate3874(.O (g21406), .I (g17955));
INVX1 gate3875(.O (g16684), .I (g14223));
INVX1 gate3876(.O (g11948), .I (g10224));
INVX1 gate3877(.O (I21776), .I (g21308));
INVX1 gate3878(.O (I15702), .I (g12217));
INVX1 gate3879(.O (g14262), .I (g10838));
INVX1 gate3880(.O (g12944), .I (g12659));
INVX1 gate3881(.O (I18810), .I (g13716));
INVX1 gate3882(.O (g23406), .I (g20330));
INVX1 gate3883(.O (g9792), .I (g5401));
INVX1 gate3884(.O (g32641), .I (g30614));
INVX1 gate3885(.O (g6832), .I (I11665));
INVX1 gate3886(.O (g32797), .I (g30825));
INVX1 gate3887(.O (g23962), .I (g19147));
INVX1 gate3888(.O (g31815), .I (g29385));
INVX1 gate3889(.O (g23361), .I (I22464));
INVX1 gate3890(.O (g28032), .I (g26365));
INVX1 gate3891(.O (I32482), .I (g34304));
INVX1 gate3892(.O (g11702), .I (g6928));
INVX1 gate3893(.O (g7778), .I (g1339));
INVX1 gate3894(.O (g15579), .I (I17159));
INVX1 gate3895(.O (g31601), .I (I29207));
INVX1 gate3896(.O (g8654), .I (g1087));
INVX1 gate3897(.O (I16452), .I (g11182));
INVX1 gate3898(.O (I18879), .I (g13267));
INVX1 gate3899(.O (g9621), .I (g6423));
INVX1 gate3900(.O (g10191), .I (g6386));
INVX1 gate3901(.O (g23500), .I (g20924));
INVX1 gate3902(.O (g24356), .I (g22594));
INVX1 gate3903(.O (g13621), .I (g10573));
INVX1 gate3904(.O (g21049), .I (g17433));
INVX1 gate3905(.O (I11896), .I (g4446));
INVX1 gate3906(.O (g25185), .I (g22228));
INVX1 gate3907(.O (g17059), .I (I18151));
INVX1 gate3908(.O (g20380), .I (g17955));
INVX1 gate3909(.O (g26083), .I (g24809));
INVX1 gate3910(.O (g14191), .I (g12381));
INVX1 gate3911(.O (g30729), .I (I28883));
INVX1 gate3912(.O (I15564), .I (g11949));
INVX1 gate3913(.O (g25092), .I (g23666));
INVX1 gate3914(.O (g24999), .I (g23626));
INVX1 gate3915(.O (g26284), .I (g24875));
INVX1 gate3916(.O (I18337), .I (g1422));
INVX1 gate3917(.O (g34501), .I (g34400));
INVX1 gate3918(.O (g27730), .I (g26424));
INVX1 gate3919(.O (g10521), .I (I13889));
INVX1 gate3920(.O (g12857), .I (I15474));
INVX1 gate3921(.O (I19348), .I (g15084));
INVX1 gate3922(.O (g21048), .I (g17533));
INVX1 gate3923(.O (g25154), .I (g22457));
INVX1 gate3924(.O (g20090), .I (g17433));
INVX1 gate3925(.O (g17058), .I (I18148));
INVX1 gate3926(.O (g32635), .I (g31542));
INVX1 gate3927(.O (g8880), .I (I12861));
INVX1 gate3928(.O (g31937), .I (g30991));
INVX1 gate3929(.O (g8595), .I (I12666));
INVX1 gate3930(.O (g24090), .I (g19935));
INVX1 gate3931(.O (g19489), .I (g16449));
INVX1 gate3932(.O (g20233), .I (g17873));
INVX1 gate3933(.O (g33937), .I (I31823));
INVX1 gate3934(.O (g12793), .I (g10287));
INVX1 gate3935(.O (I11716), .I (g4054));
INVX1 gate3936(.O (g20182), .I (g16897));
INVX1 gate3937(.O (g20651), .I (g15483));
INVX1 gate3938(.O (g20672), .I (g15277));
INVX1 gate3939(.O (I17876), .I (g13070));
INVX1 gate3940(.O (g23004), .I (g20283));
INVX1 gate3941(.O (I27495), .I (g27961));
INVX1 gate3942(.O (g7475), .I (g896));
INVX1 gate3943(.O (g21221), .I (g15680));
INVX1 gate3944(.O (g24182), .I (I23390));
INVX1 gate3945(.O (g19559), .I (g16129));
INVX1 gate3946(.O (g23221), .I (g20785));
INVX1 gate3947(.O (I14644), .I (g7717));
INVX1 gate3948(.O (g11183), .I (g8135));
INVX1 gate3949(.O (g29942), .I (g28867));
INVX1 gate3950(.O (g22957), .I (I22143));
INVX1 gate3951(.O (g31791), .I (I29363));
INVX1 gate3952(.O (g7627), .I (g4311));
INVX1 gate3953(.O (g19558), .I (g15938));
INVX1 gate3954(.O (g6905), .I (I11708));
INVX1 gate3955(.O (g16523), .I (g14041));
INVX1 gate3956(.O (g8612), .I (g2775));
INVX1 gate3957(.O (g23613), .I (I22748));
INVX1 gate3958(.O (g9518), .I (g6219));
INVX1 gate3959(.O (g15615), .I (I17181));
INVX1 gate3960(.O (I17763), .I (g13191));
INVX1 gate3961(.O (I31607), .I (g33164));
INVX1 gate3962(.O (g13062), .I (g10981));
INVX1 gate3963(.O (g7526), .I (I12013));
INVX1 gate3964(.O (g7998), .I (g392));
INVX1 gate3965(.O (g11509), .I (g7632));
INVX1 gate3966(.O (g22146), .I (g18997));
INVX1 gate3967(.O (g26653), .I (g25337));
INVX1 gate3968(.O (g20513), .I (g18065));
INVX1 gate3969(.O (g17301), .I (g14454));
INVX1 gate3970(.O (g20449), .I (g15277));
INVX1 gate3971(.O (g28162), .I (I26679));
INVX1 gate3972(.O (g10389), .I (g6986));
INVX1 gate3973(.O (g32891), .I (g30825));
INVX1 gate3974(.O (I15872), .I (g11236));
INVX1 gate3975(.O (g13933), .I (g11419));
INVX1 gate3976(.O (g23947), .I (g19210));
INVX1 gate3977(.O (g31479), .I (I29139));
INVX1 gate3978(.O (g31666), .I (I29248));
INVX1 gate3979(.O (I27954), .I (g28803));
INVX1 gate3980(.O (g18097), .I (I18897));
INVX1 gate3981(.O (g21273), .I (I21006));
INVX1 gate3982(.O (g17120), .I (g14262));
INVX1 gate3983(.O (g19544), .I (g16349));
INVX1 gate3984(.O (g23273), .I (g21070));
INVX1 gate3985(.O (g19865), .I (g15885));
INVX1 gate3986(.O (g17739), .I (I18728));
INVX1 gate3987(.O (g10612), .I (g10233));
INVX1 gate3988(.O (g11872), .I (I14684));
INVX1 gate3989(.O (g23605), .I (g20739));
INVX1 gate3990(.O (g9776), .I (g5073));
INVX1 gate3991(.O (g10099), .I (g6682));
INVX1 gate3992(.O (g15746), .I (g13121));
INVX1 gate3993(.O (g16475), .I (g14107));
INVX1 gate3994(.O (g20448), .I (g15509));
INVX1 gate3995(.O (g34304), .I (I32309));
INVX1 gate3996(.O (I12954), .I (g4358));
INVX1 gate3997(.O (g10388), .I (g6983));
INVX1 gate3998(.O (I32651), .I (g34375));
INVX1 gate3999(.O (g32575), .I (g31170));
INVX1 gate4000(.O (g32474), .I (g31194));
INVX1 gate4001(.O (g19713), .I (g16816));
INVX1 gate4002(.O (g7439), .I (g6351));
INVX1 gate4003(.O (g29930), .I (I28162));
INVX1 gate4004(.O (g22698), .I (I22009));
INVX1 gate4005(.O (g29993), .I (g29018));
INVX1 gate4006(.O (g16727), .I (g14454));
INVX1 gate4007(.O (g17738), .I (g14813));
INVX1 gate4008(.O (g17645), .I (g15018));
INVX1 gate4009(.O (g20505), .I (g15426));
INVX1 gate4010(.O (g21463), .I (g15588));
INVX1 gate4011(.O (g23812), .I (g18997));
INVX1 gate4012(.O (g32711), .I (g31070));
INVX1 gate4013(.O (g8130), .I (g4515));
INVX1 gate4014(.O (g14701), .I (g12351));
INVX1 gate4015(.O (I17456), .I (g13680));
INVX1 gate4016(.O (I23318), .I (g21689));
INVX1 gate4017(.O (g8542), .I (I12644));
INVX1 gate4018(.O (g24505), .I (g22689));
INVX1 gate4019(.O (g8330), .I (g2587));
INVX1 gate4020(.O (g24404), .I (g22908));
INVX1 gate4021(.O (g10272), .I (I13705));
INVX1 gate4022(.O (g9965), .I (g127));
INVX1 gate4023(.O (g29965), .I (g28903));
INVX1 gate4024(.O (I33034), .I (g34769));
INVX1 gate4025(.O (g14251), .I (g12308));
INVX1 gate4026(.O (I17916), .I (g13087));
INVX1 gate4027(.O (g20026), .I (g17271));
INVX1 gate4028(.O (g32537), .I (g30825));
INVX1 gate4029(.O (I18078), .I (g13350));
INVX1 gate4030(.O (g20212), .I (g17194));
INVX1 gate4031(.O (g23234), .I (g20375));
INVX1 gate4032(.O (g24026), .I (g19919));
INVX1 gate4033(.O (g9264), .I (g5396));
INVX1 gate4034(.O (g15806), .I (I17302));
INVX1 gate4035(.O (I21058), .I (g17747));
INVX1 gate4036(.O (g25438), .I (g22763));
INVX1 gate4037(.O (g6973), .I (I11743));
INVX1 gate4038(.O (I17314), .I (g14078));
INVX1 gate4039(.O (I32449), .I (g34127));
INVX1 gate4040(.O (g19679), .I (g16782));
INVX1 gate4041(.O (I18086), .I (g13856));
INVX1 gate4042(.O (g27245), .I (g26209));
INVX1 gate4043(.O (g34653), .I (I32763));
INVX1 gate4044(.O (g9360), .I (g3372));
INVX1 gate4045(.O (g9933), .I (g5759));
INVX1 gate4046(.O (g32606), .I (g30673));
INVX1 gate4047(.O (g10032), .I (g562));
INVX1 gate4048(.O (I29236), .I (g29498));
INVX1 gate4049(.O (g32492), .I (g31376));
INVX1 gate4050(.O (g19678), .I (g16752));
INVX1 gate4051(.O (I15205), .I (g10139));
INVX1 gate4052(.O (g14032), .I (g11048));
INVX1 gate4053(.O (g10140), .I (g19));
INVX1 gate4054(.O (g29210), .I (I27546));
INVX1 gate4055(.O (g9050), .I (g1087));
INVX1 gate4056(.O (g17427), .I (I18364));
INVX1 gate4057(.O (I13802), .I (g6971));
INVX1 gate4058(.O (g13574), .I (I16024));
INVX1 gate4059(.O (I25514), .I (g25073));
INVX1 gate4060(.O (I13857), .I (g9780));
INVX1 gate4061(.O (g17366), .I (g14454));
INVX1 gate4062(.O (g7952), .I (g3774));
INVX1 gate4063(.O (g25083), .I (g23782));
INVX1 gate4064(.O (g25348), .I (g22763));
INVX1 gate4065(.O (g9450), .I (g5817));
INVX1 gate4066(.O (I14450), .I (g4191));
INVX1 gate4067(.O (g16600), .I (I17780));
INVX1 gate4068(.O (g19686), .I (g17062));
INVX1 gate4069(.O (g25284), .I (I24474));
INVX1 gate4070(.O (g21514), .I (I21189));
INVX1 gate4071(.O (I11793), .I (g6049));
INVX1 gate4072(.O (g11912), .I (g8989));
INVX1 gate4073(.O (g26576), .I (I25399));
INVX1 gate4074(.O (I26682), .I (g27774));
INVX1 gate4075(.O (g28147), .I (I26654));
INVX1 gate4076(.O (I27558), .I (g28155));
INVX1 gate4077(.O (g32750), .I (g30937));
INVX1 gate4078(.O (I12016), .I (g772));
INVX1 gate4079(.O (I18125), .I (g13191));
INVX1 gate4080(.O (g10061), .I (I13581));
INVX1 gate4081(.O (g13311), .I (I15878));
INVX1 gate4082(.O (g28754), .I (I27238));
INVX1 gate4083(.O (g32381), .I (I29909));
INVX1 gate4084(.O (g7616), .I (I12086));
INVX1 gate4085(.O (I19484), .I (g15122));
INVX1 gate4086(.O (g23507), .I (g21562));
INVX1 gate4087(.O (g34852), .I (g34845));
INVX1 gate4088(.O (g20433), .I (g17929));
INVX1 gate4089(.O (g25566), .I (g22550));
INVX1 gate4090(.O (g18896), .I (g16031));
INVX1 gate4091(.O (g24149), .I (g19338));
INVX1 gate4092(.O (g20387), .I (g15426));
INVX1 gate4093(.O (g28370), .I (g27528));
INVX1 gate4094(.O (I28866), .I (g29730));
INVX1 gate4095(.O (I22180), .I (g21366));
INVX1 gate4096(.O (g16821), .I (I18031));
INVX1 gate4097(.O (g21421), .I (g15171));
INVX1 gate4098(.O (g27737), .I (g26718));
INVX1 gate4099(.O (I12893), .I (g4226));
INVX1 gate4100(.O (g7004), .I (I11777));
INVX1 gate4101(.O (g9379), .I (g5424));
INVX1 gate4102(.O (g23421), .I (g21562));
INVX1 gate4103(.O (g13051), .I (g11964));
INVX1 gate4104(.O (g20097), .I (g17691));
INVX1 gate4105(.O (g32796), .I (g31376));
INVX1 gate4106(.O (g7527), .I (I12016));
INVX1 gate4107(.O (I33164), .I (g34894));
INVX1 gate4108(.O (g24097), .I (g19935));
INVX1 gate4109(.O (g26608), .I (g25334));
INVX1 gate4110(.O (g11592), .I (I14537));
INVX1 gate4111(.O (g20104), .I (g17433));
INVX1 gate4112(.O (g7647), .I (I12132));
INVX1 gate4113(.O (g34664), .I (I32782));
INVX1 gate4114(.O (I27713), .I (g28224));
INVX1 gate4115(.O (I13548), .I (g94));
INVX1 gate4116(.O (g10360), .I (g6836));
INVX1 gate4117(.O (g23012), .I (g20330));
INVX1 gate4118(.O (g24104), .I (g19890));
INVX1 gate4119(.O (g17226), .I (I18252));
INVX1 gate4120(.O (g25139), .I (g22472));
INVX1 gate4121(.O (g17715), .I (I18700));
INVX1 gate4122(.O (g6875), .I (I11697));
INVX1 gate4123(.O (g9777), .I (g5112));
INVX1 gate4124(.O (g17481), .I (g15005));
INVX1 gate4125(.O (I25541), .I (g25180));
INVX1 gate4126(.O (g32840), .I (g30825));
INVX1 gate4127(.O (I28597), .I (g29374));
INVX1 gate4128(.O (g28367), .I (I26880));
INVX1 gate4129(.O (I31474), .I (g33212));
INVX1 gate4130(.O (g24971), .I (g23590));
INVX1 gate4131(.O (g27880), .I (I26427));
INVX1 gate4132(.O (g25138), .I (g22472));
INVX1 gate4133(.O (g34576), .I (I32654));
INVX1 gate4134(.O (g16873), .I (I18063));
INVX1 gate4135(.O (g23541), .I (g21514));
INVX1 gate4136(.O (g31800), .I (g29385));
INVX1 gate4137(.O (g12995), .I (g11820));
INVX1 gate4138(.O (g7503), .I (g1351));
INVX1 gate4139(.O (g7970), .I (g4688));
INVX1 gate4140(.O (g13350), .I (I15906));
INVX1 gate4141(.O (g23473), .I (g20785));
INVX1 gate4142(.O (g33800), .I (I31642));
INVX1 gate4143(.O (g8056), .I (g1246));
INVX1 gate4144(.O (I13317), .I (g6144));
INVX1 gate4145(.O (g11820), .I (I14644));
INVX1 gate4146(.O (g33936), .I (I31820));
INVX1 gate4147(.O (g8456), .I (g56));
INVX1 gate4148(.O (g12880), .I (g10387));
INVX1 gate4149(.O (I22131), .I (g19984));
INVX1 gate4150(.O (I24078), .I (g22360));
INVX1 gate4151(.O (g23789), .I (g21308));
INVX1 gate4152(.O (I17839), .I (g13412));
INVX1 gate4153(.O (g32192), .I (g31262));
INVX1 gate4154(.O (I33109), .I (g34851));
INVX1 gate4155(.O (I15846), .I (g11183));
INVX1 gate4156(.O (I16357), .I (g884));
INVX1 gate4157(.O (I25359), .I (g24715));
INVX1 gate4158(.O (I19799), .I (g17817));
INVX1 gate4159(.O (g30312), .I (g28970));
INVX1 gate4160(.O (I12189), .I (g5869));
INVX1 gate4161(.O (I19813), .I (g17952));
INVX1 gate4162(.O (g24368), .I (g22228));
INVX1 gate4163(.O (g21724), .I (I21291));
INVX1 gate4164(.O (g23788), .I (g18997));
INVX1 gate4165(.O (g8155), .I (g3380));
INVX1 gate4166(.O (g34312), .I (g34098));
INVX1 gate4167(.O (g26973), .I (g26105));
INVX1 gate4168(.O (g34200), .I (g33895));
INVX1 gate4169(.O (g7224), .I (g4601));
INVX1 gate4170(.O (g32522), .I (g30735));
INVX1 gate4171(.O (g23359), .I (I22458));
INVX1 gate4172(.O (g32663), .I (g30673));
INVX1 gate4173(.O (g8355), .I (I12534));
INVX1 gate4174(.O (g8851), .I (g590));
INVX1 gate4175(.O (I13057), .I (g112));
INVX1 gate4176(.O (g14451), .I (I16606));
INVX1 gate4177(.O (I23366), .I (g23321));
INVX1 gate4178(.O (I18364), .I (g13009));
INVX1 gate4179(.O (I22619), .I (g21193));
INVX1 gate4180(.O (I17131), .I (g14384));
INVX1 gate4181(.O (I22502), .I (g19376));
INVX1 gate4182(.O (g22980), .I (I22153));
INVX1 gate4183(.O (g21434), .I (g17248));
INVX1 gate4184(.O (I22557), .I (g20695));
INVX1 gate4185(.O (g21358), .I (g16307));
INVX1 gate4186(.O (g6839), .I (g1858));
INVX1 gate4187(.O (g23434), .I (g21611));
INVX1 gate4188(.O (g24850), .I (I24022));
INVX1 gate4189(.O (g30052), .I (g29018));
INVX1 gate4190(.O (I19674), .I (g15932));
INVX1 gate4191(.O (g8964), .I (g4269));
INVX1 gate4192(.O (I29913), .I (g30605));
INVX1 gate4193(.O (g27831), .I (I26406));
INVX1 gate4194(.O (I11626), .I (g31));
INVX1 gate4195(.O (g11413), .I (g9100));
INVX1 gate4196(.O (g34921), .I (I33155));
INVX1 gate4197(.O (g13413), .I (g11737));
INVX1 gate4198(.O (g34052), .I (g33635));
INVX1 gate4199(.O (g23946), .I (g19210));
INVX1 gate4200(.O (g24133), .I (g19935));
INVX1 gate4201(.O (g29169), .I (g27886));
INVX1 gate4202(.O (g18096), .I (I18894));
INVX1 gate4203(.O (g18944), .I (g15938));
INVX1 gate4204(.O (g20229), .I (g17015));
INVX1 gate4205(.O (g32483), .I (g30673));
INVX1 gate4206(.O (g19617), .I (g16349));
INVX1 gate4207(.O (g19470), .I (g16000));
INVX1 gate4208(.O (g22181), .I (g19277));
INVX1 gate4209(.O (g11691), .I (I14570));
INVX1 gate4210(.O (g19915), .I (g16349));
INVX1 gate4211(.O (g12831), .I (g9569));
INVX1 gate4212(.O (g26732), .I (g25389));
INVX1 gate4213(.O (I16803), .I (g6369));
INVX1 gate4214(.O (I12030), .I (g595));
INVX1 gate4215(.O (I17557), .I (g14510));
INVX1 gate4216(.O (g9541), .I (g2012));
INVX1 gate4217(.O (g32553), .I (g31170));
INVX1 gate4218(.O (g32862), .I (g30825));
INVX1 gate4219(.O (g7617), .I (I12089));
INVX1 gate4220(.O (g16726), .I (g14454));
INVX1 gate4221(.O (I26649), .I (g27675));
INVX1 gate4222(.O (g34813), .I (I33027));
INVX1 gate4223(.O (g10776), .I (I14033));
INVX1 gate4224(.O (g19277), .I (I19813));
INVX1 gate4225(.O (g32949), .I (g30825));
INVX1 gate4226(.O (g9332), .I (g64));
INVX1 gate4227(.O (g14591), .I (I16709));
INVX1 gate4228(.O (g14785), .I (g12629));
INVX1 gate4229(.O (I21226), .I (g16540));
INVX1 gate4230(.O (I22286), .I (g19446));
INVX1 gate4231(.O (g7516), .I (I12003));
INVX1 gate4232(.O (g21682), .I (g16540));
INVX1 gate4233(.O (I18224), .I (g13793));
INVX1 gate4234(.O (g9680), .I (I13276));
INVX1 gate4235(.O (g9153), .I (I12991));
INVX1 gate4236(.O (g10147), .I (g728));
INVX1 gate4237(.O (g20716), .I (g15277));
INVX1 gate4238(.O (g27989), .I (g26759));
INVX1 gate4239(.O (g29217), .I (I27567));
INVX1 gate4240(.O (g34973), .I (I33235));
INVX1 gate4241(.O (g25554), .I (g22550));
INVX1 gate4242(.O (I15929), .I (g10430));
INVX1 gate4243(.O (I18571), .I (g13074));
INVX1 gate4244(.O (g21291), .I (g16620));
INVX1 gate4245(.O (g32536), .I (g31376));
INVX1 gate4246(.O (g14147), .I (I16357));
INVX1 gate4247(.O (g30184), .I (g28144));
INVX1 gate4248(.O (I31796), .I (g33176));
INVX1 gate4249(.O (g10355), .I (g6816));
INVX1 gate4250(.O (g32948), .I (g30735));
INVX1 gate4251(.O (g23291), .I (g21070));
INVX1 gate4252(.O (g16607), .I (g13960));
INVX1 gate4253(.O (g19494), .I (g16349));
INVX1 gate4254(.O (g11929), .I (I14745));
INVX1 gate4255(.O (I11737), .I (g4467));
INVX1 gate4256(.O (g34674), .I (I32806));
INVX1 gate4257(.O (g8279), .I (I12487));
INVX1 gate4258(.O (g16320), .I (g14454));
INVX1 gate4259(.O (g20582), .I (g17873));
INVX1 gate4260(.O (g32702), .I (g30735));
INVX1 gate4261(.O (g9744), .I (g6486));
INVX1 gate4262(.O (g10370), .I (g7095));
INVX1 gate4263(.O (g31000), .I (g29737));
INVX1 gate4264(.O (g32757), .I (g30937));
INVX1 gate4265(.O (g32904), .I (g30735));
INVX1 gate4266(.O (g6988), .I (g4765));
INVX1 gate4267(.O (I14866), .I (g9748));
INVX1 gate4268(.O (g16530), .I (g14454));
INVX1 gate4269(.O (g26400), .I (I25351));
INVX1 gate4270(.O (g11928), .I (I14742));
INVX1 gate4271(.O (g25115), .I (I24281));
INVX1 gate4272(.O (g13583), .I (I16028));
INVX1 gate4273(.O (g32621), .I (g31542));
INVX1 gate4274(.O (g8872), .I (g4258));
INVX1 gate4275(.O (g22520), .I (g19801));
INVX1 gate4276(.O (I22601), .I (g21127));
INVX1 gate4277(.O (g10151), .I (g1992));
INVX1 gate4278(.O (g28120), .I (g27108));
INVX1 gate4279(.O (I32228), .I (g34122));
INVX1 gate4280(.O (I11697), .I (g3352));
INVX1 gate4281(.O (g10172), .I (g6459));
INVX1 gate4282(.O (g20627), .I (g17433));
INVX1 gate4283(.O (I12837), .I (g4222));
INVX1 gate4284(.O (g7892), .I (g4801));
INVX1 gate4285(.O (g34934), .I (g34918));
INVX1 gate4286(.O (g9558), .I (g5841));
INVX1 gate4287(.O (g20379), .I (g17821));
INVX1 gate4288(.O (g8057), .I (g3068));
INVX1 gate4289(.O (g32564), .I (g31376));
INVX1 gate4290(.O (I13995), .I (g8744));
INVX1 gate4291(.O (g24379), .I (g22550));
INVX1 gate4292(.O (g8457), .I (g225));
INVX1 gate4293(.O (g8989), .I (I12935));
INVX1 gate4294(.O (g19352), .I (g15758));
INVX1 gate4295(.O (g22546), .I (I21918));
INVX1 gate4296(.O (g23760), .I (I22889));
INVX1 gate4297(.O (g20050), .I (I20321));
INVX1 gate4298(.O (g23029), .I (g20453));
INVX1 gate4299(.O (g6804), .I (g490));
INVX1 gate4300(.O (g24112), .I (g19935));
INVX1 gate4301(.O (g10367), .I (g6870));
INVX1 gate4302(.O (g10394), .I (g6994));
INVX1 gate4303(.O (I25028), .I (g24484));
INVX1 gate4304(.O (g24050), .I (g20841));
INVX1 gate4305(.O (g9901), .I (g84));
INVX1 gate4306(.O (g34692), .I (I32846));
INVX1 gate4307(.O (I22143), .I (g20189));
INVX1 gate4308(.O (I21784), .I (g19638));
INVX1 gate4309(.O (g23506), .I (g21514));
INVX1 gate4310(.O (g23028), .I (g20391));
INVX1 gate4311(.O (I18752), .I (g6358));
INVX1 gate4312(.O (I28480), .I (g28652));
INVX1 gate4313(.O (g31814), .I (g29385));
INVX1 gate4314(.O (g32673), .I (g31376));
INVX1 gate4315(.O (g32847), .I (g30735));
INVX1 gate4316(.O (g20386), .I (g15224));
INVX1 gate4317(.O (I21297), .I (g18597));
INVX1 gate4318(.O (g8971), .I (I12927));
INVX1 gate4319(.O (g22860), .I (g20000));
INVX1 gate4320(.O (g24386), .I (g22594));
INVX1 gate4321(.O (g20603), .I (g17873));
INVX1 gate4322(.O (g9511), .I (g5881));
INVX1 gate4323(.O (g27736), .I (I26356));
INVX1 gate4324(.O (g7738), .I (I12176));
INVX1 gate4325(.O (g31807), .I (g29385));
INVX1 gate4326(.O (g8686), .I (g2819));
INVX1 gate4327(.O (g13302), .I (g12321));
INVX1 gate4328(.O (g20096), .I (g16782));
INVX1 gate4329(.O (g24603), .I (g23108));
INVX1 gate4330(.O (g33772), .I (I31622));
INVX1 gate4331(.O (g7991), .I (g4878));
INVX1 gate4332(.O (I23354), .I (g23277));
INVX1 gate4333(.O (g24096), .I (g19890));
INVX1 gate4334(.O (g29922), .I (g28837));
INVX1 gate4335(.O (g34400), .I (g34142));
INVX1 gate4336(.O (g7244), .I (g4408));
INVX1 gate4337(.O (g12887), .I (g10394));
INVX1 gate4338(.O (g10420), .I (g9239));
INVX1 gate4339(.O (I17143), .I (g14412));
INVX1 gate4340(.O (g22497), .I (g19513));
INVX1 gate4341(.O (g25184), .I (g22763));
INVX1 gate4342(.O (g32509), .I (g31070));
INVX1 gate4343(.O (g31639), .I (I29225));
INVX1 gate4344(.O (g10319), .I (I13740));
INVX1 gate4345(.O (g17088), .I (I18160));
INVX1 gate4346(.O (g32933), .I (g31376));
INVX1 gate4347(.O (g30329), .I (I28588));
INVX1 gate4348(.O (g9492), .I (g2759));
INVX1 gate4349(.O (I21181), .I (g17413));
INVX1 gate4350(.O (g16136), .I (I17491));
INVX1 gate4351(.O (g7340), .I (g4443));
INVX1 gate4352(.O (g20681), .I (g15483));
INVX1 gate4353(.O (g9600), .I (g3632));
INVX1 gate4354(.O (I23671), .I (g23202));
INVX1 gate4355(.O (g32508), .I (g30825));
INVX1 gate4356(.O (g9574), .I (g6462));
INVX1 gate4357(.O (g31638), .I (g29689));
INVX1 gate4358(.O (g9864), .I (I13424));
INVX1 gate4359(.O (g32634), .I (g30673));
INVX1 gate4360(.O (g32851), .I (g31327));
INVX1 gate4361(.O (g32872), .I (g31327));
INVX1 gate4362(.O (g33638), .I (I31469));
INVX1 gate4363(.O (g35001), .I (I33297));
INVX1 gate4364(.O (g30328), .I (I28585));
INVX1 gate4365(.O (g7907), .I (g3072));
INVX1 gate4366(.O (g11640), .I (I14550));
INVX1 gate4367(.O (g11769), .I (g8626));
INVX1 gate4368(.O (g34539), .I (g34354));
INVX1 gate4369(.O (g9714), .I (g4012));
INVX1 gate4370(.O (g12843), .I (g10359));
INVX1 gate4371(.O (g17497), .I (g14879));
INVX1 gate4372(.O (g22987), .I (g20391));
INVX1 gate4373(.O (g34328), .I (g34096));
INVX1 gate4374(.O (g10059), .I (g6451));
INVX1 gate4375(.O (g23927), .I (g19074));
INVX1 gate4376(.O (I18842), .I (g13809));
INVX1 gate4377(.O (g24429), .I (g22722));
INVX1 gate4378(.O (g19524), .I (g15695));
INVX1 gate4379(.O (I29891), .I (g31578));
INVX1 gate4380(.O (g7517), .I (g962));
INVX1 gate4381(.O (g22658), .I (I21969));
INVX1 gate4382(.O (g29953), .I (g28907));
INVX1 gate4383(.O (g10540), .I (g9392));
INVX1 gate4384(.O (g10058), .I (g6497));
INVX1 gate4385(.O (g31841), .I (g29385));
INVX1 gate4386(.O (g24428), .I (g22722));
INVX1 gate4387(.O (I32096), .I (g33641));
INVX1 gate4388(.O (g33391), .I (g32384));
INVX1 gate4389(.O (g19477), .I (g16431));
INVX1 gate4390(.O (g12869), .I (g10376));
INVX1 gate4391(.O (g16164), .I (I17507));
INVX1 gate4392(.O (g23649), .I (g18833));
INVX1 gate4393(.O (g26683), .I (g25514));
INVX1 gate4394(.O (g7876), .I (g1495));
INVX1 gate4395(.O (g25692), .I (I24839));
INVX1 gate4396(.O (g15614), .I (g14914));
INVX1 gate4397(.O (g22339), .I (g19801));
INVX1 gate4398(.O (g20765), .I (g17748));
INVX1 gate4399(.O (g8938), .I (g4899));
INVX1 gate4400(.O (I19235), .I (g15078));
INVX1 gate4401(.O (I20495), .I (g16283));
INVX1 gate4402(.O (g29800), .I (g28363));
INVX1 gate4403(.O (g10203), .I (g2393));
INVX1 gate4404(.O (g12868), .I (g10377));
INVX1 gate4405(.O (g21903), .I (I21480));
INVX1 gate4406(.O (g14203), .I (g12381));
INVX1 gate4407(.O (g20549), .I (g15277));
INVX1 gate4408(.O (g23648), .I (g18833));
INVX1 gate4409(.O (g13881), .I (I16181));
INVX1 gate4410(.O (I16090), .I (g10430));
INVX1 gate4411(.O (g22338), .I (g19801));
INVX1 gate4412(.O (g23491), .I (g21514));
INVX1 gate4413(.O (I20816), .I (g17088));
INVX1 gate4414(.O (g23903), .I (g18997));
INVX1 gate4415(.O (I33252), .I (g34974));
INVX1 gate4416(.O (I32681), .I (g34429));
INVX1 gate4417(.O (g10044), .I (g5357));
INVX1 gate4418(.O (g34241), .I (I32222));
INVX1 gate4419(.O (g27709), .I (I26337));
INVX1 gate4420(.O (g21604), .I (g15938));
INVX1 gate4421(.O (I22580), .I (g20982));
INVX1 gate4422(.O (I16651), .I (g10542));
INVX1 gate4423(.O (g20548), .I (g15426));
INVX1 gate4424(.O (g8519), .I (g287));
INVX1 gate4425(.O (g8740), .I (I12735));
INVX1 gate4426(.O (g31578), .I (I29199));
INVX1 gate4427(.O (g25013), .I (g23599));
INVX1 gate4428(.O (g31835), .I (g29385));
INVX1 gate4429(.O (g32574), .I (g31070));
INVX1 gate4430(.O (I20985), .I (g16300));
INVX1 gate4431(.O (g24548), .I (g22942));
INVX1 gate4432(.O (I31564), .I (g33204));
INVX1 gate4433(.O (g17296), .I (I18280));
INVX1 gate4434(.O (g25214), .I (g22228));
INVX1 gate4435(.O (g27708), .I (I26334));
INVX1 gate4436(.O (I12418), .I (g55));
INVX1 gate4437(.O (g17644), .I (g15002));
INVX1 gate4438(.O (g20504), .I (g18008));
INVX1 gate4439(.O (g30100), .I (g29131));
INVX1 gate4440(.O (g23563), .I (g20682));
INVX1 gate4441(.O (g10377), .I (g6940));
INVX1 gate4442(.O (g32912), .I (g30735));
INVX1 gate4443(.O (g8606), .I (g4653));
INVX1 gate4444(.O (I18865), .I (g14314));
INVX1 gate4445(.O (I20954), .I (g16228));
INVX1 gate4446(.O (g19748), .I (g17015));
INVX1 gate4447(.O (g10120), .I (g1902));
INVX1 gate4448(.O (g22197), .I (g19074));
INVX1 gate4449(.O (g14377), .I (g12201));
INVX1 gate4450(.O (I11753), .I (g4492));
INVX1 gate4451(.O (g22855), .I (g20391));
INVX1 gate4452(.O (g19276), .I (g17367));
INVX1 gate4453(.O (g9889), .I (g6128));
INVX1 gate4454(.O (g13027), .I (I15647));
INVX1 gate4455(.O (g7110), .I (g6682));
INVX1 gate4456(.O (I14660), .I (g9746));
INVX1 gate4457(.O (g33442), .I (g31937));
INVX1 gate4458(.O (g22870), .I (g20887));
INVX1 gate4459(.O (g22527), .I (g19546));
INVX1 gate4460(.O (I21860), .I (g19638));
INVX1 gate4461(.O (g34683), .I (I32827));
INVX1 gate4462(.O (g28127), .I (g27102));
INVX1 gate4463(.O (g25538), .I (g22594));
INVX1 gate4464(.O (g29216), .I (I27564));
INVX1 gate4465(.O (I32690), .I (g34432));
INVX1 gate4466(.O (g11249), .I (g8405));
INVX1 gate4467(.O (I28838), .I (g29372));
INVX1 gate4468(.O (I13031), .I (g6747));
INVX1 gate4469(.O (g14738), .I (I16821));
INVX1 gate4470(.O (g13249), .I (g10590));
INVX1 gate4471(.O (g14562), .I (g12036));
INVX1 gate4472(.O (g14645), .I (I16755));
INVX1 gate4473(.O (I30861), .I (g32383));
INVX1 gate4474(.O (g20129), .I (g17328));
INVX1 gate4475(.O (g16606), .I (g14110));
INVX1 gate4476(.O (g17197), .I (I18233));
INVX1 gate4477(.O (g18880), .I (g15656));
INVX1 gate4478(.O (g23767), .I (g18997));
INVX1 gate4479(.O (g23794), .I (g19147));
INVX1 gate4480(.O (g21395), .I (g17873));
INVX1 gate4481(.O (g24129), .I (g20857));
INVX1 gate4482(.O (g32592), .I (g30673));
INVX1 gate4483(.O (g20057), .I (g16349));
INVX1 gate4484(.O (g32756), .I (g31021));
INVX1 gate4485(.O (g23395), .I (I22502));
INVX1 gate4486(.O (g24057), .I (g20841));
INVX1 gate4487(.O (g20128), .I (g17533));
INVX1 gate4488(.O (I12167), .I (g5176));
INVX1 gate4489(.O (g14290), .I (I16460));
INVX1 gate4490(.O (g17870), .I (I18842));
INVX1 gate4491(.O (g17411), .I (g14454));
INVX1 gate4492(.O (g17527), .I (g14741));
INVX1 gate4493(.O (g23899), .I (g19277));
INVX1 gate4494(.O (g7002), .I (g5160));
INVX1 gate4495(.O (g13003), .I (I15609));
INVX1 gate4496(.O (g24128), .I (g20720));
INVX1 gate4497(.O (g11204), .I (I14271));
INVX1 gate4498(.O (I14550), .I (g10072));
INVX1 gate4499(.O (g7824), .I (g4169));
INVX1 gate4500(.O (g30991), .I (I28925));
INVX1 gate4501(.O (g6996), .I (g4955));
INVX1 gate4502(.O (g25241), .I (g23651));
INVX1 gate4503(.O (g11779), .I (g9602));
INVX1 gate4504(.O (I18270), .I (g13191));
INVX1 gate4505(.O (g16750), .I (g14454));
INVX1 gate4506(.O (g22867), .I (g20391));
INVX1 gate4507(.O (g34991), .I (I33273));
INVX1 gate4508(.O (g7236), .I (g4608));
INVX1 gate4509(.O (g9285), .I (g2715));
INVX1 gate4510(.O (g20626), .I (g15483));
INVX1 gate4511(.O (g27774), .I (I26381));
INVX1 gate4512(.O (I27401), .I (g27051));
INVX1 gate4513(.O (I11843), .I (g111));
INVX1 gate4514(.O (g23898), .I (g19277));
INVX1 gate4515(.O (g9500), .I (g5495));
INVX1 gate4516(.O (g20323), .I (g17873));
INVX1 gate4517(.O (I21250), .I (g16540));
INVX1 gate4518(.O (g29117), .I (g27886));
INVX1 gate4519(.O (g24626), .I (g23139));
INVX1 gate4520(.O (g33430), .I (g32421));
INVX1 gate4521(.O (g23191), .I (I22289));
INVX1 gate4522(.O (g20533), .I (g17271));
INVX1 gate4523(.O (g10427), .I (g10053));
INVX1 gate4524(.O (g12955), .I (I15577));
INVX1 gate4525(.O (g32820), .I (g31672));
INVX1 gate4526(.O (I18460), .I (g5276));
INVX1 gate4527(.O (g8341), .I (g3119));
INVX1 gate4528(.O (g10366), .I (g6895));
INVX1 gate4529(.O (g24533), .I (g22876));
INVX1 gate4530(.O (g25100), .I (g22384));
INVX1 gate4531(.O (g12879), .I (g10381));
INVX1 gate4532(.O (g22714), .I (g20436));
INVX1 gate4533(.O (g11786), .I (g7549));
INVX1 gate4534(.O (g14366), .I (I16526));
INVX1 gate4535(.O (g17503), .I (g14892));
INVX1 gate4536(.O (I14054), .I (g10028));
INVX1 gate4537(.O (g9184), .I (g6120));
INVX1 gate4538(.O (g23521), .I (g21468));
INVX1 gate4539(.O (g28181), .I (I26700));
INVX1 gate4540(.O (g25771), .I (I24920));
INVX1 gate4541(.O (g20775), .I (g18008));
INVX1 gate4542(.O (g18831), .I (g15224));
INVX1 gate4543(.O (I15647), .I (g12109));
INVX1 gate4544(.O (I23339), .I (g23232));
INVX1 gate4545(.O (g32846), .I (g31376));
INVX1 gate4546(.O (g9339), .I (g2295));
INVX1 gate4547(.O (I19759), .I (g17767));
INVX1 gate4548(.O (g19733), .I (g16856));
INVX1 gate4549(.O (I24558), .I (g23777));
INVX1 gate4550(.O (g12878), .I (g10386));
INVX1 gate4551(.O (g26758), .I (g25389));
INVX1 gate4552(.O (I27749), .I (g28917));
INVX1 gate4553(.O (I20830), .I (g17657));
INVX1 gate4554(.O (g12337), .I (g9340));
INVX1 gate4555(.O (g32731), .I (g31376));
INVX1 gate4556(.O (g31806), .I (g29385));
INVX1 gate4557(.O (g22202), .I (I21784));
INVX1 gate4558(.O (g33806), .I (I31650));
INVX1 gate4559(.O (g9024), .I (g4358));
INVX1 gate4560(.O (I12749), .I (g4575));
INVX1 gate4561(.O (g11826), .I (I14650));
INVX1 gate4562(.O (g17714), .I (g14930));
INVX1 gate4563(.O (g12886), .I (g10393));
INVX1 gate4564(.O (g22979), .I (g20453));
INVX1 gate4565(.O (g20737), .I (g15656));
INVX1 gate4566(.O (g22496), .I (g19510));
INVX1 gate4567(.O (g10403), .I (g7040));
INVX1 gate4568(.O (I21969), .I (g21370));
INVX1 gate4569(.O (g23440), .I (I22557));
INVX1 gate4570(.O (g13999), .I (g11048));
INVX1 gate4571(.O (g7222), .I (g4427));
INVX1 gate4572(.O (g27967), .I (I26479));
INVX1 gate4573(.O (g27994), .I (g26793));
INVX1 gate4574(.O (g33142), .I (g32072));
INVX1 gate4575(.O (g19630), .I (g16897));
INVX1 gate4576(.O (g9809), .I (g6082));
INVX1 gate4577(.O (g20232), .I (g16931));
INVX1 gate4578(.O (I14773), .I (g9581));
INVX1 gate4579(.O (g29814), .I (I28062));
INVX1 gate4580(.O (g17819), .I (I18825));
INVX1 gate4581(.O (g17707), .I (g14758));
INVX1 gate4582(.O (I33047), .I (g34776));
INVX1 gate4583(.O (g30206), .I (g28436));
INVX1 gate4584(.O (g7928), .I (g4776));
INVX1 gate4585(.O (g26744), .I (g25400));
INVX1 gate4586(.O (g12967), .I (g11790));
INVX1 gate4587(.O (g23861), .I (g19147));
INVX1 gate4588(.O (g23573), .I (g20248));
INVX1 gate4589(.O (g32691), .I (g30673));
INVX1 gate4590(.O (g18989), .I (g16000));
INVX1 gate4591(.O (g8879), .I (I12858));
INVX1 gate4592(.O (g8607), .I (g37));
INVX1 gate4593(.O (g11233), .I (g9664));
INVX1 gate4594(.O (I18875), .I (g13782));
INVX1 gate4595(.O (g21247), .I (g15171));
INVX1 gate4596(.O (g23247), .I (g20924));
INVX1 gate4597(.O (g11182), .I (I14241));
INVX1 gate4598(.O (I11708), .I (g3703));
INVX1 gate4599(.O (g7064), .I (g5990));
INVX1 gate4600(.O (g17818), .I (I18822));
INVX1 gate4601(.O (g9672), .I (g5390));
INVX1 gate4602(.O (I13708), .I (g136));
INVX1 gate4603(.O (g20697), .I (g17433));
INVX1 gate4604(.O (g14226), .I (g11618));
INVX1 gate4605(.O (g9077), .I (g504));
INVX1 gate4606(.O (g17496), .I (g14683));
INVX1 gate4607(.O (I19345), .I (g15083));
INVX1 gate4608(.O (g22986), .I (g20330));
INVX1 gate4609(.O (g8659), .I (g2815));
INVX1 gate4610(.O (g25882), .I (g25026));
INVX1 gate4611(.O (g23926), .I (g19074));
INVX1 gate4612(.O (g8358), .I (I12541));
INVX1 gate4613(.O (g18988), .I (g15979));
INVX1 gate4614(.O (I32775), .I (g34512));
INVX1 gate4615(.O (g9477), .I (I13149));
INVX1 gate4616(.O (g8506), .I (g3782));
INVX1 gate4617(.O (I30766), .I (g32363));
INVX1 gate4618(.O (g9523), .I (g6419));
INVX1 gate4619(.O (g24995), .I (g22763));
INVX1 gate4620(.O (g34759), .I (I32935));
INVX1 gate4621(.O (g7785), .I (g4621));
INVX1 gate4622(.O (g16522), .I (g13889));
INVX1 gate4623(.O (g23612), .I (I22745));
INVX1 gate4624(.O (g10572), .I (g10233));
INVX1 gate4625(.O (I25534), .I (g25448));
INVX1 gate4626(.O (I17964), .I (g3661));
INVX1 gate4627(.O (g23388), .I (g21070));
INVX1 gate4628(.O (I15932), .I (g12381));
INVX1 gate4629(.O (g17590), .I (I18523));
INVX1 gate4630(.O (g19476), .I (g16326));
INVX1 gate4631(.O (g12919), .I (I15536));
INVX1 gate4632(.O (I12808), .I (g4322));
INVX1 gate4633(.O (g6799), .I (g199));
INVX1 gate4634(.O (g26804), .I (g25400));
INVX1 gate4635(.O (g20512), .I (g18062));
INVX1 gate4636(.O (g34435), .I (I32476));
INVX1 gate4637(.O (g23777), .I (I22918));
INVX1 gate4638(.O (g23534), .I (I22665));
INVX1 gate4639(.O (I26451), .I (g26862));
INVX1 gate4640(.O (g13932), .I (g11534));
INVX1 gate4641(.O (g32929), .I (g31710));
INVX1 gate4642(.O (g8587), .I (g3689));
INVX1 gate4643(.O (I14839), .I (g9689));
INVX1 gate4644(.O (g23272), .I (g20924));
INVX1 gate4645(.O (g11513), .I (g7948));
INVX1 gate4646(.O (g19454), .I (g16349));
INVX1 gate4647(.O (g7563), .I (g6322));
INVX1 gate4648(.O (g17741), .I (g12972));
INVX1 gate4649(.O (g12918), .I (I15533));
INVX1 gate4650(.O (I18160), .I (g14441));
INVX1 gate4651(.O (I15448), .I (g10877));
INVX1 gate4652(.O (g17384), .I (I18323));
INVX1 gate4653(.O (g32583), .I (g30614));
INVX1 gate4654(.O (g32928), .I (g31672));
INVX1 gate4655(.O (g19570), .I (g16349));
INVX1 gate4656(.O (g19712), .I (g17096));
INVX1 gate4657(.O (g6997), .I (g4578));
INVX1 gate4658(.O (g22150), .I (g21280));
INVX1 gate4659(.O (g11897), .I (I14705));
INVX1 gate4660(.O (I22000), .I (g20277));
INVX1 gate4661(.O (g10490), .I (g9274));
INVX1 gate4662(.O (g9551), .I (g3281));
INVX1 gate4663(.O (g9742), .I (g6144));
INVX1 gate4664(.O (g9104), .I (I12987));
INVX1 gate4665(.O (g23462), .I (I22589));
INVX1 gate4666(.O (g9099), .I (g3706));
INVX1 gate4667(.O (g34345), .I (I32352));
INVX1 gate4668(.O (g9499), .I (g5152));
INVX1 gate4669(.O (g11404), .I (g7596));
INVX1 gate4670(.O (g15750), .I (g13291));
INVX1 gate4671(.O (g34940), .I (g34924));
INVX1 gate4672(.O (g13505), .I (g10981));
INVX1 gate4673(.O (I15717), .I (g6346));
INVX1 gate4674(.O (g16326), .I (I17658));
INVX1 gate4675(.O (g18887), .I (g15373));
INVX1 gate4676(.O (g20445), .I (g15224));
INVX1 gate4677(.O (I31820), .I (g33323));
INVX1 gate4678(.O (I12064), .I (g617));
INVX1 gate4679(.O (g23032), .I (I22211));
INVX1 gate4680(.O (g10376), .I (g6923));
INVX1 gate4681(.O (g10385), .I (I13805));
INVX1 gate4682(.O (g25206), .I (g23613));
INVX1 gate4683(.O (g12598), .I (g7004));
INVX1 gate4684(.O (g14376), .I (g12126));
INVX1 gate4685(.O (g14385), .I (I16541));
INVX1 gate4686(.O (g34848), .I (I33070));
INVX1 gate4687(.O (g19074), .I (I19772));
INVX1 gate4688(.O (g17735), .I (g14807));
INVX1 gate4689(.O (g14297), .I (g10869));
INVX1 gate4690(.O (g20499), .I (g15483));
INVX1 gate4691(.O (g7394), .I (g5637));
INVX1 gate4692(.O (g10980), .I (g9051));
INVX1 gate4693(.O (g11026), .I (g8434));
INVX1 gate4694(.O (I26785), .I (g27013));
INVX1 gate4695(.O (g12086), .I (g9654));
INVX1 gate4696(.O (g32787), .I (g30937));
INVX1 gate4697(.O (g13026), .I (g11018));
INVX1 gate4698(.O (g31863), .I (I29447));
INVX1 gate4699(.O (I14619), .I (g4185));
INVX1 gate4700(.O (g10354), .I (g6811));
INVX1 gate4701(.O (I23315), .I (g21685));
INVX1 gate4702(.O (I33152), .I (g34900));
INVX1 gate4703(.O (g19567), .I (g16164));
INVX1 gate4704(.O (g14095), .I (g11326));
INVX1 gate4705(.O (g29014), .I (g27742));
INVX1 gate4706(.O (g22526), .I (g19801));
INVX1 gate4707(.O (I17569), .I (g14564));
INVX1 gate4708(.O (g9754), .I (g2020));
INVX1 gate4709(.O (g21061), .I (I20929));
INVX1 gate4710(.O (g28126), .I (g27122));
INVX1 gate4711(.O (g18528), .I (I19348));
INVX1 gate4712(.O (g20498), .I (g15348));
INVX1 gate4713(.O (g6802), .I (g468));
INVX1 gate4714(.O (g8284), .I (g5002));
INVX1 gate4715(.O (g23061), .I (g20283));
INVX1 gate4716(.O (g8239), .I (g1056));
INVX1 gate4717(.O (g28250), .I (g27074));
INVX1 gate4718(.O (g10181), .I (g2551));
INVX1 gate4719(.O (g25114), .I (I24278));
INVX1 gate4720(.O (g7557), .I (g1500));
INVX1 gate4721(.O (g8180), .I (g262));
INVX1 gate4722(.O (I17747), .I (g13298));
INVX1 gate4723(.O (g12322), .I (I15162));
INVX1 gate4724(.O (g27977), .I (g26105));
INVX1 gate4725(.O (g32743), .I (g30937));
INVX1 gate4726(.O (g32827), .I (g31672));
INVX1 gate4727(.O (g25082), .I (g22342));
INVX1 gate4728(.O (g8591), .I (g3763));
INVX1 gate4729(.O (g30332), .I (I28597));
INVX1 gate4730(.O (g24056), .I (g20014));
INVX1 gate4731(.O (g9613), .I (g5062));
INVX1 gate4732(.O (g12901), .I (g10404));
INVX1 gate4733(.O (g20611), .I (g18008));
INVX1 gate4734(.O (g17526), .I (I18469));
INVX1 gate4735(.O (g12977), .I (I15590));
INVX1 gate4736(.O (g20080), .I (g17328));
INVX1 gate4737(.O (g7471), .I (g6012));
INVX1 gate4738(.O (g9044), .I (g604));
INVX1 gate4739(.O (g20924), .I (I20895));
INVX1 gate4740(.O (g19519), .I (g16795));
INVX1 gate4741(.O (g24080), .I (g21143));
INVX1 gate4742(.O (g19675), .I (g16987));
INVX1 gate4743(.O (g9444), .I (g5535));
INVX1 gate4744(.O (g9269), .I (g5517));
INVX1 gate4745(.O (g22866), .I (g20330));
INVX1 gate4746(.O (I17814), .I (g3274));
INVX1 gate4747(.O (g32640), .I (g31154));
INVX1 gate4748(.O (g20432), .I (g17847));
INVX1 gate4749(.O (g32769), .I (g31672));
INVX1 gate4750(.O (g23360), .I (I22461));
INVX1 gate4751(.O (g29116), .I (g27837));
INVX1 gate4752(.O (g19518), .I (g16239));
INVX1 gate4753(.O (g8507), .I (g3712));
INVX1 gate4754(.O (g9983), .I (g4239));
INVX1 gate4755(.O (g12656), .I (g7028));
INVX1 gate4756(.O (I15620), .I (g12038));
INVX1 gate4757(.O (I17772), .I (g14888));
INVX1 gate4758(.O (g25849), .I (g24491));
INVX1 gate4759(.O (g9862), .I (g5413));
INVX1 gate4760(.O (I27555), .I (g28142));
INVX1 gate4761(.O (g23447), .I (g21562));
INVX1 gate4762(.O (g32768), .I (g30825));
INVX1 gate4763(.O (g32803), .I (g31376));
INVX1 gate4764(.O (g25399), .I (g22763));
INVX1 gate4765(.O (g12295), .I (g7139));
INVX1 gate4766(.O (I23384), .I (g23362));
INVX1 gate4767(.O (g10190), .I (g6044));
INVX1 gate4768(.O (g29041), .I (I27385));
INVX1 gate4769(.O (g13620), .I (g10556));
INVX1 gate4770(.O (g12823), .I (g9206));
INVX1 gate4771(.O (I17639), .I (g13350));
INVX1 gate4772(.O (I27570), .I (g28262));
INVX1 gate4773(.O (I15811), .I (g11128));
INVX1 gate4774(.O (I21067), .I (g15573));
INVX1 gate4775(.O (I18822), .I (g13745));
INVX1 gate4776(.O (g16509), .I (g13873));
INVX1 gate4777(.O (I32056), .I (g33641));
INVX1 gate4778(.O (g11811), .I (g9724));
INVX1 gate4779(.O (I12712), .I (g59));
INVX1 gate4780(.O (g20145), .I (g17533));
INVX1 gate4781(.O (g34833), .I (I33047));
INVX1 gate4782(.O (g34049), .I (g33678));
INVX1 gate4783(.O (I13010), .I (g6749));
INVX1 gate4784(.O (g31821), .I (g29385));
INVX1 gate4785(.O (g32881), .I (g30673));
INVX1 gate4786(.O (I32988), .I (g34755));
INVX1 gate4787(.O (g24031), .I (g21193));
INVX1 gate4788(.O (I33020), .I (g34781));
INVX1 gate4789(.O (g16508), .I (I17704));
INVX1 gate4790(.O (I24455), .I (g22541));
INVX1 gate4791(.O (g26605), .I (g25293));
INVX1 gate4792(.O (g20650), .I (g15348));
INVX1 gate4793(.O (g23629), .I (g21514));
INVX1 gate4794(.O (g21451), .I (I21162));
INVX1 gate4795(.O (g16872), .I (I18060));
INVX1 gate4796(.O (I12907), .I (g4322));
INVX1 gate4797(.O (g22923), .I (I22124));
INVX1 gate4798(.O (I17416), .I (g13806));
INVX1 gate4799(.O (g23472), .I (g21062));
INVX1 gate4800(.O (g15483), .I (I17128));
INVX1 gate4801(.O (g9534), .I (g90));
INVX1 gate4802(.O (g9729), .I (g5138));
INVX1 gate4803(.O (g9961), .I (g6404));
INVX1 gate4804(.O (g7438), .I (g5983));
INVX1 gate4805(.O (g25263), .I (g22763));
INVX1 gate4806(.O (g29983), .I (g28977));
INVX1 gate4807(.O (g20529), .I (g15509));
INVX1 gate4808(.O (g22300), .I (I21815));
INVX1 gate4809(.O (g26812), .I (g25439));
INVX1 gate4810(.O (I21019), .I (g17325));
INVX1 gate4811(.O (g27017), .I (g25895));
INVX1 gate4812(.O (I27567), .I (g28181));
INVX1 gate4813(.O (g15862), .I (I17355));
INVX1 gate4814(.O (g8515), .I (I12631));
INVX1 gate4815(.O (g34221), .I (I32192));
INVX1 gate4816(.O (g8630), .I (g4843));
INVX1 gate4817(.O (g21246), .I (I20985));
INVX1 gate4818(.O (I27238), .I (g27320));
INVX1 gate4819(.O (g23246), .I (g20785));
INVX1 gate4820(.O (g20528), .I (g15224));
INVX1 gate4821(.O (g20696), .I (g17533));
INVX1 gate4822(.O (g25135), .I (g22457));
INVX1 gate4823(.O (g20330), .I (I20542));
INVX1 gate4824(.O (g9927), .I (g5689));
INVX1 gate4825(.O (g32662), .I (g30614));
INVX1 gate4826(.O (g8300), .I (g1242));
INVX1 gate4827(.O (g32027), .I (I29585));
INVX1 gate4828(.O (I32461), .I (g34244));
INVX1 gate4829(.O (g19577), .I (g16129));
INVX1 gate4830(.O (g17688), .I (I18667));
INVX1 gate4831(.O (g9014), .I (g3004));
INVX1 gate4832(.O (g20764), .I (I20819));
INVX1 gate4833(.O (g10497), .I (g10102));
INVX1 gate4834(.O (I25591), .I (g25380));
INVX1 gate4835(.O (g32890), .I (g30735));
INVX1 gate4836(.O (I33282), .I (g34987));
INVX1 gate4837(.O (I27941), .I (g28803));
INVX1 gate4838(.O (g9414), .I (g2004));
INVX1 gate4839(.O (g7212), .I (g6411));
INVX1 gate4840(.O (g19439), .I (g15885));
INVX1 gate4841(.O (g9660), .I (g3267));
INVX1 gate4842(.O (g9946), .I (g6093));
INVX1 gate4843(.O (g20132), .I (g16931));
INVX1 gate4844(.O (g24365), .I (g22594));
INVX1 gate4845(.O (g20869), .I (g15615));
INVX1 gate4846(.O (g13412), .I (g11963));
INVX1 gate4847(.O (g23776), .I (g21177));
INVX1 gate4848(.O (g34947), .I (g34938));
INVX1 gate4849(.O (I12382), .I (g47));
INVX1 gate4850(.O (g24132), .I (g19890));
INVX1 gate4851(.O (g32482), .I (g30614));
INVX1 gate4852(.O (g24869), .I (I24041));
INVX1 gate4853(.O (g24960), .I (g23716));
INVX1 gate4854(.O (g19438), .I (g16249));
INVX1 gate4855(.O (I12519), .I (g3447));
INVX1 gate4856(.O (g17157), .I (g13350));
INVX1 gate4857(.O (I12176), .I (g5523));
INVX1 gate4858(.O (g9903), .I (g681));
INVX1 gate4859(.O (g13133), .I (g11330));
INVX1 gate4860(.O (g32710), .I (g30825));
INVX1 gate4861(.O (I12092), .I (g790));
INVX1 gate4862(.O (g14700), .I (g12512));
INVX1 gate4863(.O (g21355), .I (g17821));
INVX1 gate4864(.O (g32552), .I (g30825));
INVX1 gate4865(.O (g31834), .I (g29385));
INVX1 gate4866(.O (g23355), .I (g21070));
INVX1 gate4867(.O (g34812), .I (I33024));
INVX1 gate4868(.O (g10658), .I (I13979));
INVX1 gate4869(.O (g21370), .I (g16323));
INVX1 gate4870(.O (g23859), .I (g19074));
INVX1 gate4871(.O (g28819), .I (I27271));
INVX1 gate4872(.O (g16311), .I (g13273));
INVX1 gate4873(.O (g32779), .I (g30937));
INVX1 gate4874(.O (I17442), .I (g13638));
INVX1 gate4875(.O (g18878), .I (g15426));
INVX1 gate4876(.O (g24161), .I (I23327));
INVX1 gate4877(.O (g29130), .I (g27907));
INVX1 gate4878(.O (I32696), .I (g34434));
INVX1 gate4879(.O (I32843), .I (g34499));
INVX1 gate4880(.O (g7993), .I (I12333));
INVX1 gate4881(.O (g20709), .I (g15426));
INVX1 gate4882(.O (g11011), .I (g10274));
INVX1 gate4883(.O (g22854), .I (g20330));
INVX1 gate4884(.O (g34951), .I (g34941));
INVX1 gate4885(.O (g34972), .I (I33232));
INVX1 gate4886(.O (g23858), .I (g18997));
INVX1 gate4887(.O (g13011), .I (I15623));
INVX1 gate4888(.O (I12935), .I (g6753));
INVX1 gate4889(.O (g32778), .I (g31021));
INVX1 gate4890(.O (g18886), .I (g16000));
INVX1 gate4891(.O (I31803), .I (g33176));
INVX1 gate4892(.O (g9036), .I (g5084));
INVX1 gate4893(.O (I18313), .I (g13350));
INVX1 gate4894(.O (g25221), .I (g23653));
INVX1 gate4895(.O (I22275), .I (g20127));
INVX1 gate4896(.O (g8440), .I (g3431));
INVX1 gate4897(.O (g20708), .I (g15426));
INVX1 gate4898(.O (g22763), .I (I22046));
INVX1 gate4899(.O (g9679), .I (g5475));
INVX1 gate4900(.O (g23172), .I (I22275));
INVX1 gate4901(.O (g13716), .I (I16090));
INVX1 gate4902(.O (I17615), .I (g13251));
INVX1 gate4903(.O (g20087), .I (g17249));
INVX1 gate4904(.O (g32786), .I (g31021));
INVX1 gate4905(.O (g33726), .I (I31581));
INVX1 gate4906(.O (I32960), .I (g34653));
INVX1 gate4907(.O (g8123), .I (g3808));
INVX1 gate4908(.O (g19566), .I (g16136));
INVX1 gate4909(.O (g14338), .I (I16502));
INVX1 gate4910(.O (g24087), .I (g21143));
INVX1 gate4911(.O (I18276), .I (g1075));
INVX1 gate4912(.O (I18285), .I (g13638));
INVX1 gate4913(.O (g28590), .I (g27724));
INVX1 gate4914(.O (g23844), .I (g21308));
INVX1 gate4915(.O (g32647), .I (g31154));
INVX1 gate4916(.O (g23394), .I (I22499));
INVX1 gate4917(.O (I32868), .I (g34579));
INVX1 gate4918(.O (g9831), .I (g2269));
INVX1 gate4919(.O (g32945), .I (g30937));
INVX1 gate4920(.O (g33436), .I (I30962));
INVX1 gate4921(.O (g22660), .I (g19140));
INVX1 gate4922(.O (g15509), .I (I17136));
INVX1 gate4923(.O (I19012), .I (g15060));
INVX1 gate4924(.O (g17763), .I (g15011));
INVX1 gate4925(.O (g8666), .I (g3703));
INVX1 gate4926(.O (g10060), .I (g6541));
INVX1 gate4927(.O (I18900), .I (g16767));
INVX1 gate4928(.O (g27976), .I (g26703));
INVX1 gate4929(.O (g27985), .I (g26131));
INVX1 gate4930(.O (I32161), .I (g33791));
INVX1 gate4931(.O (g32826), .I (g30825));
INVX1 gate4932(.O (g25273), .I (g23978));
INVX1 gate4933(.O (g29863), .I (g28410));
INVX1 gate4934(.O (g24043), .I (g20982));
INVX1 gate4935(.O (g10197), .I (g31));
INVX1 gate4936(.O (I21300), .I (g18598));
INVX1 gate4937(.O (g22456), .I (g19801));
INVX1 gate4938(.O (g12976), .I (I15587));
INVX1 gate4939(.O (g15634), .I (I17188));
INVX1 gate4940(.O (I23688), .I (g23244));
INVX1 gate4941(.O (I23300), .I (g21665));
INVX1 gate4942(.O (g14197), .I (g12160));
INVX1 gate4943(.O (g32090), .I (g31003));
INVX1 gate4944(.O (g9805), .I (g5485));
INVX1 gate4945(.O (g9916), .I (g3625));
INVX1 gate4946(.O (g19653), .I (g16897));
INVX1 gate4947(.O (g33346), .I (g32132));
INVX1 gate4948(.O (I18101), .I (g13416));
INVX1 gate4949(.O (I32225), .I (g34121));
INVX1 gate4950(.O (g10527), .I (I13892));
INVX1 gate4951(.O (I12577), .I (g1227));
INVX1 gate4952(.O (g10411), .I (g7086));
INVX1 gate4953(.O (g23420), .I (g21514));
INVX1 gate4954(.O (g9749), .I (g1691));
INVX1 gate4955(.O (I18177), .I (g13191));
INVX1 gate4956(.O (I18560), .I (g5969));
INVX1 gate4957(.O (g32651), .I (g31376));
INVX1 gate4958(.O (g18918), .I (I19704));
INVX1 gate4959(.O (g32672), .I (g31579));
INVX1 gate4960(.O (I19789), .I (g17793));
INVX1 gate4961(.O (g24069), .I (g19968));
INVX1 gate4962(.O (g22550), .I (I21922));
INVX1 gate4963(.O (I33027), .I (g34767));
INVX1 gate4964(.O (g26788), .I (g25349));
INVX1 gate4965(.O (g26724), .I (g25341));
INVX1 gate4966(.O (g20657), .I (g17433));
INVX1 gate4967(.O (g20774), .I (g18008));
INVX1 gate4968(.O (I26427), .I (g26859));
INVX1 gate4969(.O (g8655), .I (g2787));
INVX1 gate4970(.O (g23446), .I (g21562));
INVX1 gate4971(.O (I16057), .I (g10430));
INVX1 gate4972(.O (I28908), .I (g30182));
INVX1 gate4973(.O (g19636), .I (g16987));
INVX1 gate4974(.O (g23227), .I (g20924));
INVX1 gate4975(.O (g30012), .I (I28241));
INVX1 gate4976(.O (g19415), .I (g15758));
INVX1 gate4977(.O (g24068), .I (g19919));
INVX1 gate4978(.O (g24375), .I (g22722));
INVX1 gate4979(.O (g21059), .I (g15509));
INVX1 gate4980(.O (I33249), .I (g34971));
INVX1 gate4981(.O (g7462), .I (g2599));
INVX1 gate4982(.O (g23059), .I (g20453));
INVX1 gate4983(.O (g31797), .I (g29385));
INVX1 gate4984(.O (g6838), .I (g1724));
INVX1 gate4985(.O (g13096), .I (I15727));
INVX1 gate4986(.O (g33641), .I (I31474));
INVX1 gate4987(.O (g32932), .I (g31327));
INVX1 gate4988(.O (g33797), .I (g33306));
INVX1 gate4989(.O (I31482), .I (g33204));
INVX1 gate4990(.O (g19852), .I (g17015));
INVX1 gate4991(.O (g22721), .I (I22028));
INVX1 gate4992(.O (g10503), .I (g8879));
INVX1 gate4993(.O (I16626), .I (g11986));
INVX1 gate4994(.O (g21058), .I (g15426));
INVX1 gate4995(.O (g6809), .I (g341));
INVX1 gate4996(.O (g32513), .I (g31376));
INVX1 gate4997(.O (I20864), .I (g16960));
INVX1 gate4998(.O (g23058), .I (g20453));
INVX1 gate4999(.O (g32449), .I (I29977));
INVX1 gate5000(.O (g14503), .I (g12256));
INVX1 gate5001(.O (g16691), .I (g14160));
INVX1 gate5002(.O (I24022), .I (g22182));
INVX1 gate5003(.O (g19963), .I (g16326));
INVX1 gate5004(.O (g12842), .I (g10355));
INVX1 gate5005(.O (g34473), .I (g34426));
INVX1 gate5006(.O (I12083), .I (g568));
INVX1 gate5007(.O (g17085), .I (g14238));
INVX1 gate5008(.O (I31779), .I (g33212));
INVX1 gate5009(.O (g24171), .I (I23357));
INVX1 gate5010(.O (g32897), .I (g30735));
INVX1 gate5011(.O (g32961), .I (g31376));
INVX1 gate5012(.O (g23203), .I (g20073));
INVX1 gate5013(.O (g8839), .I (I12819));
INVX1 gate5014(.O (g34789), .I (I32997));
INVX1 gate5015(.O (g7788), .I (g4674));
INVX1 gate5016(.O (g11429), .I (g7616));
INVX1 gate5017(.O (g17721), .I (g12915));
INVX1 gate5018(.O (g29372), .I (I27738));
INVX1 gate5019(.O (g10581), .I (g9529));
INVX1 gate5020(.O (I16775), .I (g12183));
INVX1 gate5021(.O (g13857), .I (I16163));
INVX1 gate5022(.O (g32505), .I (g31566));
INVX1 gate5023(.O (g20994), .I (g15615));
INVX1 gate5024(.O (g9095), .I (g3368));
INVX1 gate5025(.O (g32404), .I (I29936));
INVX1 gate5026(.O (I14800), .I (g10107));
INVX1 gate5027(.O (g33136), .I (g32057));
INVX1 gate5028(.O (g9037), .I (g164));
INVX1 gate5029(.O (g14714), .I (g11405));
INVX1 gate5030(.O (g33635), .I (g33436));
INVX1 gate5031(.O (g24994), .I (g22432));
INVX1 gate5032(.O (g14315), .I (I16479));
INVX1 gate5033(.O (g30325), .I (I28576));
INVX1 gate5034(.O (g34788), .I (I32994));
INVX1 gate5035(.O (g11793), .I (I14633));
INVX1 gate5036(.O (g11428), .I (g7615));
INVX1 gate5037(.O (g26682), .I (g25309));
INVX1 gate5038(.O (g9653), .I (g2441));
INVX1 gate5039(.O (g17431), .I (I18376));
INVX1 gate5040(.O (g13793), .I (I16120));
INVX1 gate5041(.O (g22341), .I (g19801));
INVX1 gate5042(.O (g32717), .I (g30735));
INVX1 gate5043(.O (g34325), .I (g34092));
INVX1 gate5044(.O (I15765), .I (g10823));
INVX1 gate5045(.O (I18009), .I (g13680));
INVX1 gate5046(.O (g21281), .I (g16286));
INVX1 gate5047(.O (g18977), .I (g16100));
INVX1 gate5048(.O (I31786), .I (g33197));
INVX1 gate5049(.O (I32970), .I (g34716));
INVX1 gate5050(.O (g22156), .I (g19147));
INVX1 gate5051(.O (g27830), .I (g26802));
INVX1 gate5052(.O (g21902), .I (I21477));
INVX1 gate5053(.O (g34920), .I (I33152));
INVX1 gate5054(.O (g8172), .I (g3873));
INVX1 gate5055(.O (g8278), .I (g3096));
INVX1 gate5056(.O (g34434), .I (I32473));
INVX1 gate5057(.O (g23902), .I (g21468));
INVX1 gate5058(.O (g23301), .I (g21037));
INVX1 gate5059(.O (g34358), .I (I32364));
INVX1 gate5060(.O (g28917), .I (I27314));
INVX1 gate5061(.O (g23377), .I (g21070));
INVX1 gate5062(.O (I32878), .I (g34501));
INVX1 gate5063(.O (g22180), .I (g19210));
INVX1 gate5064(.O (g24425), .I (g22722));
INVX1 gate5065(.O (g19554), .I (g16861));
INVX1 gate5066(.O (g10111), .I (g1858));
INVX1 gate5067(.O (g12830), .I (g9995));
INVX1 gate5068(.O (g12893), .I (g10391));
INVX1 gate5069(.O (I11816), .I (g93));
INVX1 gate5070(.O (g16583), .I (g14069));
INVX1 gate5071(.O (g7392), .I (g4438));
INVX1 gate5072(.O (g20919), .I (g15224));
INVX1 gate5073(.O (g15756), .I (g13315));
INVX1 gate5074(.O (I25146), .I (g24911));
INVX1 gate5075(.O (g34946), .I (g34934));
INVX1 gate5076(.O (I25562), .I (g25250));
INVX1 gate5077(.O (g19609), .I (g16264));
INVX1 gate5078(.O (g8235), .I (I12463));
INVX1 gate5079(.O (g8343), .I (g3447));
INVX1 gate5080(.O (I18476), .I (g14031));
INVX1 gate5081(.O (g34121), .I (I32056));
INVX1 gate5082(.O (I14964), .I (g10230));
INVX1 gate5083(.O (g19200), .I (I19789));
INVX1 gate5084(.O (g21562), .I (I21199));
INVX1 gate5085(.O (g9752), .I (g1840));
INVX1 gate5086(.O (g12865), .I (g10372));
INVX1 gate5087(.O (g20010), .I (g17226));
INVX1 gate5088(.O (g8282), .I (g3841));
INVX1 gate5089(.O (g20918), .I (g15224));
INVX1 gate5090(.O (g23645), .I (g20875));
INVX1 gate5091(.O (g8566), .I (g3831));
INVX1 gate5092(.O (I18555), .I (g5630));
INVX1 gate5093(.O (g24010), .I (g21562));
INVX1 gate5094(.O (g9917), .I (I13473));
INVX1 gate5095(.O (I32967), .I (g34648));
INVX1 gate5096(.O (I32994), .I (g34739));
INVX1 gate5097(.O (g10741), .I (g8411));
INVX1 gate5098(.O (I21480), .I (g18696));
INVX1 gate5099(.O (g7854), .I (g1152));
INVX1 gate5100(.O (g13504), .I (g11303));
INVX1 gate5101(.O (g25541), .I (g22763));
INVX1 gate5102(.O (g20545), .I (g15373));
INVX1 gate5103(.O (g20079), .I (g17328));
INVX1 gate5104(.O (g20444), .I (g15373));
INVX1 gate5105(.O (g21290), .I (I21029));
INVX1 gate5106(.O (g32723), .I (g31327));
INVX1 gate5107(.O (I31672), .I (g33149));
INVX1 gate5108(.O (g10384), .I (I13802));
INVX1 gate5109(.O (g8134), .I (I12415));
INVX1 gate5110(.O (g23290), .I (g20924));
INVX1 gate5111(.O (I33182), .I (g34910));
INVX1 gate5112(.O (I13374), .I (g6490));
INVX1 gate5113(.O (g8334), .I (g3034));
INVX1 gate5114(.O (g24079), .I (g20998));
INVX1 gate5115(.O (g21698), .I (g18562));
INVX1 gate5116(.O (g14384), .I (I16538));
INVX1 gate5117(.O (g22667), .I (g21156));
INVX1 gate5118(.O (g34682), .I (I32824));
INVX1 gate5119(.O (g29209), .I (I27543));
INVX1 gate5120(.O (g20599), .I (g18065));
INVX1 gate5121(.O (g6926), .I (g3853));
INVX1 gate5122(.O (I16512), .I (g12811));
INVX1 gate5123(.O (g23698), .I (g21611));
INVX1 gate5124(.O (I12415), .I (g48));
INVX1 gate5125(.O (g11317), .I (I14346));
INVX1 gate5126(.O (g20078), .I (g16846));
INVX1 gate5127(.O (I12333), .I (g45));
INVX1 gate5128(.O (g32433), .I (I29961));
INVX1 gate5129(.O (g19745), .I (g16877));
INVX1 gate5130(.O (g24078), .I (g20857));
INVX1 gate5131(.O (g6754), .I (I11617));
INVX1 gate5132(.O (g12705), .I (g7051));
INVX1 gate5133(.O (g20598), .I (g17929));
INVX1 gate5134(.O (g32620), .I (g30673));
INVX1 gate5135(.O (I28579), .I (g29474));
INVX1 gate5136(.O (g20086), .I (I20355));
INVX1 gate5137(.O (g19799), .I (g17062));
INVX1 gate5138(.O (g25325), .I (g22228));
INVX1 gate5139(.O (I32458), .I (g34243));
INVX1 gate5140(.O (g11129), .I (g7994));
INVX1 gate5141(.O (I25366), .I (g24477));
INVX1 gate5142(.O (g8804), .I (g4035));
INVX1 gate5143(.O (g10150), .I (g1700));
INVX1 gate5144(.O (g24086), .I (g20998));
INVX1 gate5145(.O (g16743), .I (g13986));
INVX1 gate5146(.O (g21427), .I (g17367));
INVX1 gate5147(.O (g15731), .I (g13326));
INVX1 gate5148(.O (g9364), .I (g5041));
INVX1 gate5149(.O (g10877), .I (I14079));
INVX1 gate5150(.O (g23427), .I (I22542));
INVX1 gate5151(.O (g25535), .I (g22763));
INVX1 gate5152(.O (g32811), .I (g30735));
INVX1 gate5153(.O (I12963), .I (g640));
INVX1 gate5154(.O (g14150), .I (g12381));
INVX1 gate5155(.O (g21366), .I (I21100));
INVX1 gate5156(.O (g32646), .I (g31070));
INVX1 gate5157(.O (g8792), .I (I12790));
INVX1 gate5158(.O (g7219), .I (g4405));
INVX1 gate5159(.O (g19798), .I (g17200));
INVX1 gate5160(.O (I28014), .I (g28158));
INVX1 gate5161(.O (g11128), .I (g7993));
INVX1 gate5162(.O (g7640), .I (I12128));
INVX1 gate5163(.O (I18238), .I (g13144));
INVX1 gate5164(.O (g10019), .I (g6479));
INVX1 gate5165(.O (g28157), .I (I26670));
INVX1 gate5166(.O (I15626), .I (g12041));
INVX1 gate5167(.O (g22210), .I (I21792));
INVX1 gate5168(.O (g20322), .I (g17873));
INVX1 gate5169(.O (g32971), .I (g31672));
INVX1 gate5170(.O (g7431), .I (g2555));
INVX1 gate5171(.O (I32079), .I (g33937));
INVX1 gate5172(.O (g7252), .I (g1592));
INVX1 gate5173(.O (g16640), .I (I17834));
INVX1 gate5174(.O (g29913), .I (g28840));
INVX1 gate5175(.O (g34760), .I (I32938));
INVX1 gate5176(.O (g7812), .I (I12214));
INVX1 gate5177(.O (g16769), .I (g13530));
INVX1 gate5178(.O (g20159), .I (g17533));
INVX1 gate5179(.O (g34134), .I (I32079));
INVX1 gate5180(.O (g25121), .I (g22432));
INVX1 gate5181(.O (g20901), .I (I20867));
INVX1 gate5182(.O (g13626), .I (g11273));
INVX1 gate5183(.O (g20532), .I (g15277));
INVX1 gate5184(.O (g17487), .I (I18414));
INVX1 gate5185(.O (I27576), .I (g28173));
INVX1 gate5186(.O (I15533), .I (g11867));
INVX1 gate5187(.O (g24159), .I (I23321));
INVX1 gate5188(.O (g13323), .I (g11048));
INVX1 gate5189(.O (g24125), .I (g19890));
INVX1 gate5190(.O (g6983), .I (g4698));
INVX1 gate5191(.O (I18382), .I (g13350));
INVX1 gate5192(.O (g21661), .I (I21222));
INVX1 gate5193(.O (g17502), .I (g14697));
INVX1 gate5194(.O (g16768), .I (g13223));
INVX1 gate5195(.O (I19927), .I (g17408));
INVX1 gate5196(.O (g20158), .I (g16971));
INVX1 gate5197(.O (g8113), .I (g3466));
INVX1 gate5198(.O (g12938), .I (I15556));
INVX1 gate5199(.O (I16498), .I (g10430));
INVX1 gate5200(.O (g23403), .I (I22512));
INVX1 gate5201(.O (g23547), .I (g21611));
INVX1 gate5202(.O (g23895), .I (g19147));
INVX1 gate5203(.O (I13424), .I (g5689));
INVX1 gate5204(.O (g24158), .I (I23318));
INVX1 gate5205(.O (g33750), .I (I31607));
INVX1 gate5206(.O (I18092), .I (g3668));
INVX1 gate5207(.O (g7405), .I (g1936));
INVX1 gate5208(.O (g13298), .I (I15862));
INVX1 gate5209(.O (g19732), .I (g17096));
INVX1 gate5210(.O (I22264), .I (g20100));
INVX1 gate5211(.O (I30980), .I (g32132));
INVX1 gate5212(.O (I24008), .I (g22182));
INVX1 gate5213(.O (g29905), .I (g28783));
INVX1 gate5214(.O (g20561), .I (g17873));
INVX1 gate5215(.O (g20656), .I (g17249));
INVX1 gate5216(.O (g9553), .I (I13202));
INVX1 gate5217(.O (I18518), .I (g13835));
INVX1 gate5218(.O (I18154), .I (g13177));
INVX1 gate5219(.O (g23226), .I (g20924));
INVX1 gate5220(.O (g7765), .I (g4165));
INVX1 gate5221(.O (g20680), .I (g15348));
INVX1 gate5222(.O (g26648), .I (g25115));
INVX1 gate5223(.O (g20144), .I (g17533));
INVX1 gate5224(.O (g10402), .I (g7023));
INVX1 gate5225(.O (g23715), .I (g20764));
INVX1 gate5226(.O (g23481), .I (I22604));
INVX1 gate5227(.O (g32850), .I (g30937));
INVX1 gate5228(.O (g31796), .I (g29385));
INVX1 gate5229(.O (g19761), .I (g17015));
INVX1 gate5230(.O (I12608), .I (g1582));
INVX1 gate5231(.O (g12875), .I (I15494));
INVX1 gate5232(.O (I21734), .I (g19268));
INVX1 gate5233(.O (g6961), .I (I11734));
INVX1 gate5234(.O (g8567), .I (g4082));
INVX1 gate5235(.O (I21930), .I (g21297));
INVX1 gate5236(.O (g34927), .I (I33173));
INVX1 gate5237(.O (g7733), .I (g4093));
INVX1 gate5238(.O (I22422), .I (g19330));
INVX1 gate5239(.O (I15697), .I (g6000));
INVX1 gate5240(.O (I17873), .I (g15017));
INVX1 gate5241(.O (g31840), .I (g29385));
INVX1 gate5242(.O (I32158), .I (g33791));
INVX1 gate5243(.O (g12218), .I (I15073));
INVX1 gate5244(.O (g32896), .I (g31376));
INVX1 gate5245(.O (g12837), .I (g10354));
INVX1 gate5246(.O (g23127), .I (g21163));
INVX1 gate5247(.O (g6927), .I (g3845));
INVX1 gate5248(.O (I21838), .I (g19263));
INVX1 gate5249(.O (g25134), .I (g22417));
INVX1 gate5250(.O (g10001), .I (g6105));
INVX1 gate5251(.O (g22975), .I (g20391));
INVX1 gate5252(.O (g13856), .I (I16160));
INVX1 gate5253(.O (I23694), .I (g23252));
INVX1 gate5254(.O (I29248), .I (g29491));
INVX1 gate5255(.O (g9888), .I (g5831));
INVX1 gate5256(.O (g10077), .I (g1724));
INVX1 gate5257(.O (g13995), .I (g11261));
INVX1 gate5258(.O (I33149), .I (g34900));
INVX1 gate5259(.O (g8593), .I (g3759));
INVX1 gate5260(.O (g29153), .I (g27937));
INVX1 gate5261(.O (g24966), .I (g22763));
INVX1 gate5262(.O (g7073), .I (g6191));
INVX1 gate5263(.O (I12799), .I (g59));
INVX1 gate5264(.O (g20631), .I (g15171));
INVX1 gate5265(.O (g17815), .I (g14348));
INVX1 gate5266(.O (g10597), .I (g10233));
INVX1 gate5267(.O (g23490), .I (g21514));
INVX1 gate5268(.O (g25506), .I (g22228));
INVX1 gate5269(.O (g9429), .I (g3723));
INVX1 gate5270(.O (I13705), .I (g63));
INVX1 gate5271(.O (I29204), .I (g29505));
INVX1 gate5272(.O (g32716), .I (g31376));
INVX1 gate5273(.O (g7473), .I (g6697));
INVX1 gate5274(.O (g16249), .I (I17590));
INVX1 gate5275(.O (g18976), .I (g16100));
INVX1 gate5276(.O (g14597), .I (I16713));
INVX1 gate5277(.O (g19539), .I (g16129));
INVX1 gate5278(.O (g6946), .I (I11721));
INVX1 gate5279(.O (g24017), .I (g18833));
INVX1 gate5280(.O (g11512), .I (g7634));
INVX1 gate5281(.O (g34648), .I (I32752));
INVX1 gate5282(.O (g24364), .I (g22722));
INVX1 gate5283(.O (g17677), .I (g14882));
INVX1 gate5284(.O (g34491), .I (I32550));
INVX1 gate5285(.O (I22542), .I (g19773));
INVX1 gate5286(.O (g16482), .I (g13464));
INVX1 gate5287(.O (I17834), .I (g14977));
INVX1 gate5288(.O (g31522), .I (I29185));
INVX1 gate5289(.O (g32582), .I (g31170));
INVX1 gate5290(.O (g7980), .I (g3161));
INVX1 gate5291(.O (g21297), .I (I21042));
INVX1 gate5292(.O (g18954), .I (g17427));
INVX1 gate5293(.O (g23376), .I (g21070));
INVX1 gate5294(.O (g23385), .I (I22488));
INVX1 gate5295(.O (I25095), .I (g25265));
INVX1 gate5296(.O (g19538), .I (g16100));
INVX1 gate5297(.O (g6903), .I (g3502));
INVX1 gate5298(.O (g7069), .I (g6137));
INVX1 gate5299(.O (g9281), .I (I13057));
INVX1 gate5300(.O (I12805), .I (g4098));
INVX1 gate5301(.O (g26990), .I (g26105));
INVX1 gate5302(.O (g34755), .I (I32929));
INVX1 gate5303(.O (g23889), .I (g20682));
INVX1 gate5304(.O (I13124), .I (g2729));
INVX1 gate5305(.O (I18728), .I (g6012));
INVX1 gate5306(.O (I21210), .I (g17526));
INVX1 gate5307(.O (g23354), .I (g20453));
INVX1 gate5308(.O (I14579), .I (g8792));
INVX1 gate5309(.O (g22169), .I (g19147));
INVX1 gate5310(.O (I26700), .I (g27956));
INVX1 gate5311(.O (g34770), .I (I32956));
INVX1 gate5312(.O (g12470), .I (I15284));
INVX1 gate5313(.O (g7540), .I (I12026));
INVX1 gate5314(.O (g8160), .I (g3423));
INVX1 gate5315(.O (g22884), .I (g20453));
INVX1 gate5316(.O (g34981), .I (g34973));
INVX1 gate5317(.O (g23888), .I (g18997));
INVX1 gate5318(.O (g23824), .I (g21271));
INVX1 gate5319(.O (I15831), .I (g10416));
INVX1 gate5320(.O (g32627), .I (g30673));
INVX1 gate5321(.O (g28307), .I (g27306));
INVX1 gate5322(.O (g32959), .I (g30937));
INVX1 gate5323(.O (g32925), .I (g31327));
INVX1 gate5324(.O (g21181), .I (g15426));
INVX1 gate5325(.O (g22168), .I (g19147));
INVX1 gate5326(.O (g10102), .I (g6727));
INVX1 gate5327(.O (g10157), .I (g2036));
INVX1 gate5328(.O (g31862), .I (I29444));
INVX1 gate5329(.O (g32958), .I (g31710));
INVX1 gate5330(.O (I15316), .I (g10087));
INVX1 gate5331(.O (I19719), .I (g17431));
INVX1 gate5332(.O (g8450), .I (g3821));
INVX1 gate5333(.O (g24023), .I (g21127));
INVX1 gate5334(.O (g26718), .I (g25168));
INVX1 gate5335(.O (I32364), .I (g34208));
INVX1 gate5336(.O (g17791), .I (g14950));
INVX1 gate5337(.O (g20571), .I (g15277));
INVX1 gate5338(.O (g9684), .I (g6191));
INVX1 gate5339(.O (g11316), .I (g8967));
INVX1 gate5340(.O (g9745), .I (g6537));
INVX1 gate5341(.O (g12075), .I (I14935));
INVX1 gate5342(.O (I17436), .I (g13416));
INVX1 gate5343(.O (g28431), .I (I26925));
INVX1 gate5344(.O (g9639), .I (g1752));
INVX1 gate5345(.O (I18906), .I (g16963));
INVX1 gate5346(.O (g9338), .I (g1870));
INVX1 gate5347(.O (g24571), .I (g22942));
INVX1 gate5348(.O (g10231), .I (g2661));
INVX1 gate5349(.O (I18083), .I (g13394));
INVX1 gate5350(.O (g9963), .I (g7));
INVX1 gate5351(.O (I26296), .I (g26820));
INVX1 gate5352(.O (g33326), .I (g32318));
INVX1 gate5353(.O (g17410), .I (g12955));
INVX1 gate5354(.O (I12761), .I (g4188));
INVX1 gate5355(.O (g11498), .I (I14475));
INVX1 gate5356(.O (g34767), .I (I32947));
INVX1 gate5357(.O (g14231), .I (g12246));
INVX1 gate5358(.O (g26832), .I (g24850));
INVX1 gate5359(.O (g34845), .I (g34773));
INVX1 gate5360(.O (g32603), .I (g31070));
INVX1 gate5361(.O (g6831), .I (g1413));
INVX1 gate5362(.O (I22464), .I (g21222));
INVX1 gate5363(.O (g23931), .I (g20875));
INVX1 gate5364(.O (g32742), .I (g31021));
INVX1 gate5365(.O (I29233), .I (g30295));
INVX1 gate5366(.O (g9309), .I (g5462));
INVX1 gate5367(.O (I23306), .I (g21673));
INVX1 gate5368(.O (g30990), .I (g29676));
INVX1 gate5369(.O (I18304), .I (g14790));
INVX1 gate5370(.O (g19771), .I (g17096));
INVX1 gate5371(.O (g25240), .I (g23650));
INVX1 gate5372(.O (g32944), .I (g31021));
INVX1 gate5373(.O (I29182), .I (g30012));
INVX1 gate5374(.O (g29474), .I (I27758));
INVX1 gate5375(.O (g34990), .I (I33270));
INVX1 gate5376(.O (g11989), .I (I14839));
INVX1 gate5377(.O (I25190), .I (g25423));
INVX1 gate5378(.O (g16826), .I (I18034));
INVX1 gate5379(.O (g17479), .I (g14855));
INVX1 gate5380(.O (g21426), .I (g15277));
INVX1 gate5381(.O (g8179), .I (g4999));
INVX1 gate5382(.O (g12037), .I (I14893));
INVX1 gate5383(.O (g20495), .I (g17926));
INVX1 gate5384(.O (g23426), .I (I22539));
INVX1 gate5385(.O (g25903), .I (I25005));
INVX1 gate5386(.O (g27984), .I (g26737));
INVX1 gate5387(.O (I13875), .I (g1233));
INVX1 gate5388(.O (g33702), .I (I31545));
INVX1 gate5389(.O (g9808), .I (g5827));
INVX1 gate5390(.O (g19683), .I (g16931));
INVX1 gate5391(.O (g23190), .I (I22286));
INVX1 gate5392(.O (I16709), .I (g10430));
INVX1 gate5393(.O (g11988), .I (I14836));
INVX1 gate5394(.O (I21815), .I (g21308));
INVX1 gate5395(.O (g17478), .I (g14996));
INVX1 gate5396(.O (g28156), .I (I26667));
INVX1 gate5397(.O (I12013), .I (g590));
INVX1 gate5398(.O (g17015), .I (I18143));
INVX1 gate5399(.O (g32681), .I (g30735));
INVX1 gate5400(.O (I32309), .I (g34210));
INVX1 gate5401(.O (I12214), .I (g6561));
INVX1 gate5402(.O (g16182), .I (g13846));
INVX1 gate5403(.O (g16651), .I (g14005));
INVX1 gate5404(.O (I22153), .I (g20014));
INVX1 gate5405(.O (g23520), .I (g21468));
INVX1 gate5406(.O (g27155), .I (g26131));
INVX1 gate5407(.O (g9759), .I (g2265));
INVX1 gate5408(.O (g18830), .I (g18008));
INVX1 gate5409(.O (I16471), .I (g12367));
INVX1 gate5410(.O (g17486), .I (I18411));
INVX1 gate5411(.O (g7898), .I (g4991));
INVX1 gate5412(.O (g25563), .I (g22594));
INVX1 gate5413(.O (g32802), .I (g31327));
INVX1 gate5414(.O (g32857), .I (g30937));
INVX1 gate5415(.O (g22223), .I (g19210));
INVX1 gate5416(.O (g13271), .I (I15834));
INVX1 gate5417(.O (g34718), .I (I32884));
INVX1 gate5418(.O (g24985), .I (g23586));
INVX1 gate5419(.O (g34521), .I (g34270));
INVX1 gate5420(.O (g32730), .I (g31327));
INVX1 gate5421(.O (g23546), .I (g21611));
INVX1 gate5422(.O (I24215), .I (g22360));
INVX1 gate5423(.O (g32793), .I (g31021));
INVX1 gate5424(.O (I18653), .I (g5681));
INVX1 gate5425(.O (g20374), .I (g18065));
INVX1 gate5426(.O (g23211), .I (g21308));
INVX1 gate5427(.O (I30644), .I (g32024));
INVX1 gate5428(.O (g19882), .I (g16540));
INVX1 gate5429(.O (g19414), .I (g16349));
INVX1 gate5430(.O (g26701), .I (g25341));
INVX1 gate5431(.O (g7245), .I (I11896));
INVX1 gate5432(.O (g17580), .I (I18509));
INVX1 gate5433(.O (g11753), .I (g8587));
INVX1 gate5434(.O (I29961), .I (g30984));
INVX1 gate5435(.O (I12538), .I (g58));
INVX1 gate5436(.O (g26777), .I (g25439));
INVX1 gate5437(.O (g20643), .I (g15962));
INVX1 gate5438(.O (I18138), .I (g14277));
INVX1 gate5439(.O (g9049), .I (g640));
INVX1 gate5440(.O (g23088), .I (I22240));
INVX1 gate5441(.O (g31847), .I (g29385));
INVX1 gate5442(.O (g32765), .I (g31327));
INVX1 gate5443(.O (g19407), .I (g16268));
INVX1 gate5444(.O (g9449), .I (g5770));
INVX1 gate5445(.O (g16449), .I (I17679));
INVX1 gate5446(.O (g11031), .I (g8609));
INVX1 gate5447(.O (g22922), .I (g20330));
INVX1 gate5448(.O (g23860), .I (g19074));
INVX1 gate5449(.O (I15650), .I (g12110));
INVX1 gate5450(.O (g32690), .I (g31070));
INVX1 gate5451(.O (g9575), .I (g6509));
INVX1 gate5452(.O (g32549), .I (g31554));
INVX1 gate5453(.O (I15736), .I (g12322));
INVX1 gate5454(.O (I14684), .I (g7717));
INVX1 gate5455(.O (I18333), .I (g1083));
INVX1 gate5456(.O (g22179), .I (g19210));
INVX1 gate5457(.O (I29717), .I (g30931));
INVX1 gate5458(.O (g25262), .I (g22763));
INVX1 gate5459(.O (I11617), .I (g1));
INVX1 gate5460(.O (g11736), .I (g8165));
INVX1 gate5461(.O (g20669), .I (g15426));
INVX1 gate5462(.O (I17136), .I (g14398));
INVX1 gate5463(.O (g16897), .I (I18083));
INVX1 gate5464(.O (I26503), .I (g26811));
INVX1 gate5465(.O (g34573), .I (I32645));
INVX1 gate5466(.O (g7344), .I (g5659));
INVX1 gate5467(.O (g25899), .I (g24997));
INVX1 gate5468(.O (g13736), .I (g11313));
INVX1 gate5469(.O (g32548), .I (g30673));
INVX1 gate5470(.O (I18852), .I (g13716));
INVX1 gate5471(.O (I32687), .I (g34431));
INVX1 gate5472(.O (g34247), .I (I32240));
INVX1 gate5473(.O (I32976), .I (g34699));
INVX1 gate5474(.O (I32985), .I (g34736));
INVX1 gate5475(.O (g22178), .I (g19147));
INVX1 gate5476(.O (g9498), .I (g5101));
INVX1 gate5477(.O (g6873), .I (g3151));
INVX1 gate5478(.O (g20668), .I (g15426));
INVX1 gate5479(.O (g34926), .I (I33170));
INVX1 gate5480(.O (g32504), .I (g30673));
INVX1 gate5481(.O (g31851), .I (g29385));
INVX1 gate5482(.O (I15843), .I (g11181));
INVX1 gate5483(.O (I32752), .I (g34510));
INVX1 gate5484(.O (g9833), .I (g2449));
INVX1 gate5485(.O (g10287), .I (I13715));
INVX1 gate5486(.O (g7259), .I (g4375));
INVX1 gate5487(.O (g21659), .I (g17727));
INVX1 gate5488(.O (I33050), .I (g34777));
INVX1 gate5489(.O (g14314), .I (I16476));
INVX1 gate5490(.O (g16717), .I (g13951));
INVX1 gate5491(.O (g17531), .I (I18476));
INVX1 gate5492(.O (g12836), .I (g10351));
INVX1 gate5493(.O (g20195), .I (g16931));
INVX1 gate5494(.O (I26581), .I (g26942));
INVX1 gate5495(.O (g8997), .I (g577));
INVX1 gate5496(.O (g23987), .I (g19277));
INVX1 gate5497(.O (g10085), .I (g1768));
INVX1 gate5498(.O (g8541), .I (g3498));
INVX1 gate5499(.O (g23250), .I (g21070));
INVX1 gate5500(.O (g24489), .I (I23694));
INVX1 gate5501(.O (I23363), .I (g23385));
INVX1 gate5502(.O (g14307), .I (I16468));
INVX1 gate5503(.O (I27235), .I (g27320));
INVX1 gate5504(.O (g17178), .I (I18214));
INVX1 gate5505(.O (g6869), .I (I11691));
INVX1 gate5506(.O (g34777), .I (I32973));
INVX1 gate5507(.O (g12477), .I (I15295));
INVX1 gate5508(.O (g20525), .I (g17955));
INVX1 gate5509(.O (I15869), .I (g11234));
INVX1 gate5510(.O (g18939), .I (g16077));
INVX1 gate5511(.O (g8132), .I (I12411));
INVX1 gate5512(.O (g28443), .I (I26936));
INVX1 gate5513(.O (g34272), .I (g34229));
INVX1 gate5514(.O (g24525), .I (g22670));
INVX1 gate5515(.O (g24424), .I (g22722));
INVX1 gate5516(.O (I11623), .I (g28));
INVX1 gate5517(.O (g13132), .I (g10632));
INVX1 gate5518(.O (g17685), .I (I18662));
INVX1 gate5519(.O (g17676), .I (g12941));
INVX1 gate5520(.O (g13869), .I (g10831));
INVX1 gate5521(.O (g20558), .I (I20650));
INVX1 gate5522(.O (g8680), .I (g686));
INVX1 gate5523(.O (g22936), .I (g20283));
INVX1 gate5524(.O (I13623), .I (g4294));
INVX1 gate5525(.O (I21486), .I (g18727));
INVX1 gate5526(.O (g17953), .I (I18861));
INVX1 gate5527(.O (I22327), .I (g19367));
INVX1 gate5528(.O (g23339), .I (g21070));
INVX1 gate5529(.O (g8353), .I (I12530));
INVX1 gate5530(.O (g18938), .I (g16053));
INVX1 gate5531(.O (g23943), .I (g19147));
INVX1 gate5532(.O (g18093), .I (I18885));
INVX1 gate5533(.O (I13037), .I (g4304));
INVX1 gate5534(.O (I29149), .I (g29384));
INVX1 gate5535(.O (g14431), .I (g12208));
INVX1 gate5536(.O (g31213), .I (I29013));
INVX1 gate5537(.O (g11868), .I (g9185));
INVX1 gate5538(.O (g12864), .I (g10373));
INVX1 gate5539(.O (g13868), .I (g11493));
INVX1 gate5540(.O (g6917), .I (g3684));
INVX1 gate5541(.O (g8744), .I (g691));
INVX1 gate5542(.O (g23338), .I (g20453));
INVX1 gate5543(.O (g18065), .I (I18875));
INVX1 gate5544(.O (g24893), .I (I24060));
INVX1 gate5545(.O (g12749), .I (g7074));
INVX1 gate5546(.O (g19435), .I (g16449));
INVX1 gate5547(.O (g9162), .I (g622));
INVX1 gate5548(.O (g9019), .I (I12950));
INVX1 gate5549(.O (g17417), .I (g14804));
INVX1 gate5550(.O (I18609), .I (g5976));
INVX1 gate5551(.O (g7886), .I (g1442));
INVX1 gate5552(.O (g20544), .I (g15171));
INVX1 gate5553(.O (g23969), .I (g19277));
INVX1 gate5554(.O (g32626), .I (g30614));
INVX1 gate5555(.O (g28039), .I (g26365));
INVX1 gate5556(.O (I32195), .I (g33628));
INVX1 gate5557(.O (I13352), .I (g4146));
INVX1 gate5558(.O (g11709), .I (I14584));
INVX1 gate5559(.O (g30997), .I (g29702));
INVX1 gate5560(.O (g10156), .I (g2675));
INVX1 gate5561(.O (g20713), .I (g15277));
INVX1 gate5562(.O (g21060), .I (g15509));
INVX1 gate5563(.O (g34997), .I (I33291));
INVX1 gate5564(.O (I12991), .I (g6752));
INVX1 gate5565(.O (g23060), .I (g19908));
INVX1 gate5566(.O (g23968), .I (g18833));
INVX1 gate5567(.O (g18875), .I (g15171));
INVX1 gate5568(.O (g32533), .I (g30614));
INVX1 gate5569(.O (g8558), .I (g3787));
INVX1 gate5570(.O (g28038), .I (g26365));
INVX1 gate5571(.O (I32525), .I (g34285));
INVX1 gate5572(.O (g13259), .I (I15824));
INVX1 gate5573(.O (g33912), .I (I31770));
INVX1 gate5574(.O (g19744), .I (g15885));
INVX1 gate5575(.O (g16620), .I (I17808));
INVX1 gate5576(.O (g7314), .I (g1740));
INVX1 gate5577(.O (g10180), .I (g2259));
INVX1 gate5578(.O (I14006), .I (g9104));
INVX1 gate5579(.O (I17108), .I (g13782));
INVX1 gate5580(.O (I14475), .I (g10175));
INVX1 gate5581(.O (g11471), .I (g7626));
INVX1 gate5582(.O (g19345), .I (g17591));
INVX1 gate5583(.O (g25099), .I (g22369));
INVX1 gate5584(.O (g13087), .I (g12012));
INVX1 gate5585(.O (g32775), .I (g30825));
INVX1 gate5586(.O (g25388), .I (g22763));
INVX1 gate5587(.O (g25324), .I (g22228));
INVX1 gate5588(.O (I14727), .I (g7753));
INVX1 gate5589(.O (g13258), .I (I15821));
INVX1 gate5590(.O (g12900), .I (g10406));
INVX1 gate5591(.O (g19399), .I (g16489));
INVX1 gate5592(.O (g20610), .I (g18008));
INVX1 gate5593(.O (g7870), .I (g1193));
INVX1 gate5594(.O (g21411), .I (g15426));
INVX1 gate5595(.O (g17762), .I (g13000));
INVX1 gate5596(.O (g20705), .I (I20793));
INVX1 gate5597(.O (g34766), .I (g34703));
INVX1 gate5598(.O (g23870), .I (g21293));
INVX1 gate5599(.O (I16010), .I (g11148));
INVX1 gate5600(.O (g23411), .I (g20734));
INVX1 gate5601(.O (g23527), .I (g21611));
INVX1 gate5602(.O (g28187), .I (I26710));
INVX1 gate5603(.O (I14222), .I (g8286));
INVX1 gate5604(.O (I21922), .I (g21335));
INVX1 gate5605(.O (g25534), .I (g22763));
INVX1 gate5606(.O (g15932), .I (I17395));
INVX1 gate5607(.O (g25098), .I (g22369));
INVX1 gate5608(.O (g10335), .I (g4483));
INVX1 gate5609(.O (I23321), .I (g21693));
INVX1 gate5610(.O (g7650), .I (g4064));
INVX1 gate5611(.O (g27101), .I (g26770));
INVX1 gate5612(.O (g25272), .I (g23715));
INVX1 gate5613(.O (g29862), .I (g28406));
INVX1 gate5614(.O (g24042), .I (g20014));
INVX1 gate5615(.O (g33072), .I (g31945));
INVX1 gate5616(.O (g20189), .I (I20447));
INVX1 gate5617(.O (g19398), .I (g16489));
INVX1 gate5618(.O (g20679), .I (g15634));
INVX1 gate5619(.O (I29368), .I (g30321));
INVX1 gate5620(.O (g17423), .I (I18360));
INVX1 gate5621(.O (g16971), .I (I18131));
INVX1 gate5622(.O (g11043), .I (g8561));
INVX1 gate5623(.O (g12036), .I (g9245));
INVX1 gate5624(.O (g9086), .I (g847));
INVX1 gate5625(.O (g32737), .I (g31327));
INVX1 gate5626(.O (I18813), .I (g5673));
INVX1 gate5627(.O (g17216), .I (g14454));
INVX1 gate5628(.O (g20270), .I (g15277));
INVX1 gate5629(.O (g9728), .I (g5109));
INVX1 gate5630(.O (g19652), .I (g16897));
INVX1 gate5631(.O (I30986), .I (g32437));
INVX1 gate5632(.O (I17750), .I (g14383));
INVX1 gate5633(.O (g22543), .I (g19801));
INVX1 gate5634(.O (g17587), .I (I18518));
INVX1 gate5635(.O (g9730), .I (g5436));
INVX1 gate5636(.O (I31504), .I (g33164));
INVX1 gate5637(.O (g24124), .I (g21209));
INVX1 gate5638(.O (g8092), .I (g1589));
INVX1 gate5639(.O (g14694), .I (I16795));
INVX1 gate5640(.O (g29948), .I (g28853));
INVX1 gate5641(.O (g8492), .I (g3396));
INVX1 gate5642(.O (g9185), .I (I13007));
INVX1 gate5643(.O (g23503), .I (g21468));
INVX1 gate5644(.O (g23894), .I (g19074));
INVX1 gate5645(.O (g19263), .I (I19799));
INVX1 gate5646(.O (g32697), .I (g31070));
INVX1 gate5647(.O (g27064), .I (I25786));
INVX1 gate5648(.O (I18674), .I (g13101));
INVX1 gate5649(.O (g25032), .I (g23639));
INVX1 gate5650(.O (g20383), .I (g15373));
INVX1 gate5651(.O (g32856), .I (g31021));
INVX1 gate5652(.O (I28913), .I (g30322));
INVX1 gate5653(.O (g11810), .I (g9664));
INVX1 gate5654(.O (g25140), .I (g22228));
INVX1 gate5655(.O (g9070), .I (g5428));
INVX1 gate5656(.O (g8714), .I (g4859));
INVX1 gate5657(.O (g7594), .I (I12064));
INVX1 gate5658(.O (g31820), .I (g29385));
INVX1 gate5659(.O (g10487), .I (g10233));
INVX1 gate5660(.O (g32880), .I (g30614));
INVX1 gate5661(.O (g13068), .I (I15697));
INVX1 gate5662(.O (g25997), .I (I25095));
INVX1 gate5663(.O (g7972), .I (g1046));
INVX1 gate5664(.O (g24030), .I (g21127));
INVX1 gate5665(.O (g20267), .I (g17955));
INVX1 gate5666(.O (g24093), .I (g20998));
INVX1 gate5667(.O (g10502), .I (g8876));
INVX1 gate5668(.O (g26776), .I (g25498));
INVX1 gate5669(.O (g23714), .I (g20751));
INVX1 gate5670(.O (I27758), .I (g28119));
INVX1 gate5671(.O (g23450), .I (I22571));
INVX1 gate5672(.O (I29228), .I (g30314));
INVX1 gate5673(.O (g32512), .I (g31566));
INVX1 gate5674(.O (g7806), .I (g4681));
INVX1 gate5675(.O (I15878), .I (g11249));
INVX1 gate5676(.O (g20065), .I (g16846));
INVX1 gate5677(.O (g31846), .I (g29385));
INVX1 gate5678(.O (g7943), .I (g1395));
INVX1 gate5679(.O (g24065), .I (g20982));
INVX1 gate5680(.O (g11878), .I (I14690));
INVX1 gate5681(.O (g19361), .I (I19843));
INVX1 gate5682(.O (I20609), .I (g16539));
INVX1 gate5683(.O (I12758), .I (g4093));
INVX1 gate5684(.O (g23819), .I (g19147));
INVX1 gate5685(.O (g12874), .I (g10383));
INVX1 gate5686(.O (g26754), .I (g25300));
INVX1 gate5687(.O (g34472), .I (I32525));
INVX1 gate5688(.O (g25766), .I (g24439));
INVX1 gate5689(.O (g28479), .I (g27654));
INVX1 gate5690(.O (I32678), .I (g34428));
INVX1 gate5691(.O (g23202), .I (I22302));
INVX1 gate5692(.O (g14443), .I (I16596));
INVX1 gate5693(.O (g23257), .I (g20924));
INVX1 gate5694(.O (g26859), .I (I25591));
INVX1 gate5695(.O (g27009), .I (g25911));
INVX1 gate5696(.O (g26825), .I (I25541));
INVX1 gate5697(.O (g21055), .I (g15224));
INVX1 gate5698(.O (g23496), .I (g20248));
INVX1 gate5699(.O (g7322), .I (g1862));
INVX1 gate5700(.O (g16228), .I (I17569));
INVX1 gate5701(.O (g20219), .I (I20495));
INVX1 gate5702(.O (g23055), .I (g20887));
INVX1 gate5703(.O (g6990), .I (g4742));
INVX1 gate5704(.O (g17242), .I (g14454));
INVX1 gate5705(.O (g34246), .I (I32237));
INVX1 gate5706(.O (g10278), .I (g4628));
INVX1 gate5707(.O (g33413), .I (g31971));
INVX1 gate5708(.O (g29847), .I (g28395));
INVX1 gate5709(.O (I29582), .I (g30591));
INVX1 gate5710(.O (g23111), .I (g20391));
INVX1 gate5711(.O (g12009), .I (I14862));
INVX1 gate5712(.O (g21070), .I (I20937));
INVX1 gate5713(.O (g6888), .I (I11701));
INVX1 gate5714(.O (g22974), .I (g20330));
INVX1 gate5715(.O (g32831), .I (g31376));
INVX1 gate5716(.O (g33691), .I (I31528));
INVX1 gate5717(.O (g32445), .I (I29973));
INVX1 gate5718(.O (I32938), .I (g34663));
INVX1 gate5719(.O (I32093), .I (g33670));
INVX1 gate5720(.O (I13276), .I (g5798));
INVX1 gate5721(.O (g16716), .I (g13948));
INVX1 gate5722(.O (g9678), .I (g5406));
INVX1 gate5723(.O (g10039), .I (g2273));
INVX1 gate5724(.O (g10306), .I (I13726));
INVX1 gate5725(.O (g32499), .I (g31376));
INVX1 gate5726(.O (g23986), .I (g18833));
INVX1 gate5727(.O (g30591), .I (I28851));
INVX1 gate5728(.O (g6956), .I (g4242));
INVX1 gate5729(.O (g18984), .I (g17486));
INVX1 gate5730(.O (g8623), .I (g3990));
INVX1 gate5731(.O (I11809), .I (g6741));
INVX1 gate5732(.O (g34591), .I (I32681));
INVX1 gate5733(.O (I18214), .I (g12918));
INVX1 gate5734(.O (g12892), .I (g10398));
INVX1 gate5735(.O (g34785), .I (I32985));
INVX1 gate5736(.O (g16582), .I (g13915));
INVX1 gate5737(.O (g17772), .I (g14297));
INVX1 gate5738(.O (g34776), .I (I32970));
INVX1 gate5739(.O (g11425), .I (g7640));
INVX1 gate5740(.O (g10038), .I (g2241));
INVX1 gate5741(.O (g32498), .I (g31566));
INVX1 gate5742(.O (g23384), .I (I22485));
INVX1 gate5743(.O (g17639), .I (I18600));
INVX1 gate5744(.O (I12141), .I (g599));
INVX1 gate5745(.O (g34147), .I (g33823));
INVX1 gate5746(.O (g9682), .I (I13280));
INVX1 gate5747(.O (g9766), .I (g2748));
INVX1 gate5748(.O (g15811), .I (g13125));
INVX1 gate5749(.O (g16310), .I (g13223));
INVX1 gate5750(.O (g7096), .I (g6537));
INVX1 gate5751(.O (g10815), .I (g9917));
INVX1 gate5752(.O (g13458), .I (g11048));
INVX1 gate5753(.O (g24160), .I (I23324));
INVX1 gate5754(.O (I15918), .I (g12381));
INVX1 gate5755(.O (g9305), .I (g5381));
INVX1 gate5756(.O (g7496), .I (g5969));
INVX1 gate5757(.O (g33929), .I (I31803));
INVX1 gate5758(.O (g16627), .I (I17819));
INVX1 gate5759(.O (g17638), .I (g14838));
INVX1 gate5760(.O (g22841), .I (g20391));
INVX1 gate5761(.O (g34950), .I (g34940));
INVX1 gate5762(.O (g12914), .I (g12235));
INVX1 gate5763(.O (g13010), .I (I15620));
INVX1 gate5764(.O (g32611), .I (g31154));
INVX1 gate5765(.O (g7845), .I (g1146));
INVX1 gate5766(.O (I33232), .I (g34957));
INVX1 gate5767(.O (g25451), .I (g22228));
INVX1 gate5768(.O (g32722), .I (g30937));
INVX1 gate5769(.O (g25220), .I (I24396));
INVX1 gate5770(.O (g32924), .I (g30937));
INVX1 gate5771(.O (g33928), .I (I31800));
INVX1 gate5772(.O (g19947), .I (g17226));
INVX1 gate5773(.O (g7195), .I (g25));
INVX1 gate5774(.O (g12907), .I (g10415));
INVX1 gate5775(.O (g20617), .I (g15277));
INVX1 gate5776(.O (g17416), .I (g14956));
INVX1 gate5777(.O (g7395), .I (g6005));
INVX1 gate5778(.O (g7891), .I (g2994));
INVX1 gate5779(.O (g8651), .I (g758));
INVX1 gate5780(.O (g16958), .I (g14238));
INVX1 gate5781(.O (g9748), .I (g114));
INVX1 gate5782(.O (g13545), .I (I16010));
INVX1 gate5783(.O (g23877), .I (g19147));
INVX1 gate5784(.O (g19273), .I (g16100));
INVX1 gate5785(.O (g20915), .I (I20882));
INVX1 gate5786(.O (g7913), .I (g1052));
INVX1 gate5787(.O (g27074), .I (I25790));
INVX1 gate5788(.O (g28321), .I (g27317));
INVX1 gate5789(.O (I32837), .I (g34498));
INVX1 gate5790(.O (g30996), .I (g29694));
INVX1 gate5791(.O (g25246), .I (g23828));
INVX1 gate5792(.O (g34151), .I (I32106));
INVX1 gate5793(.O (I12135), .I (g807));
INVX1 gate5794(.O (g10143), .I (g568));
INVX1 gate5795(.O (g29213), .I (I27555));
INVX1 gate5796(.O (g34996), .I (I33288));
INVX1 gate5797(.O (g23019), .I (g19866));
INVX1 gate5798(.O (I33261), .I (g34977));
INVX1 gate5799(.O (g8285), .I (I12497));
INVX1 gate5800(.O (g12074), .I (I14932));
INVX1 gate5801(.O (I25695), .I (g25690));
INVX1 gate5802(.O (g9226), .I (g1564));
INVX1 gate5803(.O (g20277), .I (g16487));
INVX1 gate5804(.O (g16603), .I (I17787));
INVX1 gate5805(.O (g16742), .I (g13983));
INVX1 gate5806(.O (g23196), .I (g20785));
INVX1 gate5807(.O (g34844), .I (g34737));
INVX1 gate5808(.O (I22564), .I (g20857));
INVX1 gate5809(.O (g16096), .I (g13530));
INVX1 gate5810(.O (g23018), .I (g19801));
INVX1 gate5811(.O (g32753), .I (g30735));
INVX1 gate5812(.O (g12238), .I (I15102));
INVX1 gate5813(.O (g32461), .I (g30614));
INVX1 gate5814(.O (I21242), .I (g16540));
INVX1 gate5815(.O (g10169), .I (g6395));
INVX1 gate5816(.O (g24075), .I (g19935));
INVX1 gate5817(.O (g17579), .I (g14959));
INVX1 gate5818(.O (g19371), .I (I19857));
INVX1 gate5819(.O (g20595), .I (g15877));
INVX1 gate5820(.O (g23526), .I (g21611));
INVX1 gate5821(.O (g6808), .I (g554));
INVX1 gate5822(.O (g20494), .I (g17847));
INVX1 gate5823(.O (g14169), .I (g12381));
INVX1 gate5824(.O (g8139), .I (g1648));
INVX1 gate5825(.O (I16289), .I (g12107));
INVX1 gate5826(.O (I32455), .I (g34242));
INVX1 gate5827(.O (g7266), .I (g35));
INVX1 gate5828(.O (g29912), .I (g28827));
INVX1 gate5829(.O (g29311), .I (g28998));
INVX1 gate5830(.O (g10410), .I (g7069));
INVX1 gate5831(.O (g20623), .I (g17929));
INVX1 gate5832(.O (g27675), .I (I26309));
INVX1 gate5833(.O (I12049), .I (g781));
INVX1 gate5834(.O (g9373), .I (g5142));
INVX1 gate5835(.O (g17014), .I (g14297));
INVX1 gate5836(.O (g27092), .I (g26737));
INVX1 gate5837(.O (g9091), .I (g1430));
INVX1 gate5838(.O (g20037), .I (g17328));
INVX1 gate5839(.O (g31827), .I (g29385));
INVX1 gate5840(.O (g32736), .I (g30937));
INVX1 gate5841(.O (I32617), .I (g34333));
INVX1 gate5842(.O (g13322), .I (g10918));
INVX1 gate5843(.O (g32887), .I (g30614));
INVX1 gate5844(.O (I32470), .I (g34247));
INVX1 gate5845(.O (g24623), .I (g23076));
INVX1 gate5846(.O (g33827), .I (I31672));
INVX1 gate5847(.O (g9491), .I (g2729));
INVX1 gate5848(.O (I14905), .I (g9822));
INVX1 gate5849(.O (g24037), .I (g21127));
INVX1 gate5850(.O (g34420), .I (g34152));
INVX1 gate5851(.O (g16429), .I (I17671));
INVX1 gate5852(.O (I11665), .I (g1589));
INVX1 gate5853(.O (g20782), .I (g15853));
INVX1 gate5854(.O (g21457), .I (g17367));
INVX1 gate5855(.O (g13901), .I (g11480));
INVX1 gate5856(.O (g23402), .I (g20875));
INVX1 gate5857(.O (I13166), .I (g5101));
INVX1 gate5858(.O (g32529), .I (g30735));
INVX1 gate5859(.O (g23457), .I (I22580));
INVX1 gate5860(.O (g25370), .I (g22228));
INVX1 gate5861(.O (g8795), .I (I12793));
INVX1 gate5862(.O (g10363), .I (I13779));
INVX1 gate5863(.O (I24400), .I (g23954));
INVX1 gate5864(.O (g10217), .I (g2102));
INVX1 gate5865(.O (I14593), .I (g9978));
INVX1 gate5866(.O (g30318), .I (g28274));
INVX1 gate5867(.O (g14363), .I (I16521));
INVX1 gate5868(.O (g14217), .I (I16417));
INVX1 gate5869(.O (g9283), .I (g1736));
INVX1 gate5870(.O (I14346), .I (g10233));
INVX1 gate5871(.O (g16428), .I (I17668));
INVX1 gate5872(.O (g9369), .I (g5084));
INVX1 gate5873(.O (g32528), .I (g31554));
INVX1 gate5874(.O (g32696), .I (g30825));
INVX1 gate5875(.O (g9007), .I (g1083));
INVX1 gate5876(.O (I21230), .I (g16540));
INVX1 gate5877(.O (g32843), .I (g31021));
INVX1 gate5878(.O (g6957), .I (g2932));
INVX1 gate5879(.O (g24419), .I (g22722));
INVX1 gate5880(.O (g32393), .I (g30922));
INVX1 gate5881(.O (g9407), .I (g6549));
INVX1 gate5882(.O (I15295), .I (g8515));
INVX1 gate5883(.O (I11892), .I (g4408));
INVX1 gate5884(.O (g34059), .I (g33658));
INVX1 gate5885(.O (g8672), .I (g4669));
INVX1 gate5886(.O (g9920), .I (g4322));
INVX1 gate5887(.O (I15144), .I (g5659));
INVX1 gate5888(.O (I13892), .I (g1576));
INVX1 gate5889(.O (g31803), .I (g29385));
INVX1 gate5890(.O (g32764), .I (g30937));
INVX1 gate5891(.O (g24155), .I (I23309));
INVX1 gate5892(.O (g24418), .I (g22722));
INVX1 gate5893(.O (I32467), .I (g34246));
INVX1 gate5894(.O (g20266), .I (g17873));
INVX1 gate5895(.O (g8477), .I (g3061));
INVX1 gate5896(.O (g34540), .I (I32607));
INVX1 gate5897(.O (g11823), .I (I14647));
INVX1 gate5898(.O (g13680), .I (I16077));
INVX1 gate5899(.O (g17615), .I (I18574));
INVX1 gate5900(.O (g12883), .I (g10390));
INVX1 gate5901(.O (g13144), .I (I15773));
INVX1 gate5902(.O (g22493), .I (g19801));
INVX1 gate5903(.O (g7097), .I (I11809));
INVX1 gate5904(.O (g23001), .I (g19801));
INVX1 gate5905(.O (g34058), .I (g33660));
INVX1 gate5906(.O (g24170), .I (I23354));
INVX1 gate5907(.O (g32869), .I (g30735));
INVX1 gate5908(.O (I18882), .I (g16580));
INVX1 gate5909(.O (g32960), .I (g31327));
INVX1 gate5910(.O (I18414), .I (g14359));
INVX1 gate5911(.O (g7497), .I (g6358));
INVX1 gate5912(.O (I14797), .I (g9636));
INVX1 gate5913(.O (g19421), .I (g16326));
INVX1 gate5914(.O (g17720), .I (g15045));
INVX1 gate5915(.O (I33056), .I (g34778));
INVX1 gate5916(.O (I25689), .I (g25688));
INVX1 gate5917(.O (g9582), .I (g703));
INVX1 gate5918(.O (g11336), .I (g7620));
INVX1 gate5919(.O (g7960), .I (g1404));
INVX1 gate5920(.O (g32868), .I (g31376));
INVX1 gate5921(.O (g8205), .I (g2208));
INVX1 gate5922(.O (I32782), .I (g34571));
INVX1 gate5923(.O (g10223), .I (g4561));
INVX1 gate5924(.O (g21689), .I (I21250));
INVX1 gate5925(.O (g23256), .I (g20785));
INVX1 gate5926(.O (I12106), .I (g626));
INVX1 gate5927(.O (I12605), .I (g1570));
INVX1 gate5928(.O (g17430), .I (I18373));
INVX1 gate5929(.O (g17746), .I (g14825));
INVX1 gate5930(.O (g20853), .I (g15595));
INVX1 gate5931(.O (g34044), .I (g33675));
INVX1 gate5932(.O (g21280), .I (g16601));
INVX1 gate5933(.O (g23923), .I (g18997));
INVX1 gate5934(.O (I14409), .I (g8364));
INVX1 gate5935(.O (g29152), .I (g27907));
INVX1 gate5936(.O (g29846), .I (g28391));
INVX1 gate5937(.O (I32352), .I (g34169));
INVX1 gate5938(.O (I29002), .I (g29675));
INVX1 gate5939(.O (g21300), .I (I21047));
INVX1 gate5940(.O (g20167), .I (g16971));
INVX1 gate5941(.O (g20194), .I (g16897));
INVX1 gate5942(.O (g20589), .I (g15224));
INVX1 gate5943(.O (g32709), .I (g30735));
INVX1 gate5944(.O (g11966), .I (I14800));
INVX1 gate5945(.O (g23300), .I (g20283));
INVX1 gate5946(.O (I12463), .I (g4812));
INVX1 gate5947(.O (g17465), .I (g12955));
INVX1 gate5948(.O (g8742), .I (g4035));
INVX1 gate5949(.O (g13966), .I (I16246));
INVX1 gate5950(.O (g10084), .I (g2837));
INVX1 gate5951(.O (g24167), .I (I23345));
INVX1 gate5952(.O (g9415), .I (g2169));
INVX1 gate5953(.O (g19541), .I (g16136));
INVX1 gate5954(.O (g30301), .I (I28548));
INVX1 gate5955(.O (g10110), .I (g661));
INVX1 gate5956(.O (g11631), .I (g8595));
INVX1 gate5957(.O (g19473), .I (g16349));
INVX1 gate5958(.O (g18101), .I (I18909));
INVX1 gate5959(.O (g11017), .I (g10289));
INVX1 gate5960(.O (g20588), .I (g18008));
INVX1 gate5961(.O (g20524), .I (g17873));
INVX1 gate5962(.O (g32708), .I (g31376));
INVX1 gate5963(.O (I32170), .I (g33638));
INVX1 gate5964(.O (I12033), .I (g776));
INVX1 gate5965(.O (g13017), .I (I15633));
INVX1 gate5966(.O (I28174), .I (g28803));
INVX1 gate5967(.O (I29245), .I (g29491));
INVX1 gate5968(.O (g32471), .I (g31376));
INVX1 gate5969(.O (g19789), .I (g17015));
INVX1 gate5970(.O (g24524), .I (g22876));
INVX1 gate5971(.O (g24836), .I (I24008));
INVX1 gate5972(.O (g16129), .I (I17488));
INVX1 gate5973(.O (g25227), .I (g22763));
INVX1 gate5974(.O (g14321), .I (g10874));
INVX1 gate5975(.O (g34739), .I (I32909));
INVX1 gate5976(.O (g10531), .I (g8925));
INVX1 gate5977(.O (g17684), .I (g15036));
INVX1 gate5978(.O (g27438), .I (I26130));
INVX1 gate5979(.O (g14179), .I (g11048));
INVX1 gate5980(.O (g25025), .I (g22498));
INVX1 gate5981(.O (g7267), .I (g1604));
INVX1 gate5982(.O (g24477), .I (I23680));
INVX1 gate5983(.O (g10178), .I (g2126));
INVX1 gate5984(.O (g26632), .I (g25473));
INVX1 gate5985(.O (g24119), .I (g19935));
INVX1 gate5986(.O (g27349), .I (g26352));
INVX1 gate5987(.O (I31650), .I (g33212));
INVX1 gate5988(.O (g23066), .I (g20330));
INVX1 gate5989(.O (I28390), .I (g29185));
INVX1 gate5990(.O (g9721), .I (g5097));
INVX1 gate5991(.O (g23231), .I (g20050));
INVX1 gate5992(.O (g34699), .I (I32855));
INVX1 gate5993(.O (g19434), .I (g16326));
INVX1 gate5994(.O (g16626), .I (g14133));
INVX1 gate5995(.O (g8273), .I (g2453));
INVX1 gate5996(.O (g10685), .I (I13995));
INVX1 gate5997(.O (I16489), .I (g12793));
INVX1 gate5998(.O (g16323), .I (I17653));
INVX1 gate5999(.O (g24118), .I (g19890));
INVX1 gate6000(.O (g10373), .I (g6917));
INVX1 gate6001(.O (g14186), .I (g11346));
INVX1 gate6002(.O (g14676), .I (I16775));
INVX1 gate6003(.O (g24022), .I (g20982));
INVX1 gate6004(.O (g34698), .I (g34550));
INVX1 gate6005(.O (g7293), .I (g4452));
INVX1 gate6006(.O (g12906), .I (g10413));
INVX1 gate6007(.O (g16533), .I (I17733));
INVX1 gate6008(.O (g20616), .I (g15277));
INVX1 gate6009(.O (I18114), .I (g14509));
INVX1 gate6010(.O (g23876), .I (g19074));
INVX1 gate6011(.O (I18758), .I (g6719));
INVX1 gate6012(.O (g13023), .I (g11897));
INVX1 gate6013(.O (g18874), .I (g15938));
INVX1 gate6014(.O (I31528), .I (g33219));
INVX1 gate6015(.O (g25044), .I (g23675));
INVX1 gate6016(.O (I19661), .I (g17587));
INVX1 gate6017(.O (g29929), .I (g28914));
INVX1 gate6018(.O (g16775), .I (I17999));
INVX1 gate6019(.O (I18107), .I (g4019));
INVX1 gate6020(.O (g10417), .I (g7117));
INVX1 gate6021(.O (I25511), .I (g25073));
INVX1 gate6022(.O (g32602), .I (g30825));
INVX1 gate6023(.O (g32810), .I (g31376));
INVX1 gate6024(.O (I13637), .I (g102));
INVX1 gate6025(.O (I20882), .I (g17619));
INVX1 gate6026(.O (g32657), .I (g31528));
INVX1 gate6027(.O (g32774), .I (g30735));
INVX1 gate6028(.O (g33778), .I (I31625));
INVX1 gate6029(.O (g7828), .I (g4871));
INVX1 gate6030(.O (g32955), .I (g30735));
INVX1 gate6031(.O (g21511), .I (g15483));
INVX1 gate6032(.O (g29928), .I (g28871));
INVX1 gate6033(.O (I26670), .I (g27709));
INVX1 gate6034(.O (g20704), .I (g15373));
INVX1 gate6035(.O (g23511), .I (I22640));
INVX1 gate6036(.O (g34427), .I (I32452));
INVX1 gate6037(.O (I32119), .I (g33648));
INVX1 gate6038(.O (g32879), .I (g31327));
INVX1 gate6039(.O (g8572), .I (I12654));
INVX1 gate6040(.O (g20053), .I (g17328));
INVX1 gate6041(.O (g32970), .I (g30825));
INVX1 gate6042(.O (g10334), .I (g4420));
INVX1 gate6043(.O (g19682), .I (g17015));
INVX1 gate6044(.O (I14537), .I (g10106));
INVX1 gate6045(.O (g24053), .I (g21256));
INVX1 gate6046(.O (g25120), .I (g22432));
INVX1 gate6047(.O (I17780), .I (g13303));
INVX1 gate6048(.O (g17523), .I (g14732));
INVX1 gate6049(.O (g20900), .I (I20864));
INVX1 gate6050(.O (g8712), .I (I12712));
INVX1 gate6051(.O (g7592), .I (g347));
INVX1 gate6052(.O (I16544), .I (g11931));
INVX1 gate6053(.O (I18849), .I (g14290));
INVX1 gate6054(.O (g18008), .I (I18868));
INVX1 gate6055(.O (g32878), .I (g30937));
INVX1 gate6056(.O (g31945), .I (g31189));
INVX1 gate6057(.O (g21660), .I (g17694));
INVX1 gate6058(.O (g24466), .I (I23671));
INVX1 gate6059(.O (I16713), .I (g5331));
INVX1 gate6060(.O (g9689), .I (g124));
INVX1 gate6061(.O (g10762), .I (g8470));
INVX1 gate6062(.O (g25562), .I (g22763));
INVX1 gate6063(.O (g18892), .I (g15680));
INVX1 gate6064(.O (g20036), .I (g17433));
INVX1 gate6065(.O (g31826), .I (g29385));
INVX1 gate6066(.O (g32886), .I (g31327));
INVX1 gate6067(.O (I33161), .I (g34894));
INVX1 gate6068(.O (I18398), .I (g13745));
INVX1 gate6069(.O (g20101), .I (g17533));
INVX1 gate6070(.O (g24036), .I (g20982));
INVX1 gate6071(.O (I12541), .I (g194));
INVX1 gate6072(.O (g20560), .I (g17328));
INVX1 gate6073(.O (g16856), .I (I18048));
INVX1 gate6074(.O (g21456), .I (g15509));
INVX1 gate6075(.O (I26667), .I (g27585));
INVX1 gate6076(.O (g11985), .I (I14827));
INVX1 gate6077(.O (g17475), .I (I18398));
INVX1 gate6078(.O (g24101), .I (g20998));
INVX1 gate6079(.O (I23684), .I (g23230));
INVX1 gate6080(.O (g32792), .I (g31710));
INVX1 gate6081(.O (g23456), .I (g21514));
INVX1 gate6082(.O (g13976), .I (g11130));
INVX1 gate6083(.O (g24177), .I (I23375));
INVX1 gate6084(.O (g24560), .I (g22942));
INVX1 gate6085(.O (I15954), .I (g12381));
INVX1 gate6086(.O (g32967), .I (g31327));
INVX1 gate6087(.O (g10216), .I (I13684));
INVX1 gate6088(.O (g14423), .I (I16579));
INVX1 gate6089(.O (g8534), .I (g3338));
INVX1 gate6090(.O (I16610), .I (g10981));
INVX1 gate6091(.O (g9671), .I (g5134));
INVX1 gate6092(.O (g20642), .I (g15277));
INVX1 gate6093(.O (g23480), .I (I22601));
INVX1 gate6094(.O (g27415), .I (g26382));
INVX1 gate6095(.O (I20584), .I (g16587));
INVX1 gate6096(.O (g23916), .I (g19277));
INVX1 gate6097(.O (g9030), .I (g4793));
INVX1 gate6098(.O (g19760), .I (g17015));
INVX1 gate6099(.O (I32305), .I (g34209));
INVX1 gate6100(.O (I14381), .I (g8300));
INVX1 gate6101(.O (g16512), .I (g14015));
INVX1 gate6102(.O (I16679), .I (g12039));
INVX1 gate6103(.O (g23550), .I (g20248));
INVX1 gate6104(.O (g26784), .I (g25341));
INVX1 gate6105(.O (g9247), .I (g1559));
INVX1 gate6106(.O (I33258), .I (g34976));
INVX1 gate6107(.O (I32809), .I (g34586));
INVX1 gate6108(.O (g18907), .I (g15979));
INVX1 gate6109(.O (g7624), .I (I12106));
INVX1 gate6110(.O (g32459), .I (g31070));
INVX1 gate6111(.O (g20064), .I (g17533));
INVX1 gate6112(.O (g7953), .I (g4966));
INVX1 gate6113(.O (g30572), .I (g29945));
INVX1 gate6114(.O (g24064), .I (g20841));
INVX1 gate6115(.O (g28579), .I (g27714));
INVX1 gate6116(.O (g9564), .I (g6120));
INVX1 gate6117(.O (I18135), .I (g13144));
INVX1 gate6118(.O (g23307), .I (g20924));
INVX1 gate6119(.O (g32919), .I (g30735));
INVX1 gate6120(.O (g23085), .I (g19957));
INVX1 gate6121(.O (g32458), .I (g30825));
INVX1 gate6122(.O (I24759), .I (g24229));
INVX1 gate6123(.O (g14543), .I (I16660));
INVX1 gate6124(.O (g33932), .I (I31810));
INVX1 gate6125(.O (g9826), .I (g1844));
INVX1 gate6126(.O (g10117), .I (g2509));
INVX1 gate6127(.O (g10000), .I (g6151));
INVX1 gate6128(.O (g26824), .I (g25298));
INVX1 gate6129(.O (I16460), .I (g10430));
INVX1 gate6130(.O (g20874), .I (g15680));
INVX1 gate6131(.O (g21054), .I (g15373));
INVX1 gate6132(.O (g32918), .I (g31327));
INVX1 gate6133(.O (g23243), .I (g21070));
INVX1 gate6134(.O (g20630), .I (g17955));
INVX1 gate6135(.O (g11842), .I (I14660));
INVX1 gate6136(.O (g21431), .I (g18065));
INVX1 gate6137(.O (g9741), .I (I13317));
INVX1 gate6138(.O (g8903), .I (g1075));
INVX1 gate6139(.O (g23431), .I (g21514));
INVX1 gate6140(.O (I13906), .I (g7620));
INVX1 gate6141(.O (g32545), .I (g31070));
INVX1 gate6142(.O (g9910), .I (g2108));
INVX1 gate6143(.O (g17600), .I (g14659));
INVX1 gate6144(.O (I19671), .I (g15932));
INVX1 gate6145(.O (g34490), .I (I32547));
INVX1 gate6146(.O (g20166), .I (g16886));
INVX1 gate6147(.O (g20009), .I (g16349));
INVX1 gate6148(.O (I22583), .I (g20998));
INVX1 gate6149(.O (g27576), .I (g26081));
INVX1 gate6150(.O (g27585), .I (g25994));
INVX1 gate6151(.O (g20665), .I (g15373));
INVX1 gate6152(.O (g25547), .I (g22550));
INVX1 gate6153(.O (g32599), .I (g30673));
INVX1 gate6154(.O (I20744), .I (g17141));
INVX1 gate6155(.O (I31810), .I (g33164));
INVX1 gate6156(.O (g9638), .I (g1620));
INVX1 gate6157(.O (g21269), .I (g15506));
INVX1 gate6158(.O (g24166), .I (I23342));
INVX1 gate6159(.O (g24665), .I (g23067));
INVX1 gate6160(.O (g7716), .I (g1199));
INVX1 gate6161(.O (g7149), .I (g4564));
INVX1 gate6162(.O (g34784), .I (I32982));
INVX1 gate6163(.O (g7349), .I (g1270));
INVX1 gate6164(.O (g30297), .I (g28758));
INVX1 gate6165(.O (g27554), .I (g26625));
INVX1 gate6166(.O (g20008), .I (g16449));
INVX1 gate6167(.O (g34956), .I (I33214));
INVX1 gate6168(.O (g17952), .I (I18858));
INVX1 gate6169(.O (g32598), .I (g30614));
INVX1 gate6170(.O (g13016), .I (g11878));
INVX1 gate6171(.O (I22046), .I (g19330));
INVX1 gate6172(.O (g23942), .I (g21562));
INVX1 gate6173(.O (I20399), .I (g16205));
INVX1 gate6174(.O (g23341), .I (g21163));
INVX1 gate6175(.O (g18092), .I (I18882));
INVX1 gate6176(.O (g21268), .I (g15680));
INVX1 gate6177(.O (I14192), .I (g10233));
INVX1 gate6178(.O (I18048), .I (g13638));
INVX1 gate6179(.O (I28062), .I (g29194));
INVX1 gate6180(.O (g25226), .I (g22763));
INVX1 gate6181(.O (g22137), .I (g21370));
INVX1 gate6182(.O (g21156), .I (g17247));
INVX1 gate6183(.O (g17821), .I (I18829));
INVX1 gate6184(.O (g8178), .I (I12437));
INVX1 gate6185(.O (g6801), .I (g391));
INVX1 gate6186(.O (I21006), .I (g15579));
INVX1 gate6187(.O (g28615), .I (g27817));
INVX1 gate6188(.O (I16875), .I (g6675));
INVX1 gate6189(.O (g25481), .I (g22228));
INVX1 gate6190(.O (I15893), .I (g10430));
INVX1 gate6191(.O (I31878), .I (g33696));
INVX1 gate6192(.O (g19649), .I (g17015));
INVX1 gate6193(.O (I32874), .I (g34504));
INVX1 gate6194(.O (g21180), .I (g18008));
INVX1 gate6195(.O (I14663), .I (g9747));
INVX1 gate6196(.O (g21670), .I (g16540));
INVX1 gate6197(.O (I18221), .I (g13605));
INVX1 gate6198(.O (g16722), .I (I17938));
INVX1 gate6199(.O (g16924), .I (I18092));
INVX1 gate6200(.O (g20555), .I (g15480));
INVX1 gate6201(.O (g32817), .I (g31376));
INVX1 gate6202(.O (I28851), .I (g29317));
INVX1 gate6203(.O (I28872), .I (g30072));
INVX1 gate6204(.O (I32693), .I (g34433));
INVX1 gate6205(.O (g8135), .I (I12418));
INVX1 gate6206(.O (I21222), .I (g18091));
INVX1 gate6207(.O (g19491), .I (g16349));
INVX1 gate6208(.O (g34181), .I (g33913));
INVX1 gate6209(.O (g34671), .I (I32797));
INVX1 gate6210(.O (g20570), .I (g15277));
INVX1 gate6211(.O (g20712), .I (g15509));
INVX1 gate6212(.O (g11865), .I (g10124));
INVX1 gate6213(.O (I22302), .I (g19353));
INVX1 gate6214(.O (g13865), .I (I16168));
INVX1 gate6215(.O (g20914), .I (g15373));
INVX1 gate6216(.O (g21335), .I (I21067));
INVX1 gate6217(.O (g18883), .I (g15938));
INVX1 gate6218(.O (g32532), .I (g31170));
INVX1 gate6219(.O (g32901), .I (g31327));
INVX1 gate6220(.O (g14639), .I (I16747));
INVX1 gate6221(.O (g10230), .I (I13694));
INVX1 gate6222(.O (g23335), .I (g20391));
INVX1 gate6223(.O (I32665), .I (g34386));
INVX1 gate6224(.O (g19755), .I (g15915));
INVX1 gate6225(.O (g6755), .I (I11620));
INVX1 gate6226(.O (g12921), .I (g12228));
INVX1 gate6227(.O (g23839), .I (g18997));
INVX1 gate6228(.O (I17787), .I (g3267));
INVX1 gate6229(.O (g17873), .I (I18849));
INVX1 gate6230(.O (g23930), .I (g19147));
INVX1 gate6231(.O (g23993), .I (g19277));
INVX1 gate6232(.O (g32783), .I (g30825));
INVX1 gate6233(.O (g19770), .I (g17062));
INVX1 gate6234(.O (I29199), .I (g30237));
INVX1 gate6235(.O (g30931), .I (I28913));
INVX1 gate6236(.O (g8805), .I (I12799));
INVX1 gate6237(.O (I14862), .I (g8092));
INVX1 gate6238(.O (g8916), .I (I12887));
INVX1 gate6239(.O (I16160), .I (g11237));
INVX1 gate6240(.O (g21694), .I (g16540));
INVX1 gate6241(.O (g23838), .I (g18997));
INVX1 gate6242(.O (g9861), .I (g5459));
INVX1 gate6243(.O (g10416), .I (g10318));
INVX1 gate6244(.O (I15705), .I (g12218));
INVX1 gate6245(.O (g9048), .I (I12963));
INVX1 gate6246(.O (I17302), .I (g14044));
INVX1 gate6247(.O (g32561), .I (g30614));
INVX1 gate6248(.O (g32656), .I (g30673));
INVX1 gate6249(.O (g23965), .I (g21611));
INVX1 gate6250(.O (I31459), .I (g33219));
INVX1 gate6251(.O (g20239), .I (g17128));
INVX1 gate6252(.O (I32476), .I (g34277));
INVX1 gate6253(.O (g11705), .I (I14576));
INVX1 gate6254(.O (I22640), .I (g21256));
INVX1 gate6255(.O (g24074), .I (g21193));
INVX1 gate6256(.O (I22769), .I (g21277));
INVX1 gate6257(.O (g26860), .I (I25594));
INVX1 gate6258(.O (I14326), .I (g8607));
INVX1 gate6259(.O (g34426), .I (I32449));
INVX1 gate6260(.O (g11042), .I (g8691));
INVX1 gate6261(.O (g16031), .I (I17436));
INVX1 gate6262(.O (g20567), .I (g15426));
INVX1 gate6263(.O (g20594), .I (g15277));
INVX1 gate6264(.O (g32680), .I (g31376));
INVX1 gate6265(.O (g10391), .I (g6988));
INVX1 gate6266(.O (I16455), .I (g11845));
INVX1 gate6267(.O (g32823), .I (g31327));
INVX1 gate6268(.O (g20238), .I (g17096));
INVX1 gate6269(.O (g25297), .I (g23746));
INVX1 gate6270(.O (g13255), .I (g10632));
INVX1 gate6271(.O (g9827), .I (g1974));
INVX1 gate6272(.O (g13189), .I (g10762));
INVX1 gate6273(.O (g22542), .I (g19801));
INVX1 gate6274(.O (g13679), .I (g10573));
INVX1 gate6275(.O (g28142), .I (I26649));
INVX1 gate6276(.O (g31811), .I (g29385));
INVX1 gate6277(.O (g23487), .I (g20924));
INVX1 gate6278(.O (g14510), .I (I16629));
INVX1 gate6279(.O (g31646), .I (I29228));
INVX1 gate6280(.O (g9333), .I (g417));
INVX1 gate6281(.O (I14702), .I (g7717));
INVX1 gate6282(.O (g19794), .I (g16489));
INVX1 gate6283(.O (g11678), .I (I14563));
INVX1 gate6284(.O (g12184), .I (I15036));
INVX1 gate6285(.O (g16529), .I (g14055));
INVX1 gate6286(.O (g29081), .I (g27837));
INVX1 gate6287(.O (g12805), .I (g9511));
INVX1 gate6288(.O (g13188), .I (g10909));
INVX1 gate6289(.O (g19395), .I (g16431));
INVX1 gate6290(.O (g23502), .I (g21070));
INVX1 gate6291(.O (I27927), .I (g28803));
INVX1 gate6292(.O (g20382), .I (g15171));
INVX1 gate6293(.O (I16201), .I (g4023));
INVX1 gate6294(.O (I23351), .I (g23263));
INVX1 gate6295(.O (I31545), .I (g33219));
INVX1 gate6296(.O (I23372), .I (g23361));
INVX1 gate6297(.O (g26700), .I (g25429));
INVX1 gate6298(.O (g7258), .I (g4414));
INVX1 gate6299(.O (I33079), .I (g34809));
INVX1 gate6300(.O (g11686), .I (I14567));
INVX1 gate6301(.O (g16528), .I (g14154));
INVX1 gate6302(.O (g7577), .I (g1263));
INVX1 gate6303(.O (g7867), .I (g1489));
INVX1 gate6304(.O (g13460), .I (I15942));
INVX1 gate6305(.O (g15831), .I (g13385));
INVX1 gate6306(.O (I26479), .I (g25771));
INVX1 gate6307(.O (I12927), .I (g4332));
INVX1 gate6308(.O (g26987), .I (g26131));
INVX1 gate6309(.O (g11383), .I (g9061));
INVX1 gate6310(.O (g10014), .I (g6439));
INVX1 gate6311(.O (g23443), .I (g21468));
INVX1 gate6312(.O (I15030), .I (g10073));
INVX1 gate6313(.O (I18795), .I (g5327));
INVX1 gate6314(.O (g21279), .I (g15680));
INVX1 gate6315(.O (g24176), .I (I23372));
INVX1 gate6316(.O (g24185), .I (I23399));
INVX1 gate6317(.O (g23279), .I (g21037));
INVX1 gate6318(.O (g32966), .I (g31021));
INVX1 gate6319(.O (g19633), .I (g16931));
INVX1 gate6320(.O (g7717), .I (I12172));
INVX1 gate6321(.O (g30088), .I (g29094));
INVX1 gate6322(.O (g24092), .I (g20857));
INVX1 gate6323(.O (I32074), .I (g33670));
INVX1 gate6324(.O (g29945), .I (I28174));
INVX1 gate6325(.O (g6868), .I (I11688));
INVX1 gate6326(.O (g11030), .I (g8292));
INVX1 gate6327(.O (g20154), .I (I20412));
INVX1 gate6328(.O (g22905), .I (I22114));
INVX1 gate6329(.O (g32631), .I (g30825));
INVX1 gate6330(.O (g19719), .I (g16897));
INVX1 gate6331(.O (g21278), .I (I21013));
INVX1 gate6332(.O (g11294), .I (g7598));
INVX1 gate6333(.O (g24154), .I (I23306));
INVX1 gate6334(.O (I32594), .I (g34298));
INVX1 gate6335(.O (g8037), .I (g405));
INVX1 gate6336(.O (g23278), .I (g20283));
INVX1 gate6337(.O (g13267), .I (I15831));
INVX1 gate6338(.O (g29999), .I (g28973));
INVX1 gate6339(.O (g32364), .I (I29894));
INVX1 gate6340(.O (g6767), .I (I11626));
INVX1 gate6341(.O (g17614), .I (I18571));
INVX1 gate6342(.O (g22593), .I (g19801));
INVX1 gate6343(.O (g9780), .I (I13360));
INVX1 gate6344(.O (g16960), .I (I18114));
INVX1 gate6345(.O (g20637), .I (g15224));
INVX1 gate6346(.O (g26943), .I (I25695));
INVX1 gate6347(.O (g8102), .I (g3072));
INVX1 gate6348(.O (g13065), .I (g10476));
INVX1 gate6349(.O (g19718), .I (g17015));
INVX1 gate6350(.O (g21286), .I (g15509));
INVX1 gate6351(.O (g8302), .I (g1926));
INVX1 gate6352(.O (g14442), .I (I16593));
INVX1 gate6353(.O (g29998), .I (g28966));
INVX1 gate6354(.O (g17607), .I (I18560));
INVX1 gate6355(.O (g21468), .I (I21181));
INVX1 gate6356(.O (g17320), .I (I18297));
INVX1 gate6357(.O (g21306), .I (g15582));
INVX1 gate6358(.O (g31850), .I (g29385));
INVX1 gate6359(.O (g8579), .I (g2771));
INVX1 gate6360(.O (g23306), .I (g20924));
INVX1 gate6361(.O (I29225), .I (g30311));
INVX1 gate6362(.O (I31817), .I (g33323));
INVX1 gate6363(.O (g7975), .I (g3040));
INVX1 gate6364(.O (g33850), .I (I31701));
INVX1 gate6365(.O (g17530), .I (g14947));
INVX1 gate6366(.O (g10116), .I (g2413));
INVX1 gate6367(.O (g9662), .I (g3983));
INVX1 gate6368(.O (g9018), .I (g4273));
INVX1 gate6369(.O (g11875), .I (I14687));
INVX1 gate6370(.O (g8719), .I (I12719));
INVX1 gate6371(.O (g27013), .I (I25743));
INVX1 gate6372(.O (g7026), .I (g5507));
INVX1 gate6373(.O (I32675), .I (g34427));
INVX1 gate6374(.O (g9467), .I (g6434));
INVX1 gate6375(.O (g19440), .I (g15915));
INVX1 gate6376(.O (g16709), .I (I17919));
INVX1 gate6377(.O (g17122), .I (g14348));
INVX1 gate6378(.O (g34126), .I (I32067));
INVX1 gate6379(.O (g34659), .I (I32775));
INVX1 gate6380(.O (I12770), .I (g4200));
INVX1 gate6381(.O (I12563), .I (g3798));
INVX1 gate6382(.O (g12013), .I (I14866));
INVX1 gate6383(.O (g23815), .I (g19074));
INVX1 gate6384(.O (g34987), .I (I33261));
INVX1 gate6385(.O (I25677), .I (g25640));
INVX1 gate6386(.O (I15837), .I (g1459));
INVX1 gate6387(.O (I33158), .I (g34897));
INVX1 gate6388(.O (g7170), .I (g5719));
INVX1 gate6389(.O (g19861), .I (g17096));
INVX1 gate6390(.O (g10275), .I (g4584));
INVX1 gate6391(.O (g19573), .I (g16877));
INVX1 gate6392(.O (g8917), .I (I12890));
INVX1 gate6393(.O (g16708), .I (I17916));
INVX1 gate6394(.O (g22153), .I (g18997));
INVX1 gate6395(.O (g21677), .I (I21238));
INVX1 gate6396(.O (g33228), .I (I30766));
INVX1 gate6397(.O (g10430), .I (I13847));
INVX1 gate6398(.O (g14275), .I (g12358));
INVX1 gate6399(.O (g25546), .I (g22550));
INVX1 gate6400(.O (g32571), .I (g31376));
INVX1 gate6401(.O (I31561), .I (g33197));
INVX1 gate6402(.O (I17249), .I (g13605));
INVX1 gate6403(.O (g25211), .I (g22763));
INVX1 gate6404(.O (I32935), .I (g34657));
INVX1 gate6405(.O (g22409), .I (I21860));
INVX1 gate6406(.O (g19389), .I (g17532));
INVX1 gate6407(.O (g17641), .I (g14845));
INVX1 gate6408(.O (g20501), .I (g17955));
INVX1 gate6409(.O (g26870), .I (I25606));
INVX1 gate6410(.O (g30296), .I (g28889));
INVX1 gate6411(.O (g20577), .I (g15483));
INVX1 gate6412(.O (g34339), .I (g34077));
INVX1 gate6413(.O (g9816), .I (g6167));
INVX1 gate6414(.O (g34943), .I (I33197));
INVX1 gate6415(.O (I20951), .I (g17782));
INVX1 gate6416(.O (g25024), .I (g22472));
INVX1 gate6417(.O (g33716), .I (I31569));
INVX1 gate6418(.O (I31823), .I (g33149));
INVX1 gate6419(.O (g19612), .I (g16897));
INVX1 gate6420(.O (g34296), .I (I32297));
INVX1 gate6421(.O (g7280), .I (g2153));
INVX1 gate6422(.O (g29897), .I (I28128));
INVX1 gate6423(.O (g7939), .I (g1280));
INVX1 gate6424(.O (g22136), .I (g20277));
INVX1 gate6425(.O (g29961), .I (g28892));
INVX1 gate6426(.O (g8442), .I (g3476));
INVX1 gate6427(.O (g22408), .I (g19483));
INVX1 gate6428(.O (g22635), .I (g19801));
INVX1 gate6429(.O (I12767), .I (g4197));
INVX1 gate6430(.O (g14237), .I (g11666));
INVX1 gate6431(.O (g8786), .I (I12770));
INVX1 gate6432(.O (g23937), .I (g19277));
INVX1 gate6433(.O (g10035), .I (g1720));
INVX1 gate6434(.O (g32495), .I (g31070));
INVX1 gate6435(.O (g29505), .I (g29186));
INVX1 gate6436(.O (g19777), .I (g17015));
INVX1 gate6437(.O (g17409), .I (I18344));
INVX1 gate6438(.O (I12899), .I (g4232));
INVX1 gate6439(.O (g7544), .I (g918));
INVX1 gate6440(.O (g8164), .I (g3484));
INVX1 gate6441(.O (g9381), .I (g5527));
INVX1 gate6442(.O (I15617), .I (g12037));
INVX1 gate6443(.O (I13805), .I (g6976));
INVX1 gate6444(.O (I18788), .I (g13138));
INVX1 gate6445(.O (g8364), .I (g1585));
INVX1 gate6446(.O (g32816), .I (g31327));
INVX1 gate6447(.O (I15915), .I (g10430));
INVX1 gate6448(.O (g24438), .I (g22722));
INVX1 gate6449(.O (g11470), .I (g7625));
INVX1 gate6450(.O (g17136), .I (g14348));
INVX1 gate6451(.O (g10142), .I (I13637));
INVX1 gate6452(.O (g17408), .I (I18341));
INVX1 gate6453(.O (g34060), .I (g33704));
INVX1 gate6454(.O (g29212), .I (I27552));
INVX1 gate6455(.O (g7636), .I (g4098));
INVX1 gate6456(.O (g9685), .I (g6533));
INVX1 gate6457(.O (I26676), .I (g27736));
INVX1 gate6458(.O (g9197), .I (g1221));
INVX1 gate6459(.O (I18829), .I (g13350));
INVX1 gate6460(.O (g32687), .I (g31376));
INVX1 gate6461(.O (g9397), .I (g6088));
INVX1 gate6462(.O (I18434), .I (g13782));
INVX1 gate6463(.O (g33959), .I (I31878));
INVX1 gate6464(.O (g9021), .I (I12954));
INVX1 gate6465(.O (I12719), .I (g365));
INVX1 gate6466(.O (g16602), .I (g14101));
INVX1 gate6467(.O (g21410), .I (g15224));
INVX1 gate6468(.O (g34197), .I (g33812));
INVX1 gate6469(.O (I27718), .I (g28231));
INVX1 gate6470(.O (I16401), .I (g869));
INVX1 gate6471(.O (g16774), .I (g14024));
INVX1 gate6472(.O (g23410), .I (g21562));
INVX1 gate6473(.O (g8770), .I (g749));
INVX1 gate6474(.O (I29337), .I (g30286));
INVX1 gate6475(.O (g34855), .I (I33079));
INVX1 gate6476(.O (I26654), .I (g27576));
INVX1 gate6477(.O (I22380), .I (g21156));
INVX1 gate6478(.O (g16955), .I (I18107));
INVX1 gate6479(.O (g32752), .I (g31376));
INVX1 gate6480(.O (g8296), .I (g246));
INVX1 gate6481(.O (g25250), .I (I24434));
INVX1 gate6482(.O (g27100), .I (g26759));
INVX1 gate6483(.O (g32954), .I (g31376));
INVX1 gate6484(.O (g8725), .I (g739));
INVX1 gate6485(.O (g24083), .I (g19984));
INVX1 gate6486(.O (g33378), .I (I30904));
INVX1 gate6487(.O (g21666), .I (g16540));
INVX1 gate6488(.O (g23479), .I (g21562));
INVX1 gate6489(.O (I26936), .I (g27599));
INVX1 gate6490(.O (g32643), .I (g31376));
INVX1 gate6491(.O (g6940), .I (g4035));
INVX1 gate6492(.O (I15494), .I (g10385));
INVX1 gate6493(.O (g13075), .I (I15705));
INVX1 gate6494(.O (g23363), .I (I22470));
INVX1 gate6495(.O (I18344), .I (g13003));
INVX1 gate6496(.O (g7187), .I (g6065));
INVX1 gate6497(.O (g7387), .I (g2421));
INVX1 gate6498(.O (g20622), .I (g15595));
INVX1 gate6499(.O (g11467), .I (g7623));
INVX1 gate6500(.O (g13595), .I (g10951));
INVX1 gate6501(.O (I17999), .I (g4012));
INVX1 gate6502(.O (g20566), .I (g15224));
INVX1 gate6503(.O (g7461), .I (g2567));
INVX1 gate6504(.O (I15623), .I (g12040));
INVX1 gate6505(.O (g23478), .I (g21514));
INVX1 gate6506(.O (g13494), .I (g11912));
INVX1 gate6507(.O (g23015), .I (g20391));
INVX1 gate6508(.O (g8553), .I (g3747));
INVX1 gate6509(.O (I26334), .I (g26834));
INVX1 gate6510(.O (I19707), .I (g17590));
INVX1 gate6511(.O (g25296), .I (g23745));
INVX1 gate6512(.O (g10130), .I (g5694));
INVX1 gate6513(.O (g16171), .I (g13530));
INVX1 gate6514(.O (g33944), .I (I31829));
INVX1 gate6515(.O (g19061), .I (I19762));
INVX1 gate6516(.O (g26818), .I (I25530));
INVX1 gate6517(.O (g16886), .I (I18078));
INVX1 gate6518(.O (I27573), .I (g28157));
INVX1 gate6519(.O (g32669), .I (g30614));
INVX1 gate6520(.O (I15782), .I (g10430));
INVX1 gate6521(.O (g23486), .I (g20785));
INVX1 gate6522(.O (g26055), .I (I25115));
INVX1 gate6523(.O (g13037), .I (g10981));
INVX1 gate6524(.O (g10362), .I (g6850));
INVX1 gate6525(.O (g29149), .I (g27837));
INVX1 gate6526(.O (g7027), .I (g5499));
INVX1 gate6527(.O (I19818), .I (g1056));
INVX1 gate6528(.O (g19766), .I (g16449));
INVX1 gate6529(.O (g21556), .I (g15669));
INVX1 gate6530(.O (I12861), .I (g4372));
INVX1 gate6531(.O (g10165), .I (g5698));
INVX1 gate6532(.O (g13782), .I (I16117));
INVX1 gate6533(.O (g17575), .I (g14921));
INVX1 gate6534(.O (g28137), .I (I26638));
INVX1 gate6535(.O (g11984), .I (g9186));
INVX1 gate6536(.O (g16967), .I (I18125));
INVX1 gate6537(.O (I22331), .I (g19417));
INVX1 gate6538(.O (g32668), .I (g31070));
INVX1 gate6539(.O (g32842), .I (g31710));
INVX1 gate6540(.O (g17711), .I (I18694));
INVX1 gate6541(.O (g7046), .I (g5791));
INVX1 gate6542(.O (I32284), .I (g34052));
INVX1 gate6543(.O (g20653), .I (I20747));
INVX1 gate6544(.O (g27991), .I (g25852));
INVX1 gate6545(.O (I33288), .I (g34989));
INVX1 gate6546(.O (g31802), .I (g29385));
INVX1 gate6547(.O (g9631), .I (g6573));
INVX1 gate6548(.O (g17327), .I (I18310));
INVX1 gate6549(.O (g25060), .I (g23708));
INVX1 gate6550(.O (g32489), .I (g30614));
INVX1 gate6551(.O (g8389), .I (g3125));
INVX1 gate6552(.O (I13329), .I (g86));
INVX1 gate6553(.O (I27388), .I (g27698));
INVX1 gate6554(.O (g31857), .I (g29385));
INVX1 gate6555(.O (g7446), .I (g1256));
INVX1 gate6556(.O (g18200), .I (I19012));
INVX1 gate6557(.O (g29811), .I (g28376));
INVX1 gate6558(.O (g23223), .I (g21308));
INVX1 gate6559(.O (g7514), .I (g6704));
INVX1 gate6560(.O (g19360), .I (g16249));
INVX1 gate6561(.O (g11418), .I (I14424));
INVX1 gate6562(.O (g34714), .I (I32874));
INVX1 gate6563(.O (g8990), .I (g146));
INVX1 gate6564(.O (g12882), .I (g10389));
INVX1 gate6565(.O (g9257), .I (g5115));
INVX1 gate6566(.O (g22492), .I (g19614));
INVX1 gate6567(.O (g25197), .I (g23958));
INVX1 gate6568(.O (g29343), .I (g28174));
INVX1 gate6569(.O (g7003), .I (g5152));
INVX1 gate6570(.O (I13539), .I (g6381));
INVX1 gate6571(.O (g22303), .I (g19277));
INVX1 gate6572(.O (I27777), .I (g29043));
INVX1 gate6573(.O (g9817), .I (I13374));
INVX1 gate6574(.O (g32559), .I (g30825));
INVX1 gate6575(.O (g34315), .I (g34085));
INVX1 gate6576(.O (g10475), .I (g8844));
INVX1 gate6577(.O (I17932), .I (g3310));
INVX1 gate6578(.O (g24138), .I (g21143));
INVX1 gate6579(.O (g32525), .I (g31170));
INVX1 gate6580(.O (g32488), .I (g31194));
INVX1 gate6581(.O (g11170), .I (g8476));
INVX1 gate6582(.O (g34910), .I (g34864));
INVX1 gate6583(.O (I29444), .I (g30928));
INVX1 gate6584(.O (g8171), .I (g3817));
INVX1 gate6585(.O (g10727), .I (I14016));
INVX1 gate6586(.O (g7345), .I (g6415));
INVX1 gate6587(.O (g7841), .I (g904));
INVX1 gate6588(.O (I12534), .I (g50));
INVX1 gate6589(.O (g20636), .I (g18008));
INVX1 gate6590(.O (I19384), .I (g15085));
INVX1 gate6591(.O (g8787), .I (I12773));
INVX1 gate6592(.O (g32558), .I (g30735));
INVX1 gate6593(.O (g34202), .I (I32161));
INVX1 gate6594(.O (g23084), .I (g19954));
INVX1 gate6595(.O (g24636), .I (g23121));
INVX1 gate6596(.O (g6826), .I (g218));
INVX1 gate6597(.O (g10222), .I (g4492));
INVX1 gate6598(.O (g7191), .I (g6398));
INVX1 gate6599(.O (g30055), .I (g29157));
INVX1 gate6600(.O (g17606), .I (g14999));
INVX1 gate6601(.O (g20852), .I (g15595));
INVX1 gate6602(.O (g32830), .I (g31327));
INVX1 gate6603(.O (g23922), .I (g18997));
INVX1 gate6604(.O (g23321), .I (I22422));
INVX1 gate6605(.O (g32893), .I (g30937));
INVX1 gate6606(.O (I18028), .I (g13638));
INVX1 gate6607(.O (g21179), .I (g15373));
INVX1 gate6608(.O (I24920), .I (g25513));
INVX1 gate6609(.O (g26801), .I (I25511));
INVX1 gate6610(.O (I24434), .I (g22763));
INVX1 gate6611(.O (g29368), .I (I27730));
INVX1 gate6612(.O (g9751), .I (g1710));
INVX1 gate6613(.O (g34070), .I (g33725));
INVX1 gate6614(.O (g8281), .I (g3494));
INVX1 gate6615(.O (g32544), .I (g30735));
INVX1 gate6616(.O (g19629), .I (g17015));
INVX1 gate6617(.O (g32865), .I (g31327));
INVX1 gate6618(.O (g19451), .I (g15938));
INVX1 gate6619(.O (g21178), .I (g17955));
INVX1 gate6620(.O (g34590), .I (I32678));
INVX1 gate6621(.O (g19472), .I (g16349));
INVX1 gate6622(.O (g24963), .I (g22342));
INVX1 gate6623(.O (g20664), .I (g15373));
INVX1 gate6624(.O (g34986), .I (I33258));
INVX1 gate6625(.O (g32713), .I (g30673));
INVX1 gate6626(.O (g7536), .I (g5976));
INVX1 gate6627(.O (g9585), .I (g1616));
INVX1 gate6628(.O (g8297), .I (g142));
INVX1 gate6629(.O (g10347), .I (I13759));
INVX1 gate6630(.O (g21685), .I (I21246));
INVX1 gate6631(.O (I16733), .I (g12026));
INVX1 gate6632(.O (I12997), .I (g351));
INVX1 gate6633(.O (g28726), .I (g27937));
INVX1 gate6634(.O (g34384), .I (I32391));
INVX1 gate6635(.O (g23953), .I (g19277));
INVX1 gate6636(.O (g30067), .I (g29060));
INVX1 gate6637(.O (g11401), .I (g7593));
INVX1 gate6638(.O (g22840), .I (g20330));
INVX1 gate6639(.O (g21654), .I (g17619));
INVX1 gate6640(.O (I29977), .I (g31596));
INVX1 gate6641(.O (g7858), .I (g947));
INVX1 gate6642(.O (g32610), .I (g31070));
INVX1 gate6643(.O (g20576), .I (g18065));
INVX1 gate6644(.O (g20585), .I (g17955));
INVX1 gate6645(.O (g23654), .I (g20248));
INVX1 gate6646(.O (I12061), .I (g562));
INVX1 gate6647(.O (g32705), .I (g30614));
INVX1 gate6648(.O (g34094), .I (g33772));
INVX1 gate6649(.O (g13477), .I (I15954));
INVX1 gate6650(.O (g8745), .I (g744));
INVX1 gate6651(.O (g28436), .I (I26929));
INVX1 gate6652(.O (g8138), .I (g1500));
INVX1 gate6653(.O (g8639), .I (g2807));
INVX1 gate6654(.O (g24585), .I (g23063));
INVX1 gate6655(.O (I22149), .I (g21036));
INVX1 gate6656(.O (g19071), .I (g15591));
INVX1 gate6657(.O (g23800), .I (g21246));
INVX1 gate6658(.O (I23711), .I (g23192));
INVX1 gate6659(.O (g20554), .I (g15348));
INVX1 gate6660(.O (g23417), .I (g20391));
INVX1 gate6661(.O (g32679), .I (g31579));
INVX1 gate6662(.O (g16322), .I (I17650));
INVX1 gate6663(.O (g8791), .I (I12787));
INVX1 gate6664(.O (g10351), .I (g6802));
INVX1 gate6665(.O (g23936), .I (g19210));
INVX1 gate6666(.O (g10372), .I (g6900));
INVX1 gate6667(.O (I23327), .I (g22647));
INVX1 gate6668(.O (g25202), .I (g23932));
INVX1 gate6669(.O (g19776), .I (g17015));
INVX1 gate6670(.O (g19785), .I (g16987));
INVX1 gate6671(.O (g34150), .I (I32103));
INVX1 gate6672(.O (I32963), .I (g34650));
INVX1 gate6673(.O (g16159), .I (g13584));
INVX1 gate6674(.O (g22192), .I (g19801));
INVX1 gate6675(.O (g20609), .I (g15373));
INVX1 gate6676(.O (g28274), .I (I26799));
INVX1 gate6677(.O (g15171), .I (I17098));
INVX1 gate6678(.O (g34877), .I (I33103));
INVX1 gate6679(.O (g10175), .I (g28));
INVX1 gate6680(.O (I17723), .I (g13177));
INVX1 gate6681(.O (g12082), .I (g9645));
INVX1 gate6682(.O (g17390), .I (g14755));
INVX1 gate6683(.O (g28593), .I (g27727));
INVX1 gate6684(.O (g32678), .I (g31528));
INVX1 gate6685(.O (g13022), .I (g11894));
INVX1 gate6686(.O (g7522), .I (g6661));
INVX1 gate6687(.O (g23334), .I (g20785));
INVX1 gate6688(.O (g25055), .I (g23590));
INVX1 gate6689(.O (g19147), .I (I19786));
INVX1 gate6690(.O (g30019), .I (g29060));
INVX1 gate6691(.O (g7115), .I (g12));
INVX1 gate6692(.O (g12107), .I (g9687));
INVX1 gate6693(.O (g8808), .I (g595));
INVX1 gate6694(.O (g19754), .I (g17062));
INVX1 gate6695(.O (g7315), .I (g1772));
INVX1 gate6696(.O (g16158), .I (g13555));
INVX1 gate6697(.O (g20608), .I (g15171));
INVX1 gate6698(.O (g25111), .I (g23699));
INVX1 gate6699(.O (g9669), .I (g5092));
INVX1 gate6700(.O (g19355), .I (g16027));
INVX1 gate6701(.O (I12360), .I (g528));
INVX1 gate6702(.O (g25070), .I (g23590));
INVX1 gate6703(.O (g32460), .I (g31194));
INVX1 gate6704(.O (g32686), .I (g31579));
INVX1 gate6705(.O (I22343), .I (g19371));
INVX1 gate6706(.O (g24115), .I (g20998));
INVX1 gate6707(.O (g32939), .I (g31327));
INVX1 gate6708(.O (I18903), .I (g16872));
INVX1 gate6709(.O (g30018), .I (g28987));
INVX1 gate6710(.O (g32383), .I (I29913));
INVX1 gate6711(.O (g19950), .I (g15885));
INVX1 gate6712(.O (g14063), .I (g11048));
INVX1 gate6713(.O (g19370), .I (g15915));
INVX1 gate6714(.O (I19917), .I (g18088));
INVX1 gate6715(.O (I14046), .I (g9900));
INVX1 gate6716(.O (I17148), .I (g14442));
INVX1 gate6717(.O (g16656), .I (I17852));
INVX1 gate6718(.O (g9772), .I (I13352));
INVX1 gate6719(.O (I26638), .I (g27965));
INVX1 gate6720(.O (g20921), .I (g15426));
INVX1 gate6721(.O (g12345), .I (g7158));
INVX1 gate6722(.O (I16476), .I (g10430));
INVX1 gate6723(.O (g14790), .I (I16855));
INVX1 gate6724(.O (g20052), .I (g17533));
INVX1 gate6725(.O (g23964), .I (g19147));
INVX1 gate6726(.O (I23303), .I (g21669));
INVX1 gate6727(.O (g32938), .I (g30937));
INVX1 gate6728(.O (g28034), .I (g26365));
INVX1 gate6729(.O (g33533), .I (I31361));
INVX1 gate6730(.O (g29310), .I (g28991));
INVX1 gate6731(.O (g16680), .I (g13223));
INVX1 gate6732(.O (g24052), .I (g21193));
INVX1 gate6733(.O (I17104), .I (g12932));
INVX1 gate6734(.O (g12940), .I (g11744));
INVX1 gate6735(.O (g17522), .I (g14927));
INVX1 gate6736(.O (g21423), .I (g15224));
INVX1 gate6737(.O (g12399), .I (g9920));
INVX1 gate6738(.O (g9743), .I (I13321));
INVX1 gate6739(.O (I16555), .I (g10430));
INVX1 gate6740(.O (g23423), .I (g20871));
INVX1 gate6741(.O (g8201), .I (g1894));
INVX1 gate6742(.O (g9890), .I (g6058));
INVX1 gate6743(.O (g13305), .I (g11048));
INVX1 gate6744(.O (g6827), .I (g1277));
INVX1 gate6745(.O (g14873), .I (I16898));
INVX1 gate6746(.O (g23216), .I (g20924));
INVX1 gate6747(.O (g11900), .I (I14708));
INVX1 gate6748(.O (g19996), .I (g17271));
INVX1 gate6749(.O (g29379), .I (I27749));
INVX1 gate6750(.O (g29925), .I (g28820));
INVX1 gate6751(.O (g13809), .I (I16135));
INVX1 gate6752(.O (I23381), .I (g23322));
INVX1 gate6753(.O (I15036), .I (g799));
INVX1 gate6754(.O (g8449), .I (g3752));
INVX1 gate6755(.O (g12804), .I (g9927));
INVX1 gate6756(.O (g9011), .I (g1422));
INVX1 gate6757(.O (g19367), .I (I19851));
INVX1 gate6758(.O (g19394), .I (g16326));
INVX1 gate6759(.O (I12451), .I (g3092));
INVX1 gate6760(.O (g6846), .I (g2152));
INVX1 gate6761(.O (g9856), .I (g5343));
INVX1 gate6762(.O (g8575), .I (g291));
INVX1 gate6763(.O (g13036), .I (g10981));
INVX1 gate6764(.O (g32875), .I (g31376));
INVX1 gate6765(.O (g30917), .I (I28897));
INVX1 gate6766(.O (I14827), .I (g9686));
INVX1 gate6767(.O (g11560), .I (g7647));
INVX1 gate6768(.O (g13101), .I (I15736));
INVX1 gate6769(.O (g14209), .I (g11415));
INVX1 gate6770(.O (g7880), .I (g1291));
INVX1 gate6771(.O (g13177), .I (I15782));
INVX1 gate6772(.O (g34917), .I (I33143));
INVX1 gate6773(.O (g8715), .I (g4927));
INVX1 gate6774(.O (g20674), .I (g15277));
INVX1 gate6775(.O (g7595), .I (I12067));
INVX1 gate6776(.O (g23543), .I (g21514));
INVX1 gate6777(.O (g6803), .I (g496));
INVX1 gate6778(.O (g16966), .I (g14291));
INVX1 gate6779(.O (g7537), .I (g311));
INVX1 gate6780(.O (g24184), .I (I23396));
INVX1 gate6781(.O (I18845), .I (g6711));
INVX1 gate6782(.O (I32921), .I (g34650));
INVX1 gate6783(.O (g16631), .I (g14454));
INVX1 gate6784(.O (g14208), .I (g11563));
INVX1 gate6785(.O (I18262), .I (g13857));
INVX1 gate6786(.O (g29944), .I (g28911));
INVX1 gate6787(.O (g22904), .I (I22111));
INVX1 gate6788(.O (g23000), .I (g20453));
INVX1 gate6789(.O (I26578), .I (g26941));
INVX1 gate6790(.O (g23908), .I (g20739));
INVX1 gate6791(.O (g17326), .I (I18307));
INVX1 gate6792(.O (g32837), .I (g31327));
INVX1 gate6793(.O (g31856), .I (g29385));
INVX1 gate6794(.O (I13206), .I (g5448));
INVX1 gate6795(.O (g8833), .I (g794));
INVX1 gate6796(.O (g30077), .I (g29057));
INVX1 gate6797(.O (g9992), .I (g5990));
INVX1 gate6798(.O (g20732), .I (g15595));
INVX1 gate6799(.O (g23569), .I (g21611));
INVX1 gate6800(.O (g25196), .I (g22763));
INVX1 gate6801(.O (g10542), .I (g7196));
INVX1 gate6802(.O (I31610), .I (g33149));
INVX1 gate6803(.O (I23390), .I (g23395));
INVX1 gate6804(.O (g13064), .I (g11705));
INVX1 gate6805(.O (g24732), .I (g23042));
INVX1 gate6806(.O (g14453), .I (I16610));
INVX1 gate6807(.O (g7017), .I (g128));
INVX1 gate6808(.O (I30992), .I (g32445));
INVX1 gate6809(.O (g7243), .I (I11892));
INVX1 gate6810(.O (g19446), .I (I19917));
INVX1 gate6811(.O (g34597), .I (I32699));
INVX1 gate6812(.O (I12776), .I (g4207));
INVX1 gate6813(.O (I13759), .I (g6754));
INVX1 gate6814(.O (I18191), .I (g14385));
INVX1 gate6815(.O (g23568), .I (g21611));
INVX1 gate6816(.O (I33255), .I (g34975));
INVX1 gate6817(.O (I33189), .I (g34929));
INVX1 gate6818(.O (g8584), .I (g3639));
INVX1 gate6819(.O (g8539), .I (g3454));
INVX1 gate6820(.O (g23242), .I (g21070));
INVX1 gate6821(.O (I32973), .I (g34714));
INVX1 gate6822(.O (I29571), .I (g31783));
INVX1 gate6823(.O (g34689), .I (I32837));
INVX1 gate6824(.O (I33270), .I (g34982));
INVX1 gate6825(.O (g34923), .I (I33161));
INVX1 gate6826(.O (g9863), .I (g5503));
INVX1 gate6827(.O (I12355), .I (g46));
INVX1 gate6828(.O (g16289), .I (g13223));
INVX1 gate6829(.O (g9480), .I (g559));
INVX1 gate6830(.O (I17228), .I (g13350));
INVX1 gate6831(.O (g6994), .I (g4933));
INVX1 gate6832(.O (g21123), .I (g15615));
INVX1 gate6833(.O (g18100), .I (I18906));
INVX1 gate6834(.O (g34688), .I (I32834));
INVX1 gate6835(.O (g9713), .I (g3618));
INVX1 gate6836(.O (g10607), .I (g10233));
INVX1 gate6837(.O (g12833), .I (I15448));
INVX1 gate6838(.O (g22847), .I (g20283));
INVX1 gate6839(.O (g16309), .I (I17639));
INVX1 gate6840(.O (I12950), .I (g4287));
INVX1 gate6841(.O (g23814), .I (g19074));
INVX1 gate6842(.O (g10320), .I (g817));
INVX1 gate6843(.O (g32617), .I (g30825));
INVX1 gate6844(.O (g28575), .I (g27711));
INVX1 gate6845(.O (g32470), .I (g31566));
INVX1 gate6846(.O (g10073), .I (g134));
INVX1 gate6847(.O (I18832), .I (g13782));
INVX1 gate6848(.O (I31686), .I (g33164));
INVX1 gate6849(.O (g7328), .I (g2197));
INVX1 gate6850(.O (g32915), .I (g31710));
INVX1 gate6851(.O (g10274), .I (g976));
INVX1 gate6852(.O (g29765), .I (I28014));
INVX1 gate6853(.O (g10530), .I (g8922));
INVX1 gate6854(.O (g7542), .I (I12030));
INVX1 gate6855(.O (I12858), .I (g4340));
INVX1 gate6856(.O (g28711), .I (g27886));
INVX1 gate6857(.O (g13009), .I (I15617));
INVX1 gate6858(.O (g16308), .I (I17636));
INVX1 gate6859(.O (g9569), .I (g6227));
INVX1 gate6860(.O (g13665), .I (g11306));
INVX1 gate6861(.O (g27004), .I (g26131));
INVX1 gate6862(.O (g30102), .I (g29157));
INVX1 gate6863(.O (g8362), .I (g194));
INVX1 gate6864(.O (I13744), .I (g3518));
INVX1 gate6865(.O (g31831), .I (g29385));
INVX1 gate6866(.O (g32201), .I (g31509));
INVX1 gate6867(.O (g24013), .I (g21611));
INVX1 gate6868(.O (I33030), .I (g34768));
INVX1 gate6869(.O (I12151), .I (g604));
INVX1 gate6870(.O (g10122), .I (I13623));
INVX1 gate6871(.O (g6816), .I (g933));
INVX1 gate6872(.O (I12172), .I (g2715));
INVX1 gate6873(.O (g17183), .I (I18221));
INVX1 gate6874(.O (g17673), .I (g14723));
INVX1 gate6875(.O (g17847), .I (I18839));
INVX1 gate6876(.O (I26430), .I (g26856));
INVX1 gate6877(.O (g13008), .I (g11855));
INVX1 gate6878(.O (g15656), .I (I17198));
INVX1 gate6879(.O (I21483), .I (g18726));
INVX1 gate6880(.O (g20329), .I (g15277));
INVX1 gate6881(.O (I33267), .I (g34979));
INVX1 gate6882(.O (g8052), .I (g1211));
INVX1 gate6883(.O (I18861), .I (g14307));
INVX1 gate6884(.O (g21293), .I (I21036));
INVX1 gate6885(.O (g20207), .I (g17015));
INVX1 gate6886(.O (g23230), .I (I22327));
INVX1 gate6887(.O (g15680), .I (I17207));
INVX1 gate6888(.O (g20539), .I (g15483));
INVX1 gate6889(.O (g25001), .I (g23666));
INVX1 gate6890(.O (g17062), .I (I18154));
INVX1 gate6891(.O (g20005), .I (g17433));
INVX1 gate6892(.O (g13485), .I (g10476));
INVX1 gate6893(.O (g20328), .I (g15867));
INVX1 gate6894(.O (g32595), .I (g30825));
INVX1 gate6895(.O (g32467), .I (g31194));
INVX1 gate6896(.O (g32494), .I (g30825));
INVX1 gate6897(.O (g19902), .I (g17200));
INVX1 gate6898(.O (g24005), .I (I23149));
INVX1 gate6899(.O (g17509), .I (I18446));
INVX1 gate6900(.O (g14034), .I (g11048));
INVX1 gate6901(.O (g19957), .I (g16540));
INVX1 gate6902(.O (g16816), .I (I18028));
INVX1 gate6903(.O (g20538), .I (g15348));
INVX1 gate6904(.O (g9688), .I (g113));
INVX1 gate6905(.O (g28606), .I (g27762));
INVX1 gate6906(.O (g6847), .I (g2283));
INVX1 gate6907(.O (g13555), .I (g12692));
INVX1 gate6908(.O (g18882), .I (I19674));
INVX1 gate6909(.O (g32623), .I (g30735));
INVX1 gate6910(.O (g18991), .I (g16136));
INVX1 gate6911(.O (I28897), .I (g30155));
INVX1 gate6912(.O (g19739), .I (g16931));
INVX1 gate6913(.O (I25391), .I (g24483));
INVX1 gate6914(.O (g9976), .I (g2537));
INVX1 gate6915(.O (g17508), .I (I18443));
INVX1 gate6916(.O (g29317), .I (I27677));
INVX1 gate6917(.O (g10153), .I (g2417));
INVX1 gate6918(.O (g23841), .I (g19074));
INVX1 gate6919(.O (I22096), .I (g19890));
INVX1 gate6920(.O (g23992), .I (g19210));
INVX1 gate6921(.O (g32782), .I (g30735));
INVX1 gate6922(.O (g23391), .I (g20645));
INVX1 gate6923(.O (g19146), .I (g15574));
INVX1 gate6924(.O (g19738), .I (g15992));
INVX1 gate6925(.O (g33080), .I (I30644));
INVX1 gate6926(.O (g21510), .I (g15647));
INVX1 gate6927(.O (g23510), .I (g18833));
INVX1 gate6928(.O (g10409), .I (g7087));
INVX1 gate6929(.O (g16752), .I (I17976));
INVX1 gate6930(.O (I21757), .I (g21308));
INVX1 gate6931(.O (I33218), .I (g34955));
INVX1 gate6932(.O (I25579), .I (g25297));
INVX1 gate6933(.O (g16954), .I (I18104));
INVX1 gate6934(.O (g29129), .I (g27858));
INVX1 gate6935(.O (g22213), .I (g19147));
INVX1 gate6936(.O (g19699), .I (I20116));
INVX1 gate6937(.O (g8504), .I (g3451));
INVX1 gate6938(.O (g34511), .I (g34419));
INVX1 gate6939(.O (g10136), .I (g6113));
INVX1 gate6940(.O (g16643), .I (I17839));
INVX1 gate6941(.O (g10408), .I (g7049));
INVX1 gate6942(.O (g9000), .I (g632));
INVX1 gate6943(.O (g32822), .I (g30937));
INVX1 gate6944(.O (g13074), .I (I15702));
INVX1 gate6945(.O (I24191), .I (g22360));
INVX1 gate6946(.O (g29128), .I (g27800));
INVX1 gate6947(.O (g14635), .I (I16741));
INVX1 gate6948(.O (I12227), .I (g34));
INVX1 gate6949(.O (g13239), .I (g10632));
INVX1 gate6950(.O (g19698), .I (g16971));
INVX1 gate6951(.O (g9326), .I (g6203));
INVX1 gate6952(.O (I15238), .I (g6351));
INVX1 gate6953(.O (g12951), .I (I15569));
INVX1 gate6954(.O (g25157), .I (g22498));
INVX1 gate6955(.O (g23578), .I (I22725));
INVX1 gate6956(.O (g8070), .I (g3518));
INVX1 gate6957(.O (g13594), .I (g11012));
INVX1 gate6958(.O (I16438), .I (g11165));
INVX1 gate6959(.O (g23014), .I (g20391));
INVX1 gate6960(.O (I25586), .I (g25537));
INVX1 gate6961(.O (g8470), .I (I12605));
INVX1 gate6962(.O (g20100), .I (I20369));
INVX1 gate6963(.O (g7512), .I (g5283));
INVX1 gate6964(.O (g34660), .I (g34473));
INVX1 gate6965(.O (I30983), .I (g32433));
INVX1 gate6966(.O (g9760), .I (g2315));
INVX1 gate6967(.O (g20771), .I (g15171));
INVX1 gate6968(.O (g22311), .I (g18935));
INVX1 gate6969(.O (g24100), .I (g20857));
INVX1 gate6970(.O (g26054), .I (g24804));
INVX1 gate6971(.O (g7490), .I (g2629));
INVX1 gate6972(.O (I15382), .I (g9071));
INVX1 gate6973(.O (I14647), .I (g7717));
INVX1 gate6974(.O (g25231), .I (g22228));
INVX1 gate6975(.O (g7166), .I (g4311));
INVX1 gate6976(.O (g20235), .I (g15277));
INVX1 gate6977(.O (g19427), .I (g16292));
INVX1 gate6978(.O (I26130), .I (g26510));
INVX1 gate6979(.O (g11941), .I (I14761));
INVX1 gate6980(.O (g19366), .I (g15885));
INVX1 gate6981(.O (I17857), .I (g3969));
INVX1 gate6982(.O (g32853), .I (g30673));
INVX1 gate6983(.O (g24683), .I (g23112));
INVX1 gate6984(.O (g33736), .I (I31597));
INVX1 gate6985(.O (g11519), .I (g8481));
INVX1 gate6986(.O (I14999), .I (g10030));
INVX1 gate6987(.O (g16195), .I (g13437));
INVX1 gate6988(.O (g34480), .I (I32535));
INVX1 gate6989(.O (g16489), .I (I17699));
INVX1 gate6990(.O (g34916), .I (I33140));
INVX1 gate6991(.O (g13675), .I (g10556));
INVX1 gate6992(.O (I20861), .I (g16960));
INVX1 gate6993(.O (g32589), .I (g31070));
INVX1 gate6994(.O (g7456), .I (g2495));
INVX1 gate6995(.O (g15224), .I (I17101));
INVX1 gate6996(.O (g7148), .I (I11835));
INVX1 gate6997(.O (g6817), .I (g956));
INVX1 gate6998(.O (g7649), .I (g1345));
INVX1 gate6999(.O (g22592), .I (I21930));
INVX1 gate7000(.O (g22756), .I (g20436));
INVX1 gate7001(.O (g16525), .I (I17723));
INVX1 gate7002(.O (g15571), .I (g13211));
INVX1 gate7003(.O (g26942), .I (I25692));
INVX1 gate7004(.O (g9924), .I (g5644));
INVX1 gate7005(.O (g10474), .I (g8841));
INVX1 gate7006(.O (g32588), .I (g30825));
INVX1 gate7007(.O (g32524), .I (g31070));
INVX1 gate7008(.O (g9220), .I (g843));
INVX1 gate7009(.O (g31843), .I (g29385));
INVX1 gate7010(.O (g32836), .I (g31021));
INVX1 gate7011(.O (g33696), .I (I31535));
INVX1 gate7012(.O (g30076), .I (g29085));
INVX1 gate7013(.O (g30085), .I (g29082));
INVX1 gate7014(.O (g7851), .I (g921));
INVX1 gate7015(.O (I33075), .I (g34843));
INVX1 gate7016(.O (g9779), .I (g5156));
INVX1 gate7017(.O (g26655), .I (g25492));
INVX1 gate7018(.O (g13637), .I (g10556));
INVX1 gate7019(.O (g20515), .I (g15483));
INVX1 gate7020(.O (g34307), .I (g34087));
INVX1 gate7021(.O (g23041), .I (g19882));
INVX1 gate7022(.O (I20388), .I (g17724));
INVX1 gate7023(.O (g32477), .I (g31566));
INVX1 gate7024(.O (I18360), .I (g1426));
INVX1 gate7025(.O (g21275), .I (g15426));
INVX1 gate7026(.O (g24515), .I (g22689));
INVX1 gate7027(.O (I31494), .I (g33283));
INVX1 gate7028(.O (g24991), .I (g22369));
INVX1 gate7029(.O (I12120), .I (g632));
INVX1 gate7030(.O (g10109), .I (g135));
INVX1 gate7031(.O (g30054), .I (g29134));
INVX1 gate7032(.O (g21430), .I (g15608));
INVX1 gate7033(.O (g27163), .I (I25869));
INVX1 gate7034(.O (g34596), .I (I32696));
INVX1 gate7035(.O (g8406), .I (g232));
INVX1 gate7036(.O (g17756), .I (g14858));
INVX1 gate7037(.O (I27738), .I (g28140));
INVX1 gate7038(.O (g23430), .I (I22547));
INVX1 gate7039(.O (g23746), .I (g20902));
INVX1 gate7040(.O (g23493), .I (g21611));
INVX1 gate7041(.O (g7964), .I (g3155));
INVX1 gate7042(.O (g7260), .I (I11908));
INVX1 gate7043(.O (g8635), .I (g2783));
INVX1 gate7044(.O (g24407), .I (g22594));
INVX1 gate7045(.O (g34243), .I (I32228));
INVX1 gate7046(.O (g29697), .I (g28336));
INVX1 gate7047(.O (g9977), .I (g2667));
INVX1 gate7048(.O (g19481), .I (g16349));
INVX1 gate7049(.O (g10108), .I (g120));
INVX1 gate7050(.O (I14932), .I (g9901));
INVX1 gate7051(.O (g29995), .I (g28955));
INVX1 gate7052(.O (I33037), .I (g34770));
INVX1 gate7053(.O (g34431), .I (I32464));
INVX1 gate7054(.O (g12012), .I (g9213));
INVX1 gate7055(.O (g32118), .I (g31008));
INVX1 gate7056(.O (g15816), .I (I17314));
INVX1 gate7057(.O (g8766), .I (g572));
INVX1 gate7058(.O (g18940), .I (I19719));
INVX1 gate7059(.O (g8087), .I (g1157));
INVX1 gate7060(.O (I31782), .I (g33219));
INVX1 gate7061(.O (g32864), .I (g30937));
INVX1 gate7062(.O (g23237), .I (g20924));
INVX1 gate7063(.O (I19734), .I (g17725));
INVX1 gate7064(.O (g7063), .I (g4831));
INVX1 gate7065(.O (g10606), .I (g10233));
INVX1 gate7066(.O (g21340), .I (I21074));
INVX1 gate7067(.O (g32749), .I (g31021));
INVX1 gate7068(.O (g32616), .I (g30735));
INVX1 gate7069(.O (g23340), .I (g21070));
INVX1 gate7070(.O (g23983), .I (g19210));
INVX1 gate7071(.O (I22128), .I (g19968));
INVX1 gate7072(.O (g34773), .I (I32963));
INVX1 gate7073(.O (g9051), .I (g1426));
INVX1 gate7074(.O (g23684), .I (I22819));
INVX1 gate7075(.O (g25480), .I (g22228));
INVX1 gate7076(.O (g34942), .I (g34928));
INVX1 gate7077(.O (g32748), .I (g31710));
INVX1 gate7078(.O (I15577), .I (g10430));
INVX1 gate7079(.O (g8748), .I (g776));
INVX1 gate7080(.O (g11215), .I (g8285));
INVX1 gate7081(.O (g19127), .I (I19775));
INVX1 gate7082(.O (g9451), .I (g5873));
INVX1 gate7083(.O (g28326), .I (g27414));
INVX1 gate7084(.O (I32991), .I (g34759));
INVX1 gate7085(.O (I14505), .I (g10140));
INVX1 gate7086(.O (I33155), .I (g34897));
INVX1 gate7087(.O (g13215), .I (g10909));
INVX1 gate7088(.O (g26131), .I (I25161));
INVX1 gate7089(.O (g34156), .I (g33907));
INVX1 gate7090(.O (g13729), .I (g10951));
INVX1 gate7091(.O (g25550), .I (g22763));
INVX1 gate7092(.O (g20441), .I (g17873));
INVX1 gate7093(.O (g20584), .I (g17873));
INVX1 gate7094(.O (g32704), .I (g31070));
INVX1 gate7095(.O (I21047), .I (g17429));
INVX1 gate7096(.O (g10381), .I (g6957));
INVX1 gate7097(.O (g28040), .I (g26365));
INVX1 gate7098(.O (g33708), .I (I31555));
INVX1 gate7099(.O (I33170), .I (g34890));
INVX1 gate7100(.O (g19490), .I (g16489));
INVX1 gate7101(.O (g25287), .I (g22228));
INVX1 gate7102(.O (g34670), .I (I32794));
INVX1 gate7103(.O (I29939), .I (g31667));
INVX1 gate7104(.O (g9999), .I (g6109));
INVX1 gate7105(.O (I17128), .I (g13835));
INVX1 gate7106(.O (g23517), .I (g21070));
INVX1 gate7107(.O (g33258), .I (g32296));
INVX1 gate7108(.O (g32809), .I (g31327));
INVX1 gate7109(.O (g32900), .I (g30937));
INVX1 gate7110(.O (g25307), .I (g22763));
INVX1 gate7111(.O (g32466), .I (g31070));
INVX1 gate7112(.O (g7118), .I (g832));
INVX1 gate7113(.O (g7619), .I (g1296));
INVX1 gate7114(.O (g16124), .I (g13555));
INVX1 gate7115(.O (I19487), .I (g15125));
INVX1 gate7116(.O (g19376), .I (g17509));
INVX1 gate7117(.O (g19385), .I (g16326));
INVX1 gate7118(.O (I17626), .I (g14582));
INVX1 gate7119(.O (g17413), .I (I18350));
INVX1 gate7120(.O (g9103), .I (g5774));
INVX1 gate7121(.O (g32808), .I (g30937));
INVX1 gate7122(.O (I26952), .I (g27972));
INVX1 gate7123(.O (g24759), .I (g23003));
INVX1 gate7124(.O (I18071), .I (g13680));
INVX1 gate7125(.O (g19980), .I (g17226));
INVX1 gate7126(.O (g25243), .I (g22763));
INVX1 gate7127(.O (g34839), .I (I33053));
INVX1 gate7128(.O (g17691), .I (I18674));
INVX1 gate7129(.O (g20114), .I (I20385));
INVX1 gate7130(.O (g16686), .I (I17892));
INVX1 gate7131(.O (g34930), .I (I33182));
INVX1 gate7132(.O (g11349), .I (I14365));
INVX1 gate7133(.O (g34993), .I (I33279));
INVX1 gate7134(.O (g12946), .I (I15564));
INVX1 gate7135(.O (g15842), .I (g13469));
INVX1 gate7136(.O (g32560), .I (g31070));
INVX1 gate7137(.O (g20435), .I (g15348));
INVX1 gate7138(.O (g8373), .I (g2485));
INVX1 gate7139(.O (I15906), .I (g10430));
INVX1 gate7140(.O (g24114), .I (g20720));
INVX1 gate7141(.O (g8091), .I (g1579));
INVX1 gate7142(.O (I33167), .I (g34890));
INVX1 gate7143(.O (g6772), .I (I11629));
INVX1 gate7144(.O (g29498), .I (I27784));
INVX1 gate7145(.O (g24082), .I (g19890));
INVX1 gate7146(.O (I15284), .I (g6697));
INVX1 gate7147(.O (g16030), .I (g13570));
INVX1 gate7148(.O (g7393), .I (g5320));
INVX1 gate7149(.O (g13906), .I (I16201));
INVX1 gate7150(.O (g10390), .I (g6987));
INVX1 gate7151(.O (g21362), .I (g17873));
INVX1 gate7152(.O (g24107), .I (g20857));
INVX1 gate7153(.O (g32642), .I (g31542));
INVX1 gate7154(.O (g9732), .I (g5481));
INVX1 gate7155(.O (g23362), .I (I22467));
INVX1 gate7156(.O (g34131), .I (I32074));
INVX1 gate7157(.O (g29056), .I (g27800));
INVX1 gate7158(.O (g22928), .I (I22131));
INVX1 gate7159(.O (g9753), .I (g1890));
INVX1 gate7160(.O (I26516), .I (g26824));
INVX1 gate7161(.O (g23523), .I (g21514));
INVX1 gate7162(.O (g31810), .I (g29385));
INVX1 gate7163(.O (g8283), .I (I12493));
INVX1 gate7164(.O (g25773), .I (g24453));
INVX1 gate7165(.O (I27481), .I (g27928));
INVX1 gate7166(.O (g18833), .I (I19661));
INVX1 gate7167(.O (g31657), .I (I29239));
INVX1 gate7168(.O (g7971), .I (g4818));
INVX1 gate7169(.O (g13304), .I (I15872));
INVX1 gate7170(.O (I20447), .I (g16244));
INVX1 gate7171(.O (I28582), .I (g30116));
INVX1 gate7172(.O (I18825), .I (g6019));
INVX1 gate7173(.O (I18370), .I (g14873));
INVX1 gate7174(.O (g24744), .I (g22202));
INVX1 gate7175(.O (I31477), .I (g33391));
INVX1 gate7176(.O (g29080), .I (g27779));
INVX1 gate7177(.O (g7686), .I (g4659));
INVX1 gate7178(.O (g33375), .I (g32377));
INVX1 gate7179(.O (g8407), .I (g1171));
INVX1 gate7180(.O (g17929), .I (I18855));
INVX1 gate7181(.O (g9072), .I (g2994));
INVX1 gate7182(.O (g25156), .I (g22498));
INVX1 gate7183(.O (I29218), .I (g30304));
INVX1 gate7184(.O (g8920), .I (I12899));
INVX1 gate7185(.O (g8059), .I (g3171));
INVX1 gate7186(.O (g32733), .I (g31672));
INVX1 gate7187(.O (I33119), .I (g34852));
INVX1 gate7188(.O (g14192), .I (g11385));
INVX1 gate7189(.O (I18858), .I (g13835));
INVX1 gate7190(.O (g9472), .I (g6555));
INVX1 gate7191(.O (g19931), .I (g17200));
INVX1 gate7192(.O (g25180), .I (g23529));
INVX1 gate7193(.O (g6856), .I (I11682));
INVX1 gate7194(.O (I12572), .I (g51));
INVX1 gate7195(.O (g15830), .I (g13432));
INVX1 gate7196(.O (g17583), .I (g14968));
INVX1 gate7197(.O (g8718), .I (g3333));
INVX1 gate7198(.O (I18151), .I (g13144));
INVX1 gate7199(.O (g34210), .I (I32173));
INVX1 gate7200(.O (g32874), .I (g30673));
INVX1 gate7201(.O (I28925), .I (g29987));
INVX1 gate7202(.O (g9443), .I (g5489));
INVX1 gate7203(.O (g21727), .I (I21300));
INVX1 gate7204(.O (I22512), .I (g19389));
INVX1 gate7205(.O (g20652), .I (I20744));
INVX1 gate7206(.O (g28508), .I (I26989));
INVX1 gate7207(.O (g32630), .I (g30735));
INVX1 gate7208(.O (g7121), .I (I11820));
INVX1 gate7209(.O (g23863), .I (g19210));
INVX1 gate7210(.O (g32693), .I (g31579));
INVX1 gate7211(.O (I31616), .I (g33219));
INVX1 gate7212(.O (g21222), .I (g17430));
INVX1 gate7213(.O (I23396), .I (g23427));
INVX1 gate7214(.O (g7670), .I (g4104));
INVX1 gate7215(.O (g23222), .I (g20785));
INVX1 gate7216(.O (I18367), .I (g13010));
INVX1 gate7217(.O (g26187), .I (I25190));
INVX1 gate7218(.O (g29342), .I (g28188));
INVX1 gate7219(.O (g9316), .I (g5742));
INVX1 gate7220(.O (g25930), .I (I25028));
INVX1 gate7221(.O (g7625), .I (I12109));
INVX1 gate7222(.O (g32665), .I (g31579));
INVX1 gate7223(.O (I31748), .I (g33228));
INVX1 gate7224(.O (I13473), .I (g4157));
INVX1 gate7225(.O (g19520), .I (g16826));
INVX1 gate7226(.O (g6992), .I (g4899));
INVX1 gate7227(.O (g12760), .I (g10272));
INVX1 gate7228(.O (g9434), .I (g5385));
INVX1 gate7229(.O (g13138), .I (I15765));
INVX1 gate7230(.O (g17787), .I (I18795));
INVX1 gate7231(.O (g7232), .I (g4411));
INVX1 gate7232(.O (g10553), .I (g8971));
INVX1 gate7233(.O (g25838), .I (g25250));
INVX1 gate7234(.O (I27784), .I (g29013));
INVX1 gate7235(.O (I15636), .I (g12075));
INVX1 gate7236(.O (I33276), .I (g34985));
INVX1 gate7237(.O (I33285), .I (g34988));
INVX1 gate7238(.O (g18947), .I (g16136));
INVX1 gate7239(.O (I27385), .I (g27438));
INVX1 gate7240(.O (g30039), .I (g29134));
INVX1 gate7241(.O (g30306), .I (g28796));
INVX1 gate7242(.O (g25131), .I (g23699));
INVX1 gate7243(.O (I33053), .I (g34778));
INVX1 gate7244(.O (g15705), .I (g13217));
INVX1 gate7245(.O (g26937), .I (I25683));
INVX1 gate7246(.O (g17302), .I (I18285));
INVX1 gate7247(.O (g32892), .I (g31021));
INVX1 gate7248(.O (g23347), .I (I22444));
INVX1 gate7249(.O (g24135), .I (g20720));
INVX1 gate7250(.O (g32476), .I (g30673));
INVX1 gate7251(.O (g32485), .I (g31376));
INVX1 gate7252(.O (g33459), .I (I30995));
INVX1 gate7253(.O (I31466), .I (g33318));
INVX1 gate7254(.O (g7909), .I (g936));
INVX1 gate7255(.O (g30038), .I (g29097));
INVX1 gate7256(.O (g23253), .I (g21037));
INVX1 gate7257(.O (I12103), .I (g572));
INVX1 gate7258(.O (g11852), .I (I14668));
INVX1 gate7259(.O (g17743), .I (I18734));
INVX1 gate7260(.O (g9681), .I (g5798));
INVX1 gate7261(.O (I22499), .I (g21160));
INVX1 gate7262(.O (g10040), .I (g2652));
INVX1 gate7263(.O (I22316), .I (g19361));
INVX1 gate7264(.O (g32555), .I (g30673));
INVX1 gate7265(.O (I18446), .I (g13028));
INVX1 gate7266(.O (g14536), .I (I16651));
INVX1 gate7267(.O (g19860), .I (g17226));
INVX1 gate7268(.O (g33458), .I (I30992));
INVX1 gate7269(.O (g7519), .I (g1157));
INVX1 gate7270(.O (g24361), .I (g22885));
INVX1 gate7271(.O (g11963), .I (g9153));
INVX1 gate7272(.O (g25557), .I (g22763));
INVX1 gate7273(.O (g32570), .I (g31554));
INVX1 gate7274(.O (g32712), .I (g30614));
INVX1 gate7275(.O (g25210), .I (g23802));
INVX1 gate7276(.O (g32914), .I (g31672));
INVX1 gate7277(.O (I25351), .I (g24466));
INVX1 gate7278(.O (g9914), .I (g2533));
INVX1 gate7279(.O (I20355), .I (g17613));
INVX1 gate7280(.O (g33918), .I (I31782));
INVX1 gate7281(.O (g23236), .I (g20785));
INVX1 gate7282(.O (g20500), .I (g17873));
INVX1 gate7283(.O (g10621), .I (g7567));
INVX1 gate7284(.O (g34677), .I (I32815));
INVX1 gate7285(.O (g29365), .I (g29067));
INVX1 gate7286(.O (g14252), .I (I16438));
INVX1 gate7287(.O (I22989), .I (g21175));
INVX1 gate7288(.O (g13664), .I (g11252));
INVX1 gate7289(.O (g20049), .I (I20318));
INVX1 gate7290(.O (g23952), .I (g19277));
INVX1 gate7291(.O (g23351), .I (g20924));
INVX1 gate7292(.O (g32907), .I (g30937));
INVX1 gate7293(.O (I31642), .I (g33204));
INVX1 gate7294(.O (g33079), .I (I30641));
INVX1 gate7295(.O (g24049), .I (g20014));
INVX1 gate7296(.O (I14896), .I (g9820));
INVX1 gate7297(.O (g29960), .I (g28885));
INVX1 gate7298(.O (g21175), .I (I20951));
INVX1 gate7299(.O (g22881), .I (I22096));
INVX1 gate7300(.O (g23821), .I (g19210));
INVX1 gate7301(.O (g10564), .I (g9462));
INVX1 gate7302(.O (g15938), .I (I17401));
INVX1 gate7303(.O (g16075), .I (g13597));
INVX1 gate7304(.O (g9413), .I (g1744));
INVX1 gate7305(.O (g19659), .I (g17062));
INVX1 gate7306(.O (g14564), .I (I16679));
INVX1 gate7307(.O (g24048), .I (g19968));
INVX1 gate7308(.O (I11682), .I (g2756));
INVX1 gate7309(.O (g11576), .I (g8542));
INVX1 gate7310(.O (I33064), .I (g34784));
INVX1 gate7311(.O (I25790), .I (g26424));
INVX1 gate7312(.O (I17989), .I (g14173));
INVX1 gate7313(.O (g20004), .I (g17249));
INVX1 gate7314(.O (g13484), .I (g10981));
INVX1 gate7315(.O (g32567), .I (g31070));
INVX1 gate7316(.O (g32594), .I (g30735));
INVX1 gate7317(.O (g19658), .I (g16987));
INVX1 gate7318(.O (g23264), .I (g21037));
INVX1 gate7319(.O (g25286), .I (g22228));
INVX1 gate7320(.O (g16623), .I (g14127));
INVX1 gate7321(.O (g10183), .I (g2595));
INVX1 gate7322(.O (I15609), .I (g12013));
INVX1 gate7323(.O (g7586), .I (I12056));
INVX1 gate7324(.O (g23516), .I (g20924));
INVX1 gate7325(.O (g25039), .I (g22498));
INVX1 gate7326(.O (I28548), .I (g28147));
INVX1 gate7327(.O (g10397), .I (g7018));
INVX1 gate7328(.O (g6976), .I (I11750));
INVX1 gate7329(.O (g14183), .I (g12381));
INVX1 gate7330(.O (g14673), .I (I16770));
INVX1 gate7331(.O (g11609), .I (g7660));
INVX1 gate7332(.O (g9820), .I (g99));
INVX1 gate7333(.O (g16782), .I (I18006));
INVX1 gate7334(.O (g12903), .I (g10411));
INVX1 gate7335(.O (g20613), .I (g15224));
INVX1 gate7336(.O (I21787), .I (g19422));
INVX1 gate7337(.O (I22461), .I (g21225));
INVX1 gate7338(.O (g31817), .I (g29385));
INVX1 gate7339(.O (g13312), .I (g11048));
INVX1 gate7340(.O (I18301), .I (g12976));
INVX1 gate7341(.O (g32941), .I (g30735));
INVX1 gate7342(.O (g32382), .I (g31657));
INVX1 gate7343(.O (g11608), .I (g7659));
INVX1 gate7344(.O (g19644), .I (g17953));
INVX1 gate7345(.O (g10509), .I (g10233));
INVX1 gate7346(.O (I18120), .I (g13350));
INVX1 gate7347(.O (g32519), .I (g30673));
INVX1 gate7348(.O (I22031), .I (g21387));
INVX1 gate7349(.O (I27546), .I (g29041));
INVX1 gate7350(.O (g32185), .I (I29717));
INVX1 gate7351(.O (g18421), .I (I19235));
INVX1 gate7352(.O (g14509), .I (I16626));
INVX1 gate7353(.O (I15921), .I (g12381));
INVX1 gate7354(.O (g32675), .I (g31070));
INVX1 gate7355(.O (g8388), .I (g3010));
INVX1 gate7356(.O (I23357), .I (g23359));
INVX1 gate7357(.O (g20273), .I (g17128));
INVX1 gate7358(.O (g20106), .I (g17328));
INVX1 gate7359(.O (g12563), .I (g9864));
INVX1 gate7360(.O (g20605), .I (g17955));
INVX1 gate7361(.O (g21422), .I (g15373));
INVX1 gate7362(.O (I26409), .I (g26187));
INVX1 gate7363(.O (g30217), .I (I28458));
INVX1 gate7364(.O (g8216), .I (g3092));
INVX1 gate7365(.O (g10851), .I (I14069));
INVX1 gate7366(.O (I12089), .I (g744));
INVX1 gate7367(.O (g10872), .I (g7567));
INVX1 gate7368(.O (g9601), .I (g4005));
INVX1 gate7369(.O (g23422), .I (g21611));
INVX1 gate7370(.O (g32518), .I (g30614));
INVX1 gate7371(.O (I16328), .I (g878));
INVX1 gate7372(.O (g24106), .I (g19984));
INVX1 gate7373(.O (g24605), .I (g23139));
INVX1 gate7374(.O (I14050), .I (g9963));
INVX1 gate7375(.O (g29043), .I (I27391));
INVX1 gate7376(.O (I16538), .I (g10417));
INVX1 gate7377(.O (g13745), .I (I16102));
INVX1 gate7378(.O (g32637), .I (g30735));
INVX1 gate7379(.O (g31656), .I (I29236));
INVX1 gate7380(.O (I20318), .I (g16920));
INVX1 gate7381(.O (g17249), .I (I18265));
INVX1 gate7382(.O (I28002), .I (g28153));
INVX1 gate7383(.O (g32935), .I (g31672));
INVX1 gate7384(.O (g24463), .I (g23578));
INVX1 gate7385(.O (I21769), .I (g19402));
INVX1 gate7386(.O (I17650), .I (g13271));
INVX1 gate7387(.O (I28128), .I (g28314));
INVX1 gate7388(.O (g20033), .I (g16579));
INVX1 gate7389(.O (g31823), .I (g29385));
INVX1 gate7390(.O (I32613), .I (g34329));
INVX1 gate7391(.O (g32883), .I (g30735));
INVX1 gate7392(.O (g17248), .I (I18262));
INVX1 gate7393(.O (I30641), .I (g32024));
INVX1 gate7394(.O (I31555), .I (g33212));
INVX1 gate7395(.O (I14742), .I (g9534));
INVX1 gate7396(.O (g19411), .I (g16489));
INVX1 gate7397(.O (g19527), .I (g16349));
INVX1 gate7398(.O (g17710), .I (g14764));
INVX1 gate7399(.O (g24033), .I (g19919));
INVX1 gate7400(.O (I17198), .I (g13809));
INVX1 gate7401(.O (g12845), .I (g10358));
INVX1 gate7402(.O (g27990), .I (g26770));
INVX1 gate7403(.O (g16853), .I (g13584));
INVX1 gate7404(.O (I12497), .I (g49));
INVX1 gate7405(.O (g23542), .I (g21514));
INVX1 gate7406(.O (g9581), .I (g91));
INVX1 gate7407(.O (g23021), .I (g20283));
INVX1 gate7408(.O (g23453), .I (I22576));
INVX1 gate7409(.O (g10213), .I (g6732));
INVX1 gate7410(.O (I32947), .I (g34659));
INVX1 gate7411(.O (g12899), .I (g10407));
INVX1 gate7412(.O (g21726), .I (I21297));
INVX1 gate7413(.O (g16589), .I (g14082));
INVX1 gate7414(.O (g25169), .I (g22763));
INVX1 gate7415(.O (g29955), .I (g28950));
INVX1 gate7416(.O (g9060), .I (g3355));
INVX1 gate7417(.O (I32106), .I (g33653));
INVX1 gate7418(.O (g23913), .I (g19147));
INVX1 gate7419(.O (g15915), .I (I17392));
INVX1 gate7420(.O (g9460), .I (g6154));
INVX1 gate7421(.O (g24795), .I (g23342));
INVX1 gate7422(.O (g29970), .I (I28199));
INVX1 gate7423(.O (g7659), .I (I12141));
INVX1 gate7424(.O (g12898), .I (g10405));
INVX1 gate7425(.O (g22647), .I (I21959));
INVX1 gate7426(.O (g17778), .I (I18778));
INVX1 gate7427(.O (g16588), .I (g13929));
INVX1 gate7428(.O (g25168), .I (I24334));
INVX1 gate7429(.O (g23614), .I (g20248));
INVX1 gate7430(.O (g25410), .I (g22228));
INVX1 gate7431(.O (g18829), .I (g15171));
INVX1 gate7432(.O (I12987), .I (g12));
INVX1 gate7433(.O (I15732), .I (g6692));
INVX1 gate7434(.O (g8741), .I (g4821));
INVX1 gate7435(.O (g10047), .I (g5421));
INVX1 gate7436(.O (I32812), .I (g34588));
INVX1 gate7437(.O (g19503), .I (g16349));
INVX1 gate7438(.O (g29878), .I (g28421));
INVX1 gate7439(.O (g15277), .I (I17104));
INVX1 gate7440(.O (g21607), .I (g17873));
INVX1 gate7441(.O (g22999), .I (g20453));
INVX1 gate7442(.O (g23607), .I (g21611));
INVX1 gate7443(.O (g21905), .I (I21486));
INVX1 gate7444(.O (g14205), .I (g12381));
INVX1 gate7445(.O (g26654), .I (g25275));
INVX1 gate7446(.O (g20514), .I (g15348));
INVX1 gate7447(.O (I25530), .I (g25222));
INVX1 gate7448(.O (g32501), .I (g30825));
INVX1 gate7449(.O (g32729), .I (g30937));
INVX1 gate7450(.O (g18828), .I (g17955));
INVX1 gate7451(.O (g31631), .I (I29221));
INVX1 gate7452(.O (g10311), .I (g4633));
INVX1 gate7453(.O (g23320), .I (I22419));
INVX1 gate7454(.O (g23905), .I (g21514));
INVX1 gate7455(.O (g9739), .I (g5752));
INVX1 gate7456(.O (g32577), .I (g31554));
INVX1 gate7457(.O (g33631), .I (I31459));
INVX1 gate7458(.O (I14730), .I (g7717));
INVX1 gate7459(.O (g18946), .I (g16100));
INVX1 gate7460(.O (g29171), .I (g27937));
INVX1 gate7461(.O (g21274), .I (g15373));
INVX1 gate7462(.O (g14912), .I (I16917));
INVX1 gate7463(.O (g30321), .I (I28572));
INVX1 gate7464(.O (g23274), .I (g21070));
INVX1 gate7465(.O (g20507), .I (g15509));
INVX1 gate7466(.O (g23530), .I (g20248));
INVX1 gate7467(.O (g22998), .I (g20391));
INVX1 gate7468(.O (g27832), .I (I26409));
INVX1 gate7469(.O (I32234), .I (g34126));
INVX1 gate7470(.O (g34922), .I (I33158));
INVX1 gate7471(.O (I24281), .I (g23440));
INVX1 gate7472(.O (g26936), .I (I25680));
INVX1 gate7473(.O (g15595), .I (I17173));
INVX1 gate7474(.O (g32728), .I (g31021));
INVX1 gate7475(.O (g21346), .I (g17821));
INVX1 gate7476(.O (g25015), .I (g23662));
INVX1 gate7477(.O (g6977), .I (I11753));
INVX1 gate7478(.O (I20957), .I (g16228));
INVX1 gate7479(.O (g19714), .I (g16821));
INVX1 gate7480(.O (I13240), .I (g5794));
INVX1 gate7481(.O (g7275), .I (g1728));
INVX1 gate7482(.O (g22182), .I (I21766));
INVX1 gate7483(.O (g29967), .I (g28946));
INVX1 gate7484(.O (g29994), .I (g29049));
INVX1 gate7485(.O (g34531), .I (I32594));
INVX1 gate7486(.O (g9995), .I (g6035));
INVX1 gate7487(.O (I12644), .I (g3689));
INVX1 gate7488(.O (I11903), .I (g4414));
INVX1 gate7489(.O (g23565), .I (g21562));
INVX1 gate7490(.O (g10072), .I (g9));
INVX1 gate7491(.O (g32438), .I (g30991));
INVX1 gate7492(.O (I14690), .I (g9340));
INVX1 gate7493(.O (g8883), .I (g4709));
INVX1 gate7494(.O (g7615), .I (I12083));
INVX1 gate7495(.O (g12440), .I (g9985));
INVX1 gate7496(.O (g27573), .I (g26667));
INVX1 gate7497(.O (I20562), .I (g16525));
INVX1 gate7498(.O (g25556), .I (g22763));
INVX1 gate7499(.O (g24163), .I (I23333));
INVX1 gate7500(.O (I33176), .I (g34887));
INVX1 gate7501(.O (g7174), .I (g6052));
INVX1 gate7502(.O (g19979), .I (g17226));
INVX1 gate7503(.O (g16748), .I (I17970));
INVX1 gate7504(.O (g7374), .I (g2227));
INVX1 gate7505(.O (g12861), .I (g10367));
INVX1 gate7506(.O (g17651), .I (g14868));
INVX1 gate7507(.O (g17672), .I (g14720));
INVX1 gate7508(.O (g34676), .I (I32812));
INVX1 gate7509(.O (g8217), .I (g3143));
INVX1 gate7510(.O (I16515), .I (g12477));
INVX1 gate7511(.O (I17471), .I (g13394));
INVX1 gate7512(.O (g9390), .I (g5808));
INVX1 gate7513(.O (g21292), .I (I21033));
INVX1 gate7514(.O (g11214), .I (g9602));
INVX1 gate7515(.O (g32906), .I (g31021));
INVX1 gate7516(.O (g7985), .I (g3506));
INVX1 gate7517(.O (g16285), .I (I17612));
INVX1 gate7518(.O (g8466), .I (g1514));
INVX1 gate7519(.O (I19762), .I (g15732));
INVX1 gate7520(.O (g22449), .I (g19597));
INVX1 gate7521(.O (g34654), .I (I32766));
INVX1 gate7522(.O (g20541), .I (g17821));
INVX1 gate7523(.O (I12855), .I (g4311));
INVX1 gate7524(.O (g16305), .I (g13346));
INVX1 gate7525(.O (g10350), .I (g6800));
INVX1 gate7526(.O (g13329), .I (I15893));
INVX1 gate7527(.O (g16053), .I (I17442));
INVX1 gate7528(.O (g9501), .I (g5731));
INVX1 gate7529(.O (g6999), .I (g86));
INVX1 gate7530(.O (g16809), .I (g14387));
INVX1 gate7531(.O (g21409), .I (g18008));
INVX1 gate7532(.O (g22897), .I (g21024));
INVX1 gate7533(.O (g7239), .I (g5033));
INVX1 gate7534(.O (I12411), .I (g4809));
INVX1 gate7535(.O (g23409), .I (g21514));
INVX1 gate7536(.O (g8165), .I (g3530));
INVX1 gate7537(.O (g32622), .I (g31376));
INVX1 gate7538(.O (g8571), .I (g57));
INVX1 gate7539(.O (g8365), .I (g2060));
INVX1 gate7540(.O (I26381), .I (g26851));
INVX1 gate7541(.O (g24789), .I (g23309));
INVX1 gate7542(.O (g32566), .I (g30825));
INVX1 gate7543(.O (g19741), .I (g16987));
INVX1 gate7544(.O (I30537), .I (g32027));
INVX1 gate7545(.O (g29079), .I (g27742));
INVX1 gate7546(.O (g7380), .I (g2331));
INVX1 gate7547(.O (g21408), .I (g15373));
INVX1 gate7548(.O (g10152), .I (g2122));
INVX1 gate7549(.O (g7591), .I (g6668));
INVX1 gate7550(.O (g23408), .I (g21468));
INVX1 gate7551(.O (g8055), .I (g1236));
INVX1 gate7552(.O (g10396), .I (g6997));
INVX1 gate7553(.O (g20325), .I (g15171));
INVX1 gate7554(.O (g24359), .I (g22550));
INVX1 gate7555(.O (g19067), .I (g15979));
INVX1 gate7556(.O (g20920), .I (g15426));
INVX1 gate7557(.O (g20535), .I (g17847));
INVX1 gate7558(.O (I13990), .I (g7636));
INVX1 gate7559(.O (g20434), .I (g18065));
INVX1 gate7560(.O (g9704), .I (g2575));
INVX1 gate7561(.O (g31816), .I (g29385));
INVX1 gate7562(.O (g8133), .I (g4809));
INVX1 gate7563(.O (g24920), .I (I24089));
INVX1 gate7564(.O (g24535), .I (g22942));
INVX1 gate7565(.O (I18376), .I (g14332));
INVX1 gate7566(.O (g24358), .I (g22550));
INVX1 gate7567(.O (I18297), .I (g1418));
INVX1 gate7568(.O (I12503), .I (g215));
INVX1 gate7569(.O (g17505), .I (g14899));
INVX1 gate7570(.O (g17404), .I (I18337));
INVX1 gate7571(.O (g10413), .I (g7110));
INVX1 gate7572(.O (g8774), .I (g781));
INVX1 gate7573(.O (g32653), .I (g30825));
INVX1 gate7574(.O (g19801), .I (I20216));
INVX1 gate7575(.O (I32473), .I (g34248));
INVX1 gate7576(.O (g17717), .I (g14937));
INVX1 gate7577(.O (I17879), .I (g14386));
INVX1 gate7578(.O (g34423), .I (g34222));
INVX1 gate7579(.O (g15588), .I (I17166));
INVX1 gate7580(.O (I22886), .I (g18926));
INVX1 gate7581(.O (g32138), .I (g31233));
INVX1 gate7582(.O (I17970), .I (g4027));
INVX1 gate7583(.O (I20895), .I (g16954));
INVX1 gate7584(.O (g24121), .I (g20720));
INVX1 gate7585(.O (I18888), .I (g16644));
INVX1 gate7586(.O (g8396), .I (g3401));
INVX1 gate7587(.O (g9250), .I (g1600));
INVX1 gate7588(.O (g34587), .I (I32671));
INVX1 gate7589(.O (I13718), .I (g890));
INVX1 gate7590(.O (g12997), .I (g11826));
INVX1 gate7591(.O (g10405), .I (g7064));
INVX1 gate7592(.O (g32636), .I (g31376));
INVX1 gate7593(.O (I23998), .I (g22182));
INVX1 gate7594(.O (I32788), .I (g34577));
INVX1 gate7595(.O (g32415), .I (g31591));
INVX1 gate7596(.O (g14405), .I (g12170));
INVX1 gate7597(.O (g19695), .I (g17015));
INVX1 gate7598(.O (g8538), .I (g3412));
INVX1 gate7599(.O (I12819), .I (g4277));
INVX1 gate7600(.O (g29977), .I (g28920));
INVX1 gate7601(.O (I12910), .I (g4340));
INVX1 gate7602(.O (g16874), .I (I18066));
INVX1 gate7603(.O (g32852), .I (g30614));
INVX1 gate7604(.O (g11235), .I (I14301));
INVX1 gate7605(.O (I32535), .I (g34296));
INVX1 gate7606(.O (I25327), .I (g24641));
INVX1 gate7607(.O (g8509), .I (g4141));
INVX1 gate7608(.O (g35002), .I (I33300));
INVX1 gate7609(.O (g19526), .I (g16349));
INVX1 gate7610(.O (g16630), .I (g14142));
INVX1 gate7611(.O (g16693), .I (I17901));
INVX1 gate7612(.O (g26814), .I (g25221));
INVX1 gate7613(.O (g34543), .I (g34359));
INVX1 gate7614(.O (I22425), .I (g19379));
INVX1 gate7615(.O (g24173), .I (I23363));
INVX1 gate7616(.O (g32963), .I (g30825));
INVX1 gate7617(.O (g22148), .I (g19074));
INVX1 gate7618(.O (g7515), .I (I12000));
INVX1 gate7619(.O (g12871), .I (g10378));
INVX1 gate7620(.O (g29353), .I (I27713));
INVX1 gate7621(.O (I12070), .I (g785));
INVX1 gate7622(.O (I22458), .I (g18954));
INVX1 gate7623(.O (g23537), .I (g20785));
INVX1 gate7624(.O (g9568), .I (g6181));
INVX1 gate7625(.O (g31842), .I (g29385));
INVX1 gate7626(.O (g32664), .I (g31528));
INVX1 gate7627(.O (g30569), .I (I28838));
INVX1 gate7628(.O (I16345), .I (g881));
INVX1 gate7629(.O (g8418), .I (g2619));
INVX1 gate7630(.O (I19772), .I (g17818));
INVX1 gate7631(.O (g34569), .I (I32639));
INVX1 gate7632(.O (g22646), .I (g19389));
INVX1 gate7633(.O (I22918), .I (g21451));
INVX1 gate7634(.O (g17433), .I (I18382));
INVX1 gate7635(.O (I25606), .I (g25465));
INVX1 gate7636(.O (g8290), .I (g218));
INVX1 gate7637(.O (I17425), .I (g13416));
INVX1 gate7638(.O (g18903), .I (g15758));
INVX1 gate7639(.O (g30568), .I (g29339));
INVX1 gate7640(.O (g23283), .I (g20785));
INVX1 gate7641(.O (g19866), .I (g16540));
INVX1 gate7642(.O (g11991), .I (g9485));
INVX1 gate7643(.O (I17919), .I (g14609));
INVX1 gate7644(.O (g13414), .I (g11048));
INVX1 gate7645(.O (I22444), .I (g19626));
INVX1 gate7646(.O (g23492), .I (g21562));
INVX1 gate7647(.O (g25423), .I (I24558));
INVX1 gate7648(.O (g23303), .I (g20785));
INVX1 gate7649(.O (I31622), .I (g33204));
INVX1 gate7650(.O (g32576), .I (g30614));
INVX1 gate7651(.O (g24134), .I (g19984));
INVX1 gate7652(.O (g8093), .I (g1624));
INVX1 gate7653(.O (g32484), .I (g31566));
INVX1 gate7654(.O (g34242), .I (I32225));
INVX1 gate7655(.O (g24029), .I (g20982));
INVX1 gate7656(.O (g33424), .I (g32415));
INVX1 gate7657(.O (I11701), .I (g4164));
INVX1 gate7658(.O (g10113), .I (g2084));
INVX1 gate7659(.O (g17811), .I (g12925));
INVX1 gate7660(.O (g17646), .I (I18609));
INVX1 gate7661(.O (I11777), .I (g5357));
INVX1 gate7662(.O (g20506), .I (g15426));
INVX1 gate7663(.O (I28199), .I (g28803));
INVX1 gate7664(.O (I25750), .I (g26823));
INVX1 gate7665(.O (g20028), .I (g15371));
INVX1 gate7666(.O (I12067), .I (g739));
INVX1 gate7667(.O (I32173), .I (g33645));
INVX1 gate7668(.O (g32554), .I (g30614));
INVX1 gate7669(.O (I18089), .I (g13144));
INVX1 gate7670(.O (g24506), .I (I23711));
INVX1 gate7671(.O (I20385), .I (g16194));
INVX1 gate7672(.O (g7750), .I (g1070));
INVX1 gate7673(.O (g24028), .I (g20841));
INVX1 gate7674(.O (I24784), .I (g24265));
INVX1 gate7675(.O (g34123), .I (I32062));
INVX1 gate7676(.O (g16712), .I (g13223));
INVX1 gate7677(.O (g26841), .I (g24893));
INVX1 gate7678(.O (g32609), .I (g30735));
INVX1 gate7679(.O (g21381), .I (g18008));
INVX1 gate7680(.O (I27735), .I (g28779));
INVX1 gate7681(.O (I29239), .I (g29498));
INVX1 gate7682(.O (g31830), .I (g29385));
INVX1 gate7683(.O (g23982), .I (g19147));
INVX1 gate7684(.O (g10357), .I (g6825));
INVX1 gate7685(.O (g26510), .I (I25369));
INVX1 gate7686(.O (g14357), .I (g12181));
INVX1 gate7687(.O (g34772), .I (I32960));
INVX1 gate7688(.O (I12735), .I (g4572));
INVX1 gate7689(.O (g8181), .I (g424));
INVX1 gate7690(.O (g28779), .I (I27253));
INVX1 gate7691(.O (g32608), .I (g31376));
INVX1 gate7692(.O (g8381), .I (g2610));
INVX1 gate7693(.O (g19689), .I (g16795));
INVX1 gate7694(.O (g7040), .I (g4821));
INVX1 gate7695(.O (g25117), .I (g22417));
INVX1 gate7696(.O (I16135), .I (g10430));
INVX1 gate7697(.O (g25000), .I (g23630));
INVX1 gate7698(.O (g8685), .I (g1430));
INVX1 gate7699(.O (g7440), .I (g329));
INVX1 gate7700(.O (g8700), .I (g4054));
INVX1 gate7701(.O (g28081), .I (I26584));
INVX1 gate7702(.O (g32921), .I (g31672));
INVX1 gate7703(.O (g33713), .I (I31564));
INVX1 gate7704(.O (g8397), .I (g3470));
INVX1 gate7705(.O (g19688), .I (g16777));
INVX1 gate7706(.O (g9626), .I (g6466));
INVX1 gate7707(.O (g8021), .I (g3512));
INVX1 gate7708(.O (g16594), .I (I17772));
INVX1 gate7709(.O (g26835), .I (I25555));
INVX1 gate7710(.O (g13584), .I (g12735));
INVX1 gate7711(.O (g18990), .I (g16136));
INVX1 gate7712(.O (g32745), .I (g31376));
INVX1 gate7713(.O (I29185), .I (g30012));
INVX1 gate7714(.O (g22896), .I (g21012));
INVX1 gate7715(.O (I18700), .I (g6027));
INVX1 gate7716(.O (g23840), .I (g19074));
INVX1 gate7717(.O (g15733), .I (I17249));
INVX1 gate7718(.O (g32799), .I (g31710));
INVX1 gate7719(.O (g18898), .I (g15566));
INVX1 gate7720(.O (g23390), .I (g21468));
INVX1 gate7721(.O (g32813), .I (g31710));
INVX1 gate7722(.O (g22228), .I (I21810));
INVX1 gate7723(.O (g6820), .I (g1070));
INVX1 gate7724(.O (g33705), .I (I31550));
INVX1 gate7725(.O (g25242), .I (g23684));
INVX1 gate7726(.O (g7666), .I (g4076));
INVX1 gate7727(.O (I17159), .I (g13350));
INVX1 gate7728(.O (g20649), .I (g18065));
INVX1 gate7729(.O (I17125), .I (g13809));
INVX1 gate7730(.O (I22561), .I (g20841));
INVX1 gate7731(.O (I23149), .I (g19061));
INVX1 gate7732(.O (g31189), .I (I29002));
INVX1 gate7733(.O (g34992), .I (I33276));
INVX1 gate7734(.O (I17901), .I (g3976));
INVX1 gate7735(.O (g34391), .I (g34200));
INVX1 gate7736(.O (g32798), .I (g31672));
INVX1 gate7737(.O (I22353), .I (g19375));
INVX1 gate7738(.O (g28380), .I (g27064));
INVX1 gate7739(.O (g20240), .I (g17847));
INVX1 gate7740(.O (I23387), .I (g23394));
INVX1 gate7741(.O (g32973), .I (g31021));
INVX1 gate7742(.O (I30904), .I (g32424));
INVX1 gate7743(.O (g34510), .I (g34418));
INVX1 gate7744(.O (g22716), .I (g19795));
INVX1 gate7745(.O (g23192), .I (g20248));
INVX1 gate7746(.O (g16675), .I (I17873));
INVX1 gate7747(.O (g20648), .I (g15615));
INVX1 gate7748(.O (g10881), .I (g7567));
INVX1 gate7749(.O (I17783), .I (g13304));
INVX1 gate7750(.O (g20903), .I (g17249));
INVX1 gate7751(.O (g32805), .I (g31672));
INVX1 gate7752(.O (g13082), .I (g10981));
INVX1 gate7753(.O (g32674), .I (g30735));
INVX1 gate7754(.O (g24648), .I (g23148));
INVX1 gate7755(.O (g7528), .I (g930));
INVX1 gate7756(.O (g12859), .I (g10366));
INVX1 gate7757(.O (g13107), .I (g10476));
INVX1 gate7758(.O (g34579), .I (I32659));
INVX1 gate7759(.O (g7648), .I (I12135));
INVX1 gate7760(.O (g26615), .I (g25432));
INVX1 gate7761(.O (g12950), .I (g12708));
INVX1 gate7762(.O (g20604), .I (g17873));
INVX1 gate7763(.O (g9683), .I (g6140));
INVX1 gate7764(.O (g23522), .I (g21514));
INVX1 gate7765(.O (g18832), .I (g15634));
INVX1 gate7766(.O (I13360), .I (g5343));
INVX1 gate7767(.O (g24604), .I (g23112));
INVX1 gate7768(.O (g30578), .I (g29956));
INVX1 gate7769(.O (g33460), .I (I30998));
INVX1 gate7770(.O (g33686), .I (g33187));
INVX1 gate7771(.O (g19885), .I (g17249));
INVX1 gate7772(.O (g26720), .I (g25275));
INVX1 gate7773(.O (g7655), .I (g4332));
INVX1 gate7774(.O (g11744), .I (I14602));
INVX1 gate7775(.O (g20770), .I (g17955));
INVX1 gate7776(.O (I26508), .I (g26814));
INVX1 gate7777(.O (g9778), .I (g5069));
INVX1 gate7778(.O (I14271), .I (g8456));
INVX1 gate7779(.O (g20563), .I (g15171));
INVX1 gate7780(.O (g27996), .I (I26508));
INVX1 gate7781(.O (g32732), .I (g30825));
INVX1 gate7782(.O (g24770), .I (g22763));
INVX1 gate7783(.O (g8631), .I (g283));
INVX1 gate7784(.O (g25230), .I (g23314));
INVX1 gate7785(.O (g32934), .I (g30735));
INVX1 gate7786(.O (g24981), .I (g22763));
INVX1 gate7787(.O (I24089), .I (g22409));
INVX1 gate7788(.O (g11849), .I (g7601));
INVX1 gate7789(.O (I16613), .I (g10430));
INVX1 gate7790(.O (g17582), .I (g14768));
INVX1 gate7791(.O (g12996), .I (g11823));
INVX1 gate7792(.O (g10027), .I (g6523));
INVX1 gate7793(.O (g23483), .I (g18833));
INVX1 gate7794(.O (I18060), .I (g14198));
INVX1 gate7795(.O (I23369), .I (g23347));
INVX1 gate7796(.O (g14662), .I (I16762));
INVX1 gate7797(.O (g8301), .I (g1399));
INVX1 gate7798(.O (g19763), .I (g16431));
INVX1 gate7799(.O (g25265), .I (I24455));
INVX1 gate7800(.O (I32240), .I (g34131));
INVX1 gate7801(.O (g29976), .I (g29018));
INVX1 gate7802(.O (g12844), .I (g10360));
INVX1 gate7803(.O (g7410), .I (g2008));
INVX1 gate7804(.O (g11398), .I (I14409));
INVX1 gate7805(.O (g23862), .I (g19147));
INVX1 gate7806(.O (g12367), .I (I15205));
INVX1 gate7807(.O (g32692), .I (g31528));
INVX1 gate7808(.O (g32761), .I (g30825));
INVX1 gate7809(.O (I32648), .I (g34371));
INVX1 gate7810(.O (g18926), .I (I19707));
INVX1 gate7811(.O (I18855), .I (g13745));
INVX1 gate7812(.O (I11629), .I (g19));
INVX1 gate7813(.O (g11652), .I (g7674));
INVX1 gate7814(.O (g9661), .I (g3661));
INVX1 gate7815(.O (g13141), .I (g11374));
INVX1 gate7816(.O (g29374), .I (I27742));
INVX1 gate7817(.O (g20767), .I (g17873));
INVX1 gate7818(.O (g26340), .I (g24953));
INVX1 gate7819(.O (g21326), .I (I21058));
INVX1 gate7820(.O (g18099), .I (I18903));
INVX1 gate7821(.O (I18411), .I (g13018));
INVX1 gate7822(.O (g30116), .I (I28349));
INVX1 gate7823(.O (I14650), .I (g9340));
INVX1 gate7824(.O (g33875), .I (I31727));
INVX1 gate7825(.O (I24497), .I (g22592));
INVX1 gate7826(.O (g10710), .I (I14006));
INVX1 gate7827(.O (g20899), .I (I20861));
INVX1 gate7828(.O (I12300), .I (g1157));
INVX1 gate7829(.O (g10003), .I (I13539));
INVX1 gate7830(.O (g23948), .I (g21012));
INVX1 gate7831(.O (I32770), .I (g34505));
INVX1 gate7832(.O (g18098), .I (I18900));
INVX1 gate7833(.O (g10204), .I (g2685));
INVX1 gate7834(.O (I29438), .I (g30610));
INVX1 gate7835(.O (g21904), .I (I21483));
INVX1 gate7836(.O (g14204), .I (g12155));
INVX1 gate7837(.O (g16577), .I (I17747));
INVX1 gate7838(.O (g20633), .I (g15171));
INVX1 gate7839(.O (g23904), .I (g18997));
INVX1 gate7840(.O (I16371), .I (g887));
INVX1 gate7841(.O (g31837), .I (g29385));
INVX1 gate7842(.O (g14779), .I (I16847));
INVX1 gate7843(.O (g21252), .I (g15656));
INVX1 gate7844(.O (I22289), .I (g19446));
INVX1 gate7845(.O (g32329), .I (g31522));
INVX1 gate7846(.O (g29669), .I (I27941));
INVX1 gate7847(.O (g34275), .I (g34047));
INVX1 gate7848(.O (g19480), .I (g16349));
INVX1 gate7849(.O (g23252), .I (I22353));
INVX1 gate7850(.O (g17603), .I (g14993));
INVX1 gate7851(.O (g20191), .I (g17821));
INVX1 gate7852(.O (g34430), .I (I32461));
INVX1 gate7853(.O (g17742), .I (g14971));
INVX1 gate7854(.O (g32539), .I (g31170));
INVX1 gate7855(.O (g10081), .I (g2279));
INVX1 gate7856(.O (g17096), .I (I18168));
INVX1 gate7857(.O (I18894), .I (g16708));
INVX1 gate7858(.O (g6995), .I (g4944));
INVX1 gate7859(.O (g7618), .I (I12092));
INVX1 gate7860(.O (g8441), .I (g3361));
INVX1 gate7861(.O (g22857), .I (g20739));
INVX1 gate7862(.O (I22571), .I (g20097));
INVX1 gate7863(.O (I11785), .I (g5703));
INVX1 gate7864(.O (g7235), .I (g4521));
INVX1 gate7865(.O (g7343), .I (g5290));
INVX1 gate7866(.O (I14365), .I (g3303));
INVX1 gate7867(.O (g30237), .I (I28480));
INVX1 gate7868(.O (I16795), .I (g5637));
INVX1 gate7869(.O (g25007), .I (g22457));
INVX1 gate7870(.O (g32538), .I (g31070));
INVX1 gate7871(.O (g24718), .I (g22182));
INVX1 gate7872(.O (I32794), .I (g34580));
INVX1 gate7873(.O (g14786), .I (g12471));
INVX1 gate7874(.O (g29195), .I (I27495));
INVX1 gate7875(.O (g9484), .I (g1612));
INVX1 gate7876(.O (g30983), .I (g29657));
INVX1 gate7877(.O (g9439), .I (g5428));
INVX1 gate7878(.O (g17681), .I (g14735));
INVX1 gate7879(.O (g7566), .I (I12049));
INVX1 gate7880(.O (g6840), .I (g1992));
INVX1 gate7881(.O (g8673), .I (g4737));
INVX1 gate7882(.O (g16349), .I (I17661));
INVX1 gate7883(.O (g34983), .I (I33249));
INVX1 gate7884(.O (g18997), .I (I19756));
INVX1 gate7885(.O (g10356), .I (g6819));
INVX1 gate7886(.O (g33455), .I (I30983));
INVX1 gate7887(.O (g21183), .I (g15509));
INVX1 gate7888(.O (g21673), .I (I21234));
INVX1 gate7889(.O (g7693), .I (g4849));
INVX1 gate7890(.O (g11833), .I (g8026));
INVX1 gate7891(.O (g17429), .I (I18370));
INVX1 gate7892(.O (g7134), .I (g5029));
INVX1 gate7893(.O (g21397), .I (g15171));
INVX1 gate7894(.O (g23847), .I (g19210));
INVX1 gate7895(.O (g13049), .I (I15677));
INVX1 gate7896(.O (g10380), .I (g6960));
INVX1 gate7897(.O (g30142), .I (g28754));
INVX1 gate7898(.O (g18061), .I (g14800));
INVX1 gate7899(.O (g16284), .I (I17609));
INVX1 gate7900(.O (g19431), .I (g16249));
INVX1 gate7901(.O (g34142), .I (I32089));
INVX1 gate7902(.O (g25116), .I (g22369));
INVX1 gate7903(.O (g17428), .I (I18367));
INVX1 gate7904(.O (I22816), .I (g19862));
INVX1 gate7905(.O (g7548), .I (g1036));
INVX1 gate7906(.O (g11048), .I (I14158));
INVX1 gate7907(.O (g8669), .I (g3767));
INVX1 gate7908(.O (g10090), .I (g5348));
INVX1 gate7909(.O (g20573), .I (g17384));
INVX1 gate7910(.O (g10233), .I (I13699));
INVX1 gate7911(.O (g20247), .I (g17015));
INVX1 gate7912(.O (g29893), .I (g28755));
INVX1 gate7913(.O (I24060), .I (g22202));
INVX1 gate7914(.O (g16622), .I (g14104));
INVX1 gate7915(.O (g23509), .I (g21611));
INVX1 gate7916(.O (g10182), .I (g2681));
INVX1 gate7917(.O (g28620), .I (g27679));
INVX1 gate7918(.O (I21959), .I (g20242));
INVX1 gate7919(.O (g20389), .I (g15277));
INVX1 gate7920(.O (g8058), .I (g3115));
INVX1 gate7921(.O (I14708), .I (g9417));
INVX1 gate7922(.O (I28458), .I (g28443));
INVX1 gate7923(.O (I29139), .I (g29382));
INVX1 gate7924(.O (g8531), .I (g3288));
INVX1 gate7925(.O (g19773), .I (g17615));
INVX1 gate7926(.O (g24389), .I (g22908));
INVX1 gate7927(.O (g8458), .I (g294));
INVX1 gate7928(.O (g24045), .I (g21193));
INVX1 gate7929(.O (g12902), .I (g10409));
INVX1 gate7930(.O (g20612), .I (g18008));
INVX1 gate7931(.O (g23508), .I (g21562));
INVX1 gate7932(.O (I16163), .I (g11930));
INVX1 gate7933(.O (I20870), .I (g16216));
INVX1 gate7934(.O (g32771), .I (g31021));
INVX1 gate7935(.O (g8743), .I (g550));
INVX1 gate7936(.O (g20388), .I (g17297));
INVX1 gate7937(.O (g20324), .I (g17955));
INVX1 gate7938(.O (g8890), .I (g376));
INVX1 gate7939(.O (I23378), .I (g23426));
INVX1 gate7940(.O (g29713), .I (I27970));
INVX1 gate7941(.O (g24099), .I (g20720));
INVX1 gate7942(.O (g24388), .I (g22885));
INVX1 gate7943(.O (g20701), .I (g17955));
INVX1 gate7944(.O (g20777), .I (g15224));
INVX1 gate7945(.O (g20534), .I (g17183));
INVX1 gate7946(.O (g22317), .I (g19801));
INVX1 gate7947(.O (g31623), .I (g29669));
INVX1 gate7948(.O (g32683), .I (g30614));
INVX1 gate7949(.O (I17976), .I (g13638));
INVX1 gate7950(.O (g25465), .I (g23824));
INVX1 gate7951(.O (g19670), .I (g16897));
INVX1 gate7952(.O (g24534), .I (g22670));
INVX1 gate7953(.O (g8505), .I (g3480));
INVX1 gate7954(.O (g20272), .I (g17239));
INVX1 gate7955(.O (g34130), .I (I32071));
INVX1 gate7956(.O (g24098), .I (g19984));
INVX1 gate7957(.O (g14331), .I (I16489));
INVX1 gate7958(.O (g12738), .I (g9374));
INVX1 gate7959(.O (I19863), .I (g16675));
INVX1 gate7960(.O (g9616), .I (g5452));
INVX1 gate7961(.O (g17504), .I (g15021));
INVX1 gate7962(.O (I16541), .I (g11929));
INVX1 gate7963(.O (g8011), .I (g3167));
INVX1 gate7964(.O (g25340), .I (g22763));
INVX1 gate7965(.O (g25035), .I (g23699));
INVX1 gate7966(.O (I17374), .I (g13638));
INVX1 gate7967(.O (g8411), .I (I12577));
INVX1 gate7968(.O (g8734), .I (g4045));
INVX1 gate7969(.O (g19734), .I (g16861));
INVX1 gate7970(.O (g13106), .I (g10981));
INVX1 gate7971(.O (g27698), .I (g26648));
INVX1 gate7972(.O (g29042), .I (I27388));
INVX1 gate7973(.O (g13605), .I (I16040));
INVX1 gate7974(.O (g10897), .I (g7601));
INVX1 gate7975(.O (I33214), .I (g34954));
INVX1 gate7976(.O (I20867), .I (g16216));
INVX1 gate7977(.O (I27314), .I (g28009));
INVX1 gate7978(.O (g6954), .I (g4138));
INVX1 gate7979(.O (g19930), .I (g17200));
INVX1 gate7980(.O (g6810), .I (g723));
INVX1 gate7981(.O (g9527), .I (g6500));
INVX1 gate7982(.O (I14069), .I (g9104));
INVX1 gate7983(.O (g11812), .I (g7567));
INVX1 gate7984(.O (g7202), .I (g4639));
INVX1 gate7985(.O (I16724), .I (g12108));
INVX1 gate7986(.O (g10404), .I (g7026));
INVX1 gate7987(.O (I12314), .I (g1500));
INVX1 gate7988(.O (g13463), .I (g10476));
INVX1 gate7989(.O (g31822), .I (g29385));
INVX1 gate7990(.O (g32515), .I (g30825));
INVX1 gate7991(.O (I31539), .I (g33212));
INVX1 gate7992(.O (g32882), .I (g31376));
INVX1 gate7993(.O (I14602), .I (g9340));
INVX1 gate7994(.O (I15033), .I (g10273));
INVX1 gate7995(.O (g19694), .I (g16429));
INVX1 gate7996(.O (g7908), .I (g4157));
INVX1 gate7997(.O (I32388), .I (g34153));
INVX1 gate7998(.O (g24032), .I (g21256));
INVX1 gate7999(.O (g22626), .I (I21941));
INVX1 gate8000(.O (I21802), .I (g21308));
INVX1 gate8001(.O (I16829), .I (g6715));
INVX1 gate8002(.O (g25517), .I (g22228));
INVX1 gate8003(.O (g11033), .I (g8500));
INVX1 gate8004(.O (g11371), .I (g7565));
INVX1 gate8005(.O (I16535), .I (g11235));
INVX1 gate8006(.O (g18911), .I (g15169));
INVX1 gate8007(.O (g23452), .I (g21468));
INVX1 gate8008(.O (g10026), .I (g6494));
INVX1 gate8009(.O (g32407), .I (I29939));
INVX1 gate8010(.O (g9546), .I (g2437));
INVX1 gate8011(.O (g13033), .I (g11917));
INVX1 gate8012(.O (g21205), .I (g15656));
INVX1 gate8013(.O (g11234), .I (g8355));
INVX1 gate8014(.O (g10212), .I (g6390));
INVX1 gate8015(.O (I14970), .I (g9965));
INVX1 gate8016(.O (g29939), .I (g28857));
INVX1 gate8017(.O (g17128), .I (I18180));
INVX1 gate8018(.O (g7518), .I (g1024));
INVX1 gate8019(.O (I17668), .I (g13279));
INVX1 gate8020(.O (I20819), .I (g17088));
INVX1 gate8021(.O (I22525), .I (g19345));
INVX1 gate8022(.O (I22488), .I (g18984));
INVX1 gate8023(.O (I17842), .I (g13051));
INVX1 gate8024(.O (I20910), .I (g17197));
INVX1 gate8025(.O (g16963), .I (I18117));
INVX1 gate8026(.O (g23912), .I (g19147));
INVX1 gate8027(.O (I17392), .I (g13680));
INVX1 gate8028(.O (g34222), .I (I32195));
INVX1 gate8029(.O (g9970), .I (g1714));
INVX1 gate8030(.O (g24061), .I (g19919));
INVX1 gate8031(.O (I29585), .I (g31655));
INVX1 gate8032(.O (g29093), .I (g27858));
INVX1 gate8033(.O (g34437), .I (I32482));
INVX1 gate8034(.O (g20766), .I (g17433));
INVX1 gate8035(.O (I26929), .I (g27980));
INVX1 gate8036(.O (g8080), .I (g3863));
INVX1 gate8037(.O (I18526), .I (g13055));
INVX1 gate8038(.O (g31853), .I (g29385));
INVX1 gate8039(.O (g19502), .I (g15674));
INVX1 gate8040(.O (g8480), .I (g3147));
INVX1 gate8041(.O (g19210), .I (I19796));
INVX1 gate8042(.O (g17533), .I (I18482));
INVX1 gate8043(.O (g25193), .I (g22763));
INVX1 gate8044(.O (g8713), .I (g4826));
INVX1 gate8045(.O (g21051), .I (g15171));
INVX1 gate8046(.O (g7593), .I (I12061));
INVX1 gate8047(.O (I17488), .I (g13394));
INVX1 gate8048(.O (g15348), .I (I17111));
INVX1 gate8049(.O (g19618), .I (g16349));
INVX1 gate8050(.O (g19443), .I (g16449));
INVX1 gate8051(.O (I14967), .I (g9964));
INVX1 gate8052(.O (g12895), .I (g10403));
INVX1 gate8053(.O (I12773), .I (g4204));
INVX1 gate8054(.O (g16585), .I (g14075));
INVX1 gate8055(.O (g13514), .I (I15987));
INVX1 gate8056(.O (g25523), .I (g22550));
INVX1 gate8057(.O (g31836), .I (g29385));
INVX1 gate8058(.O (g32441), .I (I29969));
INVX1 gate8059(.O (g32584), .I (g30673));
INVX1 gate8060(.O (I32997), .I (g34760));
INVX1 gate8061(.O (g24360), .I (g22228));
INVX1 gate8062(.O (g29219), .I (I27573));
INVX1 gate8063(.O (g15566), .I (I17143));
INVX1 gate8064(.O (g20447), .I (g15426));
INVX1 gate8065(.O (g14149), .I (g12381));
INVX1 gate8066(.O (g10387), .I (g6996));
INVX1 gate8067(.O (g16609), .I (g14454));
INVX1 gate8068(.O (g19469), .I (g16326));
INVX1 gate8069(.O (I28336), .I (g29147));
INVX1 gate8070(.O (g10620), .I (g10233));
INVX1 gate8071(.O (g17737), .I (g14810));
INVX1 gate8072(.O (g22856), .I (g20453));
INVX1 gate8073(.O (g29218), .I (I27570));
INVX1 gate8074(.O (g22995), .I (g20330));
INVX1 gate8075(.O (g32759), .I (g31376));
INVX1 gate8076(.O (g16200), .I (g13584));
INVX1 gate8077(.O (I33235), .I (g34957));
INVX1 gate8078(.O (g23350), .I (g20785));
INVX1 gate8079(.O (g25006), .I (g22417));
INVX1 gate8080(.O (g32725), .I (g30825));
INVX1 gate8081(.O (g24162), .I (I23330));
INVX1 gate8082(.O (I32766), .I (g34522));
INVX1 gate8083(.O (g7933), .I (g907));
INVX1 gate8084(.O (g16608), .I (g14116));
INVX1 gate8085(.O (g19468), .I (g15938));
INVX1 gate8086(.O (g9617), .I (I13240));
INVX1 gate8087(.O (g23820), .I (g19147));
INVX1 gate8088(.O (g34952), .I (g34942));
INVX1 gate8089(.O (g34351), .I (g34174));
INVX1 gate8090(.O (g13012), .I (I15626));
INVX1 gate8091(.O (g32758), .I (g31327));
INVX1 gate8092(.O (g7521), .I (g5630));
INVX1 gate8093(.O (I32871), .I (g34521));
INVX1 gate8094(.O (g25222), .I (I24400));
INVX1 gate8095(.O (g7050), .I (g5845));
INVX1 gate8096(.O (g20629), .I (g17955));
INVX1 gate8097(.O (g23152), .I (g20283));
INVX1 gate8098(.O (I12930), .I (g4349));
INVX1 gate8099(.O (I13699), .I (g4581));
INVX1 gate8100(.O (g9516), .I (g6116));
INVX1 gate8101(.O (I21002), .I (g16709));
INVX1 gate8102(.O (g20451), .I (g15277));
INVX1 gate8103(.O (g21396), .I (g17955));
INVX1 gate8104(.O (g31616), .I (I29214));
INVX1 gate8105(.O (I14079), .I (g7231));
INVX1 gate8106(.O (g30063), .I (g29015));
INVX1 gate8107(.O (I22124), .I (g21300));
INVX1 gate8108(.O (g9771), .I (g3969));
INVX1 gate8109(.O (I29973), .I (g31213));
INVX1 gate8110(.O (g26834), .I (I25552));
INVX1 gate8111(.O (g20911), .I (g15171));
INVX1 gate8112(.O (I16028), .I (g12381));
INVX1 gate8113(.O (g10369), .I (g6873));
INVX1 gate8114(.O (g32744), .I (g31327));
INVX1 gate8115(.O (I31515), .I (g33187));
INVX1 gate8116(.O (g24911), .I (I24078));
INVX1 gate8117(.O (g19677), .I (g17096));
INVX1 gate8118(.O (I18280), .I (g12951));
INVX1 gate8119(.O (g12490), .I (I15316));
INVX1 gate8120(.O (g17512), .I (g12983));
INVX1 gate8121(.O (I17679), .I (g13416));
INVX1 gate8122(.O (g21413), .I (g15585));
INVX1 gate8123(.O (g9299), .I (g5124));
INVX1 gate8124(.O (I15788), .I (g10430));
INVX1 gate8125(.O (g23413), .I (g21012));
INVX1 gate8126(.O (g27956), .I (I26466));
INVX1 gate8127(.O (g32849), .I (g31021));
INVX1 gate8128(.O (g9547), .I (g2735));
INVX1 gate8129(.O (g10368), .I (g6887));
INVX1 gate8130(.O (g32940), .I (g31376));
INVX1 gate8131(.O (g7379), .I (g2299));
INVX1 gate8132(.O (g8400), .I (g4836));
INVX1 gate8133(.O (g11724), .I (I14593));
INVX1 gate8134(.O (I17188), .I (g13782));
INVX1 gate8135(.O (g31809), .I (g29385));
INVX1 gate8136(.O (I12487), .I (g3443));
INVX1 gate8137(.O (g11325), .I (g7543));
INVX1 gate8138(.O (g20071), .I (g16826));
INVX1 gate8139(.O (g32848), .I (g30825));
INVX1 gate8140(.O (g9892), .I (g6428));
INVX1 gate8141(.O (g24071), .I (g20841));
INVX1 gate8142(.O (g11829), .I (I14653));
INVX1 gate8143(.O (g12889), .I (g10396));
INVX1 gate8144(.O (g11920), .I (I14730));
INVX1 gate8145(.O (I11632), .I (g16));
INVX1 gate8146(.O (g20591), .I (g15509));
INVX1 gate8147(.O (g25781), .I (g24510));
INVX1 gate8148(.O (g10412), .I (g7072));
INVX1 gate8149(.O (g20776), .I (g18008));
INVX1 gate8150(.O (g20785), .I (I20846));
INVX1 gate8151(.O (g31808), .I (g29385));
INVX1 gate8152(.O (g32652), .I (g30735));
INVX1 gate8153(.O (g32804), .I (g30735));
INVX1 gate8154(.O (g14412), .I (I16564));
INVX1 gate8155(.O (g7289), .I (g4382));
INVX1 gate8156(.O (I12618), .I (g3338));
INVX1 gate8157(.O (g12888), .I (g10395));
INVX1 gate8158(.O (g26614), .I (g25426));
INVX1 gate8159(.O (g10133), .I (g6049));
INVX1 gate8160(.O (g20147), .I (g17328));
INVX1 gate8161(.O (I17938), .I (g3676));
INVX1 gate8162(.O (g34209), .I (I32170));
INVX1 gate8163(.O (g7835), .I (g4125));
INVX1 gate8164(.O (g24147), .I (g19402));
INVX1 gate8165(.O (g10229), .I (g6736));
INVX1 gate8166(.O (I18066), .I (g3317));
INVX1 gate8167(.O (g12181), .I (g9478));
INVX1 gate8168(.O (g26607), .I (g25382));
INVX1 gate8169(.O (g17499), .I (g14885));
INVX1 gate8170(.O (g22989), .I (g20453));
INVX1 gate8171(.O (g23929), .I (g19147));
INVX1 gate8172(.O (g17316), .I (I18293));
INVX1 gate8173(.O (g11344), .I (g9015));
INVX1 gate8174(.O (g34208), .I (g33838));
INVX1 gate8175(.O (I14158), .I (g8806));
INVX1 gate8176(.O (g19410), .I (g16449));
INVX1 gate8177(.O (g24825), .I (g23204));
INVX1 gate8178(.O (g22722), .I (I22031));
INVX1 gate8179(.O (g17498), .I (g14688));
INVX1 gate8180(.O (g22988), .I (g20391));
INVX1 gate8181(.O (g8183), .I (g482));
INVX1 gate8182(.O (g23020), .I (g19869));
INVX1 gate8183(.O (I15682), .I (g12182));
INVX1 gate8184(.O (g23928), .I (g21562));
INVX1 gate8185(.O (g8608), .I (g278));
INVX1 gate8186(.O (I18885), .I (g16643));
INVX1 gate8187(.O (g30021), .I (g28994));
INVX1 gate8188(.O (I32071), .I (g33665));
INVX1 gate8189(.O (g19479), .I (g16449));
INVX1 gate8190(.O (g19666), .I (g17188));
INVX1 gate8191(.O (g6782), .I (I11632));
INVX1 gate8192(.O (g25264), .I (g23828));
INVX1 gate8193(.O (g16692), .I (g14170));
INVX1 gate8194(.O (g25790), .I (g25027));
INVX1 gate8195(.O (I29013), .I (g29705));
INVX1 gate8196(.O (g25137), .I (g22432));
INVX1 gate8197(.O (g9340), .I (I13094));
INVX1 gate8198(.O (I13715), .I (g71));
INVX1 gate8199(.O (g17056), .I (g13437));
INVX1 gate8200(.O (I29214), .I (g30300));
INVX1 gate8201(.O (g11291), .I (g7526));
INVX1 gate8202(.O (I32591), .I (g34287));
INVX1 gate8203(.O (g24172), .I (I23360));
INVX1 gate8204(.O (g23046), .I (g20283));
INVX1 gate8205(.O (g32962), .I (g30735));
INVX1 gate8206(.O (g9478), .I (I13152));
INVX1 gate8207(.O (I14823), .I (g8056));
INVX1 gate8208(.O (g19478), .I (g16000));
INVX1 gate8209(.O (g24996), .I (g22763));
INVX1 gate8210(.O (g17611), .I (g14822));
INVX1 gate8211(.O (g17722), .I (I18709));
INVX1 gate8212(.O (g9907), .I (g1959));
INVX1 gate8213(.O (g13173), .I (g10632));
INVX1 gate8214(.O (g34913), .I (I33131));
INVX1 gate8215(.O (g10582), .I (g7116));
INVX1 gate8216(.O (I16755), .I (g12377));
INVX1 gate8217(.O (I29207), .I (g30293));
INVX1 gate8218(.O (g14582), .I (I16698));
INVX1 gate8219(.O (g33874), .I (I31724));
INVX1 gate8220(.O (g9959), .I (g6177));
INVX1 gate8221(.O (g7674), .I (I12151));
INVX1 gate8222(.O (g8977), .I (g4349));
INVX1 gate8223(.O (g24367), .I (g22550));
INVX1 gate8224(.O (g24394), .I (g22228));
INVX1 gate8225(.O (I16770), .I (g6023));
INVX1 gate8226(.O (g32500), .I (g30735));
INVX1 gate8227(.O (g34436), .I (I32479));
INVX1 gate8228(.O (g9517), .I (g6163));
INVX1 gate8229(.O (g9690), .I (g732));
INVX1 gate8230(.O (g17432), .I (I18379));
INVX1 gate8231(.O (g23787), .I (g18997));
INVX1 gate8232(.O (I27677), .I (g28156));
INVX1 gate8233(.O (g29170), .I (g27907));
INVX1 gate8234(.O (g32833), .I (g30825));
INVX1 gate8235(.O (g18957), .I (I19734));
INVX1 gate8236(.O (g21282), .I (I21019));
INVX1 gate8237(.O (g16214), .I (g13437));
INVX1 gate8238(.O (g17271), .I (I18270));
INVX1 gate8239(.O (I32950), .I (g34713));
INVX1 gate8240(.O (g23282), .I (g20330));
INVX1 gate8241(.O (I26710), .I (g27511));
INVX1 gate8242(.O (g7541), .I (g344));
INVX1 gate8243(.O (g10627), .I (I13968));
INVX1 gate8244(.O (I25105), .I (g25284));
INVX1 gate8245(.O (g34320), .I (g34119));
INVX1 gate8246(.O (g27089), .I (g26703));
INVX1 gate8247(.O (g10379), .I (g6953));
INVX1 gate8248(.O (g23302), .I (g20330));
INVX1 gate8249(.O (I25743), .I (g25903));
INVX1 gate8250(.O (g31665), .I (I29245));
INVX1 gate8251(.O (g25209), .I (g22763));
INVX1 gate8252(.O (g19580), .I (g16164));
INVX1 gate8253(.O (g30593), .I (g29970));
INVX1 gate8254(.O (g33665), .I (I31500));
INVX1 gate8255(.O (g6998), .I (g4932));
INVX1 gate8256(.O (g22199), .I (g19210));
INVX1 gate8257(.O (g34530), .I (I32591));
INVX1 gate8258(.O (g10112), .I (g1988));
INVX1 gate8259(.O (g34593), .I (I32687));
INVX1 gate8260(.O (g7132), .I (g4558));
INVX1 gate8261(.O (g12546), .I (g8740));
INVX1 gate8262(.O (I22470), .I (g21326));
INVX1 gate8263(.O (g10050), .I (g6336));
INVX1 gate8264(.O (g27088), .I (g26694));
INVX1 gate8265(.O (g18562), .I (I19384));
INVX1 gate8266(.O (g34346), .I (g34162));
INVX1 gate8267(.O (g10378), .I (g6926));
INVX1 gate8268(.O (g25208), .I (g22763));
INVX1 gate8269(.O (g30565), .I (I28832));
INVX1 gate8270(.O (g7153), .I (g5373));
INVX1 gate8271(.O (g7680), .I (g4108));
INVX1 gate8272(.O (g8451), .I (g4057));
INVX1 gate8273(.O (g22198), .I (g19147));
INVX1 gate8274(.O (g22529), .I (g19549));
INVX1 gate8275(.O (g34122), .I (I32059));
INVX1 gate8276(.O (g15799), .I (g13110));
INVX1 gate8277(.O (I21831), .I (g19127));
INVX1 gate8278(.O (g13506), .I (g10808));
INVX1 gate8279(.O (g12088), .I (g7701));
INVX1 gate8280(.O (g13028), .I (I15650));
INVX1 gate8281(.O (g20446), .I (g15224));
INVX1 gate8282(.O (g10386), .I (g6982));
INVX1 gate8283(.O (g29194), .I (I27492));
INVX1 gate8284(.O (g9915), .I (g2583));
INVX1 gate8285(.O (g12860), .I (g10368));
INVX1 gate8286(.O (g22528), .I (g19801));
INVX1 gate8287(.O (g6850), .I (g2704));
INVX1 gate8288(.O (g14386), .I (I16544));
INVX1 gate8289(.O (g23769), .I (g19074));
INVX1 gate8290(.O (I11980), .I (g66));
INVX1 gate8291(.O (g22330), .I (g19801));
INVX1 gate8292(.O (I13889), .I (g7598));
INVX1 gate8293(.O (g25542), .I (g22763));
INVX1 gate8294(.O (g7802), .I (g324));
INVX1 gate8295(.O (g20059), .I (g17302));
INVX1 gate8296(.O (g32613), .I (g30673));
INVX1 gate8297(.O (g8146), .I (g1760));
INVX1 gate8298(.O (g10096), .I (g5767));
INVX1 gate8299(.O (g20025), .I (g17271));
INVX1 gate8300(.O (g8346), .I (g3845));
INVX1 gate8301(.O (g24059), .I (g21193));
INVX1 gate8302(.O (g33454), .I (I30980));
INVX1 gate8303(.O (g14096), .I (I16328));
INVX1 gate8304(.O (g24025), .I (g21256));
INVX1 gate8305(.O (g9214), .I (g617));
INVX1 gate8306(.O (g17529), .I (g15039));
INVX1 gate8307(.O (g20540), .I (g16646));
INVX1 gate8308(.O (g12497), .I (g9780));
INVX1 gate8309(.O (g30292), .I (g28736));
INVX1 gate8310(.O (I16898), .I (g10615));
INVX1 gate8311(.O (g23768), .I (g18997));
INVX1 gate8312(.O (I12884), .I (g4213));
INVX1 gate8313(.O (I22467), .I (g19662));
INVX1 gate8314(.O (g20058), .I (g16782));
INVX1 gate8315(.O (g24540), .I (g22942));
INVX1 gate8316(.O (g33712), .I (I31561));
INVX1 gate8317(.O (I26356), .I (g26843));
INVX1 gate8318(.O (I18307), .I (g12977));
INVX1 gate8319(.O (g32947), .I (g31376));
INVX1 gate8320(.O (g19531), .I (g16816));
INVX1 gate8321(.O (g24058), .I (g20982));
INVX1 gate8322(.O (g22869), .I (g20875));
INVX1 gate8323(.O (g17528), .I (g14940));
INVX1 gate8324(.O (g7558), .I (I12041));
INVX1 gate8325(.O (g32605), .I (g30614));
INVX1 gate8326(.O (g8696), .I (g3347));
INVX1 gate8327(.O (g34409), .I (g34145));
INVX1 gate8328(.O (I21722), .I (g19264));
INVX1 gate8329(.O (g22868), .I (g20453));
INVX1 gate8330(.O (I16521), .I (g10430));
INVX1 gate8331(.O (g17764), .I (I18758));
INVX1 gate8332(.O (I12666), .I (g4040));
INVX1 gate8333(.O (g10429), .I (g7148));
INVX1 gate8334(.O (g11927), .I (g10207));
INVX1 gate8335(.O (g23881), .I (g19277));
INVX1 gate8336(.O (g10857), .I (g8712));
INVX1 gate8337(.O (g32812), .I (g30825));
INVX1 gate8338(.O (g25073), .I (I24237));
INVX1 gate8339(.O (g32463), .I (g31566));
INVX1 gate8340(.O (g16100), .I (I17471));
INVX1 gate8341(.O (I32446), .I (g34127));
INVX1 gate8342(.O (g19676), .I (g17062));
INVX1 gate8343(.O (g19685), .I (g16987));
INVX1 gate8344(.O (g31239), .I (g29916));
INVX1 gate8345(.O (g25274), .I (g22763));
INVX1 gate8346(.O (g24044), .I (g21127));
INVX1 gate8347(.O (g16771), .I (g14018));
INVX1 gate8348(.O (g34408), .I (g34144));
INVX1 gate8349(.O (I22419), .I (g19638));
INVX1 gate8350(.O (g19373), .I (g16449));
INVX1 gate8351(.O (g26575), .I (g25268));
INVX1 gate8352(.O (g10428), .I (g9631));
INVX1 gate8353(.O (g32951), .I (g31021));
INVX1 gate8354(.O (g32972), .I (g31710));
INVX1 gate8355(.O (g16235), .I (g13437));
INVX1 gate8356(.O (g32033), .I (g30929));
INVX1 gate8357(.O (I32059), .I (g33648));
INVX1 gate8358(.O (g8508), .I (g3827));
INVX1 gate8359(.O (g19654), .I (g16931));
INVX1 gate8360(.O (I31361), .I (g33120));
INVX1 gate8361(.O (g9402), .I (g6209));
INVX1 gate8362(.O (g9824), .I (g1825));
INVX1 gate8363(.O (g8944), .I (g370));
INVX1 gate8364(.O (g8240), .I (g1333));
INVX1 gate8365(.O (g18661), .I (I19487));
INVX1 gate8366(.O (g20902), .I (I20870));
INVX1 gate8367(.O (g18895), .I (g16000));
INVX1 gate8368(.O (g19800), .I (g17096));
INVX1 gate8369(.O (I18341), .I (g14308));
INVX1 gate8370(.O (g19417), .I (g17178));
INVX1 gate8371(.O (g21662), .I (g16540));
INVX1 gate8372(.O (g24377), .I (g22594));
INVX1 gate8373(.O (g7092), .I (g6483));
INVX1 gate8374(.O (I31500), .I (g33176));
INVX1 gate8375(.O (g24120), .I (g19984));
INVX1 gate8376(.O (g23027), .I (g20391));
INVX1 gate8377(.O (g32795), .I (g31327));
INVX1 gate8378(.O (g25034), .I (g23695));
INVX1 gate8379(.O (I23342), .I (g23299));
INVX1 gate8380(.O (g17709), .I (g14761));
INVX1 gate8381(.O (g33382), .I (g32033));
INVX1 gate8382(.O (I12580), .I (g1239));
INVX1 gate8383(.O (g8443), .I (g3736));
INVX1 gate8384(.O (g19334), .I (I19818));
INVX1 gate8385(.O (g20146), .I (g17533));
INVX1 gate8386(.O (g20738), .I (g15483));
INVX1 gate8387(.O (I18180), .I (g13605));
INVX1 gate8388(.O (g25641), .I (I24784));
INVX1 gate8389(.O (g20562), .I (g17955));
INVX1 gate8390(.O (g9590), .I (g1882));
INVX1 gate8391(.O (g21249), .I (g15509));
INVX1 gate8392(.O (I15981), .I (g11290));
INVX1 gate8393(.O (g24146), .I (g19422));
INVX1 gate8394(.O (g6986), .I (g4743));
INVX1 gate8395(.O (g23249), .I (g21070));
INVX1 gate8396(.O (I14687), .I (g7753));
INVX1 gate8397(.O (g11770), .I (I14619));
INVX1 gate8398(.O (I21199), .I (g17501));
INVX1 gate8399(.O (I30998), .I (g32453));
INVX1 gate8400(.O (g20699), .I (g17873));
INVX1 gate8401(.O (g16515), .I (g13486));
INVX1 gate8402(.O (g10504), .I (g8763));
INVX1 gate8403(.O (g11981), .I (I14823));
INVX1 gate8404(.O (g9657), .I (g2763));
INVX1 gate8405(.O (g12968), .I (g11793));
INVX1 gate8406(.O (g17471), .I (g14454));
INVX1 gate8407(.O (g25153), .I (g23733));
INVX1 gate8408(.O (I26448), .I (g26860));
INVX1 gate8409(.O (g8316), .I (g2351));
INVX1 gate8410(.O (g17087), .I (g14321));
INVX1 gate8411(.O (g23482), .I (g18833));
INVX1 gate8412(.O (I25552), .I (g25240));
INVX1 gate8413(.O (g32514), .I (g30735));
INVX1 gate8414(.O (I18734), .I (g6373));
INVX1 gate8415(.O (g24699), .I (g23047));
INVX1 gate8416(.O (g21248), .I (g15224));
INVX1 gate8417(.O (g14504), .I (g12361));
INVX1 gate8418(.O (g19762), .I (g16326));
INVX1 gate8419(.O (g23248), .I (g20924));
INVX1 gate8420(.O (g19964), .I (g17200));
INVX1 gate8421(.O (I22589), .I (g21340));
INVX1 gate8422(.O (g20698), .I (g17873));
INVX1 gate8423(.O (g27527), .I (I26195));
INVX1 gate8424(.O (g25409), .I (g22228));
INVX1 gate8425(.O (g34575), .I (I32651));
INVX1 gate8426(.O (I25779), .I (g26424));
INVX1 gate8427(.O (g32507), .I (g30735));
INVX1 gate8428(.O (g9556), .I (g5448));
INVX1 gate8429(.O (I18839), .I (g13716));
INVX1 gate8430(.O (g23003), .I (I22180));
INVX1 gate8431(.O (g8565), .I (g3802));
INVX1 gate8432(.O (g21204), .I (g15656));
INVX1 gate8433(.O (g33637), .I (I31466));
INVX1 gate8434(.O (g29177), .I (g27937));
INVX1 gate8435(.O (g30327), .I (I28582));
INVX1 gate8436(.O (g33935), .I (I31817));
INVX1 gate8437(.O (g34711), .I (g34559));
INVX1 gate8438(.O (g12870), .I (g10374));
INVX1 gate8439(.O (I11860), .I (g43));
INVX1 gate8440(.O (g25136), .I (g22457));
INVX1 gate8441(.O (g34327), .I (g34108));
INVX1 gate8442(.O (I18667), .I (g6661));
INVX1 gate8443(.O (I18694), .I (g5666));
INVX1 gate8444(.O (g32421), .I (g31213));
INVX1 gate8445(.O (I23330), .I (g22658));
INVX1 gate8446(.O (I23393), .I (g23414));
INVX1 gate8447(.O (g10129), .I (g5352));
INVX1 gate8448(.O (I29441), .I (g30917));
INVX1 gate8449(.O (g11845), .I (I14663));
INVX1 gate8450(.O (g9064), .I (g4983));
INVX1 gate8451(.O (I18131), .I (g13350));
INVX1 gate8452(.O (g8681), .I (g763));
INVX1 gate8453(.O (g10002), .I (g6195));
INVX1 gate8454(.O (I25786), .I (g26424));
INVX1 gate8455(.O (g10057), .I (g6455));
INVX1 gate8456(.O (g9899), .I (g6513));
INVX1 gate8457(.O (I32645), .I (g34367));
INVX1 gate8458(.O (g7262), .I (g5723));
INVX1 gate8459(.O (g24366), .I (g22594));
INVX1 gate8460(.O (g20632), .I (g15171));
INVX1 gate8461(.O (I15633), .I (g12074));
INVX1 gate8462(.O (I32699), .I (g34569));
INVX1 gate8463(.O (I33273), .I (g34984));
INVX1 gate8464(.O (g30606), .I (I28866));
INVX1 gate8465(.O (g8697), .I (g3694));
INVX1 gate8466(.O (I33106), .I (g34855));
INVX1 gate8467(.O (I14668), .I (g7753));
INVX1 gate8468(.O (I25356), .I (g24374));
INVX1 gate8469(.O (g19543), .I (g16349));
INVX1 gate8470(.O (g30303), .I (g28786));
INVX1 gate8471(.O (g8914), .I (g4264));
INVX1 gate8472(.O (I19796), .I (g17870));
INVX1 gate8473(.O (g17602), .I (g14962));
INVX1 gate8474(.O (g12867), .I (g10375));
INVX1 gate8475(.O (g12894), .I (g10401));
INVX1 gate8476(.O (I17401), .I (g13394));
INVX1 gate8477(.O (g16584), .I (g13920));
INVX1 gate8478(.O (g17774), .I (g14902));
INVX1 gate8479(.O (g23647), .I (g18833));
INVX1 gate8480(.O (g18889), .I (g15509));
INVX1 gate8481(.O (g17955), .I (I18865));
INVX1 gate8482(.O (g18980), .I (g16136));
INVX1 gate8483(.O (g32541), .I (g30673));
INVX1 gate8484(.O (g7623), .I (I12103));
INVX1 gate8485(.O (g10323), .I (I13744));
INVX1 gate8486(.O (g23945), .I (g21611));
INVX1 gate8487(.O (g16206), .I (g13437));
INVX1 gate8488(.O (I25380), .I (g24481));
INVX1 gate8489(.O (g18095), .I (I18891));
INVX1 gate8490(.O (g23356), .I (g21070));
INVX1 gate8491(.O (g32473), .I (g31070));
INVX1 gate8492(.O (I31463), .I (g33318));
INVX1 gate8493(.O (g19908), .I (g16540));
INVX1 gate8494(.O (g22171), .I (g18882));
INVX1 gate8495(.O (g13191), .I (I15788));
INVX1 gate8496(.O (g26840), .I (I25562));
INVX1 gate8497(.O (g20661), .I (g15171));
INVX1 gate8498(.O (I12654), .I (g1585));
INVX1 gate8499(.O (g21380), .I (g17955));
INVX1 gate8500(.O (g10533), .I (g8795));
INVX1 gate8501(.O (g20547), .I (g15224));
INVX1 gate8502(.O (g23999), .I (g21468));
INVX1 gate8503(.O (g32789), .I (g30735));
INVX1 gate8504(.O (g18888), .I (g15426));
INVX1 gate8505(.O (g23380), .I (g20619));
INVX1 gate8506(.O (g33729), .I (I31586));
INVX1 gate8507(.O (I18443), .I (g13027));
INVX1 gate8508(.O (g19569), .I (g16349));
INVX1 gate8509(.O (I14424), .I (g4005));
INVX1 gate8510(.O (I14016), .I (g9104));
INVX1 gate8511(.O (I17118), .I (g14363));
INVX1 gate8512(.O (g16725), .I (g13963));
INVX1 gate8513(.O (I22748), .I (g19458));
INVX1 gate8514(.O (g13521), .I (g11357));
INVX1 gate8515(.O (g22994), .I (g20436));
INVX1 gate8516(.O (g34982), .I (I33246));
INVX1 gate8517(.O (g32788), .I (g31327));
INVX1 gate8518(.O (g32724), .I (g30735));
INVX1 gate8519(.O (g19747), .I (g17015));
INVX1 gate8520(.O (g23233), .I (g21037));
INVX1 gate8521(.O (g21182), .I (g15509));
INVX1 gate8522(.O (g6789), .I (I11635));
INVX1 gate8523(.O (g11832), .I (g8011));
INVX1 gate8524(.O (g23182), .I (g21389));
INVX1 gate8525(.O (g20715), .I (g15277));
INVX1 gate8526(.O (g23651), .I (g20655));
INVX1 gate8527(.O (g32829), .I (g30937));
INVX1 gate8528(.O (g28080), .I (I26581));
INVX1 gate8529(.O (g32920), .I (g30825));
INVX1 gate8530(.O (I18469), .I (g13809));
INVX1 gate8531(.O (g32535), .I (g31554));
INVX1 gate8532(.O (g25327), .I (g22161));
INVX1 gate8533(.O (g32434), .I (g31189));
INVX1 gate8534(.O (I14830), .I (g10141));
INVX1 gate8535(.O (I21258), .I (g16540));
INVX1 gate8536(.O (g24481), .I (I23684));
INVX1 gate8537(.O (I14893), .I (g9819));
INVX1 gate8538(.O (g25109), .I (g23666));
INVX1 gate8539(.O (g12818), .I (g8792));
INVX1 gate8540(.O (g20551), .I (g17302));
INVX1 gate8541(.O (g20572), .I (g15833));
INVX1 gate8542(.O (g9194), .I (g827));
INVX1 gate8543(.O (g32828), .I (g31710));
INVX1 gate8544(.O (g18931), .I (g16031));
INVX1 gate8545(.O (g6987), .I (g4754));
INVX1 gate8546(.O (g32946), .I (g31327));
INVX1 gate8547(.O (g10232), .I (g4527));
INVX1 gate8548(.O (I17276), .I (g13605));
INVX1 gate8549(.O (g7285), .I (g4643));
INVX1 gate8550(.O (g11861), .I (g8070));
INVX1 gate8551(.O (g22919), .I (g21163));
INVX1 gate8552(.O (g16744), .I (I17964));
INVX1 gate8553(.O (I17704), .I (g13144));
INVX1 gate8554(.O (g12978), .I (I15593));
INVX1 gate8555(.O (g14232), .I (g11083));
INVX1 gate8556(.O (g9731), .I (g5366));
INVX1 gate8557(.O (g23331), .I (g20905));
INVX1 gate8558(.O (I13968), .I (g7697));
INVX1 gate8559(.O (I32547), .I (g34397));
INVX1 gate8560(.O (g19751), .I (g16044));
INVX1 gate8561(.O (I24839), .I (g24298));
INVX1 gate8562(.O (g9489), .I (g2303));
INVX1 gate8563(.O (g19772), .I (g17183));
INVX1 gate8564(.O (g25283), .I (g22763));
INVX1 gate8565(.O (g34840), .I (I33056));
INVX1 gate8566(.O (g20127), .I (I20388));
INVX1 gate8567(.O (I22177), .I (g21366));
INVX1 gate8568(.O (g23449), .I (g18833));
INVX1 gate8569(.O (g26483), .I (I25359));
INVX1 gate8570(.O (g28753), .I (I27235));
INVX1 gate8571(.O (g9557), .I (g5499));
INVX1 gate8572(.O (g13926), .I (I16217));
INVX1 gate8573(.O (g24127), .I (g19984));
INVX1 gate8574(.O (g13045), .I (g11941));
INVX1 gate8575(.O (g10261), .I (g4555));
INVX1 gate8576(.O (I17808), .I (g13311));
INVX1 gate8577(.O (g9071), .I (g2831));
INVX1 gate8578(.O (g26862), .I (I25598));
INVX1 gate8579(.O (g11388), .I (I14395));
INVX1 gate8580(.O (g23897), .I (g19210));
INVX1 gate8581(.O (g13099), .I (I15732));
INVX1 gate8582(.O (g11324), .I (g7542));
INVX1 gate8583(.O (g23448), .I (g21611));
INVX1 gate8584(.O (g23961), .I (g19074));
INVX1 gate8585(.O (g32682), .I (g30825));
INVX1 gate8586(.O (g24490), .I (g22594));
INVX1 gate8587(.O (I14705), .I (g7717));
INVX1 gate8588(.O (g19638), .I (g17324));
INVX1 gate8589(.O (I17101), .I (g14338));
INVX1 gate8590(.O (g34192), .I (g33921));
INVX1 gate8591(.O (I21810), .I (g20596));
INVX1 gate8592(.O (I16629), .I (g11987));
INVX1 gate8593(.O (g16652), .I (g13892));
INVX1 gate8594(.O (g17010), .I (I18138));
INVX1 gate8595(.O (g23505), .I (g21514));
INVX1 gate8596(.O (I27543), .I (g28187));
INVX1 gate8597(.O (g26326), .I (g24872));
INVX1 gate8598(.O (g8922), .I (I12907));
INVX1 gate8599(.O (g20385), .I (g18008));
INVX1 gate8600(.O (I14679), .I (g9332));
INVX1 gate8601(.O (g13251), .I (I15814));
INVX1 gate8602(.O (I23375), .I (g23403));
INVX1 gate8603(.O (g13272), .I (I15837));
INVX1 gate8604(.O (g19416), .I (g15885));
INVX1 gate8605(.O (g20103), .I (g17433));
INVX1 gate8606(.O (g7424), .I (g2465));
INVX1 gate8607(.O (g24376), .I (g22722));
INVX1 gate8608(.O (g24385), .I (g22908));
INVX1 gate8609(.O (g34522), .I (g34271));
INVX1 gate8610(.O (g7809), .I (g4864));
INVX1 gate8611(.O (I18143), .I (g13350));
INVX1 gate8612(.O (g24103), .I (g21209));
INVX1 gate8613(.O (g23026), .I (g20391));
INVX1 gate8614(.O (g18088), .I (g13267));
INVX1 gate8615(.O (g24980), .I (g22384));
INVX1 gate8616(.O (I16246), .I (g3983));
INVX1 gate8617(.O (I30971), .I (g32015));
INVX1 gate8618(.O (I12117), .I (g586));
INVX1 gate8619(.O (g24095), .I (g21209));
INVX1 gate8620(.O (g26702), .I (g25309));
INVX1 gate8621(.O (g17599), .I (g14794));
INVX1 gate8622(.O (I12000), .I (g582));
INVX1 gate8623(.O (g25174), .I (g23890));
INVX1 gate8624(.O (g28696), .I (g27858));
INVX1 gate8625(.O (g31653), .I (g29713));
INVX1 gate8626(.O (g6991), .I (g4888));
INVX1 gate8627(.O (g33653), .I (I31486));
INVX1 gate8628(.O (I14939), .I (g10216));
INVX1 gate8629(.O (g7231), .I (g5));
INVX1 gate8630(.O (g20671), .I (g15509));
INVX1 gate8631(.O (I17733), .I (g14844));
INVX1 gate8632(.O (g27018), .I (I25750));
INVX1 gate8633(.O (g31138), .I (g29778));
INVX1 gate8634(.O (g32760), .I (g30735));
INVX1 gate8635(.O (g17086), .I (g14297));
INVX1 gate8636(.O (g24181), .I (I23387));
INVX1 gate8637(.O (g7523), .I (g305));
INVX1 gate8638(.O (g19579), .I (g16000));
INVX1 gate8639(.O (g22159), .I (I21744));
INVX1 gate8640(.O (g29941), .I (g28900));
INVX1 gate8641(.O (g13140), .I (g10632));
INVX1 gate8642(.O (g7643), .I (g4322));
INVX1 gate8643(.O (I21792), .I (g21308));
INVX1 gate8644(.O (I12568), .I (g5005));
INVX1 gate8645(.O (g12018), .I (g9538));
INVX1 gate8646(.O (I22009), .I (g21269));
INVX1 gate8647(.O (g34553), .I (I32621));
INVX1 gate8648(.O (g10499), .I (I13872));
INVX1 gate8649(.O (I22665), .I (g21308));
INVX1 gate8650(.O (I13581), .I (g6727));
INVX1 gate8651(.O (I18168), .I (g13191));
INVX1 gate8652(.O (I24278), .I (g23440));
INVX1 gate8653(.O (I14267), .I (g7835));
INVX1 gate8654(.O (g32506), .I (g31376));
INVX1 gate8655(.O (g8784), .I (I12764));
INVX1 gate8656(.O (I31724), .I (g33076));
INVX1 gate8657(.O (g33636), .I (I31463));
INVX1 gate8658(.O (g29185), .I (I27481));
INVX1 gate8659(.O (I32956), .I (g34654));
INVX1 gate8660(.O (g30326), .I (I28579));
INVX1 gate8661(.O (g21723), .I (I21288));
INVX1 gate8662(.O (g29092), .I (g27800));
INVX1 gate8663(.O (I32297), .I (g34059));
INVX1 gate8664(.O (g34949), .I (g34939));
INVX1 gate8665(.O (g10498), .I (g7161));
INVX1 gate8666(.O (I32103), .I (g33661));
INVX1 gate8667(.O (g34326), .I (g34091));
INVX1 gate8668(.O (g13061), .I (g10981));
INVX1 gate8669(.O (I31829), .I (g33454));
INVX1 gate8670(.O (I18479), .I (g13041));
INVX1 gate8671(.O (g31852), .I (g29385));
INVX1 gate8672(.O (g6959), .I (g4420));
INVX1 gate8673(.O (I31535), .I (g33377));
INVX1 gate8674(.O (g30040), .I (g29025));
INVX1 gate8675(.O (I13202), .I (g5105));
INVX1 gate8676(.O (g19586), .I (g16349));
INVX1 gate8677(.O (I12123), .I (g758));
INVX1 gate8678(.O (g17125), .I (I18177));
INVX1 gate8679(.O (g17532), .I (I18479));
INVX1 gate8680(.O (g27402), .I (I26100));
INVX1 gate8681(.O (g34536), .I (I32601));
INVX1 gate8682(.O (I17166), .I (g14536));
INVX1 gate8683(.O (g28161), .I (I26676));
INVX1 gate8684(.O (g7634), .I (I12123));
INVX1 gate8685(.O (g15758), .I (I17276));
INVX1 gate8686(.O (g21387), .I (I21115));
INVX1 gate8687(.O (I22485), .I (g21308));
INVX1 gate8688(.O (I29221), .I (g30307));
INVX1 gate8689(.O (g23433), .I (g21562));
INVX1 gate8690(.O (I28419), .I (g29195));
INVX1 gate8691(.O (I13979), .I (g7733));
INVX1 gate8692(.O (I32824), .I (g34475));
INVX1 gate8693(.O (g24426), .I (g22722));
INVX1 gate8694(.O (g8479), .I (g3057));
INVX1 gate8695(.O (g20190), .I (g16971));
INVX1 gate8696(.O (g22144), .I (g18997));
INVX1 gate8697(.O (I24038), .I (g22202));
INVX1 gate8698(.O (g23620), .I (I22769));
INVX1 gate8699(.O (g28709), .I (I27192));
INVX1 gate8700(.O (g10080), .I (g1982));
INVX1 gate8701(.O (I17008), .I (g12857));
INVX1 gate8702(.O (I32671), .I (g34388));
INVX1 gate8703(.O (g8840), .I (g4277));
INVX1 gate8704(.O (g9212), .I (g6466));
INVX1 gate8705(.O (g12866), .I (g10369));
INVX1 gate8706(.O (I21918), .I (g21290));
INVX1 gate8707(.O (I17892), .I (g3325));
INVX1 gate8708(.O (g21343), .I (g16428));
INVX1 gate8709(.O (I26925), .I (g27015));
INVX1 gate8710(.O (g8390), .I (g3385));
INVX1 gate8711(.O (g32927), .I (g30825));
INVX1 gate8712(.O (g15345), .I (I17108));
INVX1 gate8713(.O (g14432), .I (g12311));
INVX1 gate8714(.O (g17680), .I (g14889));
INVX1 gate8715(.O (g17144), .I (g14085));
INVX1 gate8716(.O (g26634), .I (g25317));
INVX1 gate8717(.O (g26851), .I (I25579));
INVX1 gate8718(.O (g11447), .I (I14450));
INVX1 gate8719(.O (g7926), .I (g3423));
INVX1 gate8720(.O (I15162), .I (g10176));
INVX1 gate8721(.O (g20546), .I (g18008));
INVX1 gate8722(.O (g20089), .I (g17533));
INVX1 gate8723(.O (g23971), .I (g20751));
INVX1 gate8724(.O (I26378), .I (g26850));
INVX1 gate8725(.O (g19720), .I (I20130));
INVX1 gate8726(.O (g20211), .I (g16931));
INVX1 gate8727(.O (I25369), .I (g24891));
INVX1 gate8728(.O (g24089), .I (g19890));
INVX1 gate8729(.O (I19851), .I (g16615));
INVX1 gate8730(.O (g27597), .I (g26745));
INVX1 gate8731(.O (g21369), .I (g16285));
INVX1 gate8732(.O (I33291), .I (g34983));
INVX1 gate8733(.O (g12077), .I (I14939));
INVX1 gate8734(.O (g32649), .I (g30673));
INVX1 gate8735(.O (g25553), .I (g22550));
INVX1 gate8736(.O (g20088), .I (g17533));
INVX1 gate8737(.O (I27391), .I (g27929));
INVX1 gate8738(.O (g8356), .I (g54));
INVX1 gate8739(.O (I20937), .I (g16967));
INVX1 gate8740(.O (g9229), .I (g5052));
INVX1 gate8741(.O (I13094), .I (g2724));
INVX1 gate8742(.O (g14753), .I (g11317));
INVX1 gate8743(.O (I33173), .I (g34887));
INVX1 gate8744(.O (g24088), .I (g21209));
INVX1 gate8745(.O (g19493), .I (g16349));
INVX1 gate8746(.O (g24024), .I (g21193));
INVX1 gate8747(.O (g14342), .I (g12163));
INVX1 gate8748(.O (g34673), .I (I32803));
INVX1 gate8749(.O (g34847), .I (I33067));
INVX1 gate8750(.O (g31609), .I (I29211));
INVX1 gate8751(.O (g29215), .I (I27561));
INVX1 gate8752(.O (g10031), .I (I13552));
INVX1 gate8753(.O (g32648), .I (g30614));
INVX1 gate8754(.O (g32491), .I (g31566));
INVX1 gate8755(.O (g32903), .I (g31376));
INVX1 gate8756(.O (g25326), .I (g22228));
INVX1 gate8757(.O (g14031), .I (I16289));
INVX1 gate8758(.O (g9822), .I (g125));
INVX1 gate8759(.O (g10199), .I (g1968));
INVX1 gate8760(.O (I11801), .I (g6395));
INVX1 gate8761(.O (I14455), .I (g10197));
INVX1 gate8762(.O (g16605), .I (g13955));
INVX1 gate8763(.O (g11472), .I (g7918));
INVX1 gate8764(.O (I27579), .I (g28184));
INVX1 gate8765(.O (I29371), .I (g30325));
INVX1 gate8766(.O (g12923), .I (I15542));
INVX1 gate8767(.O (g31608), .I (g29653));
INVX1 gate8768(.O (g18527), .I (I19345));
INVX1 gate8769(.O (g20497), .I (g18065));
INVX1 gate8770(.O (g32604), .I (g31154));
INVX1 gate8771(.O (g34062), .I (g33711));
INVX1 gate8772(.O (I28588), .I (g29368));
INVX1 gate8773(.O (g32755), .I (g31672));
INVX1 gate8774(.O (I30959), .I (g32021));
INVX1 gate8775(.O (g10198), .I (I13672));
INVX1 gate8776(.O (g12300), .I (I15144));
INVX1 gate8777(.O (g11911), .I (g10022));
INVX1 gate8778(.O (g16812), .I (g13555));
INVX1 gate8779(.O (g21412), .I (g15758));
INVX1 gate8780(.O (g32770), .I (g31710));
INVX1 gate8781(.O (g34933), .I (g34916));
INVX1 gate8782(.O (g14198), .I (g12180));
INVX1 gate8783(.O (g32563), .I (g31554));
INVX1 gate8784(.O (I32089), .I (g33665));
INVX1 gate8785(.O (I33134), .I (g34906));
INVX1 gate8786(.O (g13246), .I (g10939));
INVX1 gate8787(.O (g20700), .I (g17873));
INVX1 gate8788(.O (g20659), .I (g17873));
INVX1 gate8789(.O (g34851), .I (I33075));
INVX1 gate8790(.O (g20625), .I (g15348));
INVX1 gate8791(.O (g10393), .I (g6991));
INVX1 gate8792(.O (g24126), .I (g19935));
INVX1 gate8793(.O (g24625), .I (g23135));
INVX1 gate8794(.O (g14330), .I (I16486));
INVX1 gate8795(.O (g24987), .I (g23630));
INVX1 gate8796(.O (g8954), .I (g1079));
INVX1 gate8797(.O (g7543), .I (I12033));
INVX1 gate8798(.O (g31799), .I (g29385));
INVX1 gate8799(.O (g23896), .I (g19210));
INVX1 gate8800(.O (g25564), .I (g22312));
INVX1 gate8801(.O (g8363), .I (g239));
INVX1 gate8802(.O (g18894), .I (g16000));
INVX1 gate8803(.O (g31813), .I (g29385));
INVX1 gate8804(.O (g21228), .I (g17531));
INVX1 gate8805(.O (g33799), .I (g33299));
INVX1 gate8806(.O (g10365), .I (g6867));
INVX1 gate8807(.O (g22224), .I (g19277));
INVX1 gate8808(.O (g33813), .I (I31659));
INVX1 gate8809(.O (g8032), .I (I12355));
INVX1 gate8810(.O (g19517), .I (g16777));
INVX1 gate8811(.O (g23228), .I (g21070));
INVX1 gate8812(.O (I18373), .I (g13011));
INVX1 gate8813(.O (g29906), .I (g28793));
INVX1 gate8814(.O (g29348), .I (g28194));
INVX1 gate8815(.O (g16795), .I (I18009));
INVX1 gate8816(.O (g10960), .I (g9007));
INVX1 gate8817(.O (I17675), .I (g13394));
INVX1 gate8818(.O (g23011), .I (g20330));
INVX1 gate8819(.O (g31798), .I (g29385));
INVX1 gate8820(.O (g32767), .I (g30735));
INVX1 gate8821(.O (g32794), .I (g30937));
INVX1 gate8822(.O (I14623), .I (g8925));
INVX1 gate8823(.O (g11147), .I (g8417));
INVX1 gate8824(.O (g11754), .I (g8229));
INVX1 gate8825(.O (I17154), .I (g13605));
INVX1 gate8826(.O (I23680), .I (g23219));
INVX1 gate8827(.O (g25183), .I (g22763));
INVX1 gate8828(.O (g32899), .I (g31021));
INVX1 gate8829(.O (g7534), .I (g1367));
INVX1 gate8830(.O (g31805), .I (g29385));
INVX1 gate8831(.O (g17224), .I (I18248));
INVX1 gate8832(.O (g16514), .I (g14139));
INVX1 gate8833(.O (g12885), .I (g10382));
INVX1 gate8834(.O (g22495), .I (g19801));
INVX1 gate8835(.O (g17308), .I (g14876));
INVX1 gate8836(.O (g23582), .I (I22729));
INVX1 gate8837(.O (g32633), .I (g31154));
INVX1 gate8838(.O (g32898), .I (g30825));
INVX1 gate8839(.O (I32659), .I (g34391));
INVX1 gate8840(.O (g15048), .I (I16969));
INVX1 gate8841(.O (g9620), .I (g6187));
INVX1 gate8842(.O (g9462), .I (g6215));
INVX1 gate8843(.O (I23336), .I (g22721));
INVX1 gate8844(.O (I19756), .I (g17812));
INVX1 gate8845(.O (g19362), .I (g16072));
INVX1 gate8846(.O (g7927), .I (g4064));
INVX1 gate8847(.O (g34574), .I (I32648));
INVX1 gate8848(.O (g32719), .I (g31672));
INVX1 gate8849(.O (I12041), .I (g2741));
INVX1 gate8850(.O (g20060), .I (g16540));
INVX1 gate8851(.O (g34047), .I (g33637));
INVX1 gate8852(.O (g18979), .I (g16136));
INVX1 gate8853(.O (g19523), .I (g16100));
INVX1 gate8854(.O (g24060), .I (g21256));
INVX1 gate8855(.O (g8912), .I (g4180));
INVX1 gate8856(.O (I16120), .I (g11868));
INVX1 gate8857(.O (g33934), .I (I31814));
INVX1 gate8858(.O (g10708), .I (g7836));
INVX1 gate8859(.O (g20197), .I (g16987));
INVX1 gate8860(.O (g6928), .I (I11716));
INVX1 gate8861(.O (I12746), .I (g4087));
INVX1 gate8862(.O (g21379), .I (g17873));
INVX1 gate8863(.O (g34311), .I (g34097));
INVX1 gate8864(.O (I12493), .I (g5002));
INVX1 gate8865(.O (g22976), .I (I22149));
INVX1 gate8866(.O (g22985), .I (g20330));
INVX1 gate8867(.O (g32718), .I (g30825));
INVX1 gate8868(.O (g32521), .I (g31376));
INVX1 gate8869(.O (g10087), .I (I13597));
INVX1 gate8870(.O (g23925), .I (g21514));
INVX1 gate8871(.O (g8357), .I (I12538));
INVX1 gate8872(.O (g18978), .I (g16000));
INVX1 gate8873(.O (g7946), .I (I12314));
INVX1 gate8874(.O (g7660), .I (I12144));
INVX1 gate8875(.O (g29653), .I (I27927));
INVX1 gate8876(.O (I22729), .I (g21308));
INVX1 gate8877(.O (g26820), .I (I25534));
INVX1 gate8878(.O (g21050), .I (g17873));
INVX1 gate8879(.O (g20527), .I (g18008));
INVX1 gate8880(.O (I13597), .I (g4417));
INVX1 gate8881(.O (g11367), .I (I14381));
INVX1 gate8882(.O (g28918), .I (g27832));
INVX1 gate8883(.O (g32832), .I (g30735));
INVX1 gate8884(.O (I20321), .I (g16920));
INVX1 gate8885(.O (g23378), .I (g21070));
INVX1 gate8886(.O (g13394), .I (I15915));
INVX1 gate8887(.O (I31491), .I (g33283));
INVX1 gate8888(.O (g33761), .I (I31616));
INVX1 gate8889(.O (g24527), .I (g22670));
INVX1 gate8890(.O (g7903), .I (g969));
INVX1 gate8891(.O (g30072), .I (I28301));
INVX1 gate8892(.O (g17687), .I (g15042));
INVX1 gate8893(.O (I31604), .I (g33176));
INVX1 gate8894(.O (g28079), .I (I26578));
INVX1 gate8895(.O (g10043), .I (g1632));
INVX1 gate8896(.O (I13280), .I (g6140));
INVX1 gate8897(.O (g7513), .I (g6315));
INVX1 gate8898(.O (g26731), .I (g25470));
INVX1 gate8899(.O (g34592), .I (I32684));
INVX1 gate8900(.O (I11688), .I (g70));
INVX1 gate8901(.O (I16698), .I (g12077));
INVX1 gate8902(.O (g29333), .I (g28167));
INVX1 gate8903(.O (g16473), .I (g13977));
INVX1 gate8904(.O (I31770), .I (g33197));
INVX1 gate8905(.O (g32861), .I (g31376));
INVX1 gate8906(.O (g9842), .I (g3274));
INVX1 gate8907(.O (g23944), .I (g19147));
INVX1 gate8908(.O (g32573), .I (g30825));
INVX1 gate8909(.O (g18094), .I (I18888));
INVX1 gate8910(.O (g31013), .I (g29679));
INVX1 gate8911(.O (I14589), .I (g8818));
INVX1 gate8912(.O (g25213), .I (g23293));
INVX1 gate8913(.O (g19437), .I (g16349));
INVX1 gate8914(.O (g20503), .I (g15373));
INVX1 gate8915(.O (g9298), .I (g5080));
INVX1 gate8916(.O (g28598), .I (g27717));
INVX1 gate8917(.O (I18909), .I (g16873));
INVX1 gate8918(.O (g9392), .I (g5869));
INVX1 gate8919(.O (g32926), .I (g31376));
INVX1 gate8920(.O (I32855), .I (g34540));
INVX1 gate8921(.O (g7178), .I (g4392));
INVX1 gate8922(.O (g7436), .I (g5276));
INVX1 gate8923(.O (I14836), .I (g9688));
INVX1 gate8924(.O (g8626), .I (g4040));
INVX1 gate8925(.O (g21681), .I (I21242));
INVX1 gate8926(.O (g29963), .I (g28931));
INVX1 gate8927(.O (g16724), .I (g14079));
INVX1 gate8928(.O (g22842), .I (g19875));
INVX1 gate8929(.O (g23681), .I (g21012));
INVX1 gate8930(.O (I18117), .I (g13302));
INVX1 gate8931(.O (g32612), .I (g30614));
INVX1 gate8932(.O (g16325), .I (g13223));
INVX1 gate8933(.O (g18877), .I (g15224));
INVX1 gate8934(.O (I23309), .I (g21677));
INVX1 gate8935(.O (g25452), .I (g22228));
INVX1 gate8936(.O (g15371), .I (I17114));
INVX1 gate8937(.O (g25047), .I (g23733));
INVX1 gate8938(.O (g32099), .I (g31009));
INVX1 gate8939(.O (g10375), .I (g6941));
INVX1 gate8940(.O (I21288), .I (g18216));
INVX1 gate8941(.O (g34820), .I (I33034));
INVX1 gate8942(.O (g16920), .I (I18086));
INVX1 gate8943(.O (g20714), .I (g15277));
INVX1 gate8944(.O (g20450), .I (g15277));
INVX1 gate8945(.O (g23429), .I (g20453));
INVX1 gate8946(.O (g32701), .I (g31376));
INVX1 gate8947(.O (g12076), .I (g9280));
INVX1 gate8948(.O (g7335), .I (g2287));
INVX1 gate8949(.O (g7831), .I (I12227));
INVX1 gate8950(.O (I14119), .I (g7824));
INVX1 gate8951(.O (g32777), .I (g31710));
INVX1 gate8952(.O (g32534), .I (g30673));
INVX1 gate8953(.O (g12721), .I (g10061));
INVX1 gate8954(.O (g34152), .I (I32109));
INVX1 gate8955(.O (g20707), .I (g18008));
INVX1 gate8956(.O (g21428), .I (g15758));
INVX1 gate8957(.O (I22622), .I (g21209));
INVX1 gate8958(.O (g20910), .I (g15171));
INVX1 gate8959(.O (g34846), .I (I33064));
INVX1 gate8960(.O (g23793), .I (g19074));
INVX1 gate8961(.O (g12054), .I (g7690));
INVX1 gate8962(.O (g17392), .I (g14924));
INVX1 gate8963(.O (g19600), .I (g16164));
INVX1 gate8964(.O (g10337), .I (g5016));
INVX1 gate8965(.O (g24819), .I (I23998));
INVX1 gate8966(.O (g19781), .I (g16489));
INVX1 gate8967(.O (g17489), .I (g12955));
INVX1 gate8968(.O (I24334), .I (g22976));
INVX1 gate8969(.O (g20496), .I (g17929));
INVX1 gate8970(.O (g7805), .I (g4366));
INVX1 gate8971(.O (g7916), .I (I12300));
INVX1 gate8972(.O (g25051), .I (I24215));
INVX1 gate8973(.O (g25072), .I (g23630));
INVX1 gate8974(.O (g24818), .I (g23191));
INVX1 gate8975(.O (g32462), .I (g30673));
INVX1 gate8976(.O (I14749), .I (g10031));
INVX1 gate8977(.O (g24979), .I (g22369));
INVX1 gate8978(.O (g21690), .I (g16540));
INVX1 gate8979(.O (g22830), .I (g20283));
INVX1 gate8980(.O (g19952), .I (g15915));
INVX1 gate8981(.O (g24055), .I (g19968));
INVX1 gate8982(.O (g7749), .I (g996));
INVX1 gate8983(.O (g19351), .I (g17367));
INVX1 gate8984(.O (I12523), .I (g3794));
INVX1 gate8985(.O (g23549), .I (g18833));
INVX1 gate8986(.O (g27773), .I (I26378));
INVX1 gate8987(.O (g20070), .I (g16173));
INVX1 gate8988(.O (g20978), .I (g15595));
INVX1 gate8989(.O (g24111), .I (g19890));
INVX1 gate8990(.O (g28656), .I (g27742));
INVX1 gate8991(.O (g9708), .I (g2741));
INVX1 gate8992(.O (g24070), .I (g20014));
INVX1 gate8993(.O (g24978), .I (g22342));
INVX1 gate8994(.O (g34691), .I (I32843));
INVX1 gate8995(.O (g29312), .I (g28877));
INVX1 gate8996(.O (g20590), .I (g15426));
INVX1 gate8997(.O (g22544), .I (g19589));
INVX1 gate8998(.O (g22865), .I (g20330));
INVX1 gate8999(.O (g23548), .I (g18833));
INVX1 gate9000(.O (g8778), .I (I12758));
INVX1 gate9001(.O (g29115), .I (g27779));
INVX1 gate9002(.O (g7947), .I (g1500));
INVX1 gate9003(.O (I20216), .I (g15862));
INVX1 gate9004(.O (g24986), .I (g23590));
INVX1 gate9005(.O (I14305), .I (g8805));
INVX1 gate9006(.O (g9252), .I (g4304));
INVX1 gate9007(.O (I26880), .I (g27527));
INVX1 gate9008(.O (g23504), .I (g21468));
INVX1 gate9009(.O (g13902), .I (g11389));
INVX1 gate9010(.O (g13301), .I (g10862));
INVX1 gate9011(.O (g31771), .I (I29337));
INVX1 gate9012(.O (g19264), .I (I19802));
INVX1 gate9013(.O (g18917), .I (g16077));
INVX1 gate9014(.O (g19790), .I (g16971));
INVX1 gate9015(.O (g20384), .I (g18008));
INVX1 gate9016(.O (g12180), .I (g9477));
INVX1 gate9017(.O (g9958), .I (g6148));
INVX1 gate9018(.O (g29921), .I (g28864));
INVX1 gate9019(.O (g13120), .I (g10632));
INVX1 gate9020(.O (I18293), .I (g1079));
INVX1 gate9021(.O (g24384), .I (g22885));
INVX1 gate9022(.O (g25820), .I (g25051));
INVX1 gate9023(.O (I26512), .I (g26817));
INVX1 gate9024(.O (I17653), .I (g14276));
INVX1 gate9025(.O (g20067), .I (g17328));
INVX1 gate9026(.O (g32766), .I (g31376));
INVX1 gate9027(.O (g6955), .I (I11726));
INVX1 gate9028(.O (g29745), .I (g28500));
INVX1 gate9029(.O (g24067), .I (g21256));
INVX1 gate9030(.O (g24094), .I (g21143));
INVX1 gate9031(.O (g11562), .I (g7648));
INVX1 gate9032(.O (g17713), .I (g12947));
INVX1 gate9033(.O (I18265), .I (g13350));
INVX1 gate9034(.O (g34929), .I (I33179));
INVX1 gate9035(.O (g27930), .I (I26451));
INVX1 gate9036(.O (I12437), .I (g4999));
INVX1 gate9037(.O (g27993), .I (I26503));
INVX1 gate9038(.O (g8075), .I (g3742));
INVX1 gate9039(.O (g32871), .I (g30937));
INVX1 gate9040(.O (g30020), .I (g29097));
INVX1 gate9041(.O (g30928), .I (I28908));
INVX1 gate9042(.O (g22189), .I (I21769));
INVX1 gate9043(.O (g8475), .I (I12608));
INVX1 gate9044(.O (g26105), .I (I25146));
INVX1 gate9045(.O (g9829), .I (g2250));
INVX1 gate9046(.O (g12839), .I (g10350));
INVX1 gate9047(.O (g6814), .I (g632));
INVX1 gate9048(.O (g12930), .I (g12347));
INVX1 gate9049(.O (g7873), .I (g1266));
INVX1 gate9050(.O (g26743), .I (g25476));
INVX1 gate9051(.O (g26827), .I (g24819));
INVX1 gate9052(.O (g34583), .I (I32665));
INVX1 gate9053(.O (g7632), .I (I12117));
INVX1 gate9054(.O (g34928), .I (I33176));
INVX1 gate9055(.O (g7095), .I (g6545));
INVX1 gate9056(.O (I17636), .I (g14252));
INVX1 gate9057(.O (g21057), .I (g15426));
INVX1 gate9058(.O (g23002), .I (I22177));
INVX1 gate9059(.O (g10079), .I (g1950));
INVX1 gate9060(.O (g11290), .I (I14326));
INVX1 gate9061(.O (g24150), .I (g19268));
INVX1 gate9062(.O (g23057), .I (g20453));
INVX1 gate9063(.O (I28594), .I (g29379));
INVX1 gate9064(.O (g9911), .I (g2384));
INVX1 gate9065(.O (g7495), .I (g4375));
INVX1 gate9066(.O (g14545), .I (g12768));
INVX1 gate9067(.O (g7437), .I (g5666));
INVX1 gate9068(.O (g17610), .I (g15008));
INVX1 gate9069(.O (I27253), .I (g27996));
INVX1 gate9070(.O (I30995), .I (g32449));
INVX1 gate9071(.O (g12838), .I (g10353));
INVX1 gate9072(.O (g23128), .I (g20283));
INVX1 gate9073(.O (I20569), .I (g16486));
INVX1 gate9074(.O (I17852), .I (g3625));
INVX1 gate9075(.O (g10078), .I (g1854));
INVX1 gate9076(.O (g21245), .I (I20982));
INVX1 gate9077(.O (g24019), .I (g19968));
INVX1 gate9078(.O (g17189), .I (g14708));
INVX1 gate9079(.O (g23245), .I (g20785));
INVX1 gate9080(.O (I13287), .I (g110));
INVX1 gate9081(.O (g26769), .I (g25400));
INVX1 gate9082(.O (g8526), .I (g1526));
INVX1 gate9083(.O (g19208), .I (g17367));
INVX1 gate9084(.O (g20695), .I (I20781));
INVX1 gate9085(.O (I20747), .I (g17141));
INVX1 gate9086(.O (I31701), .I (g33164));
INVX1 gate9087(.O (g21299), .I (g16600));
INVX1 gate9088(.O (g30113), .I (g29154));
INVX1 gate9089(.O (g9733), .I (g5736));
INVX1 gate9090(.O (g10086), .I (g2193));
INVX1 gate9091(.O (g23323), .I (g20283));
INVX1 gate9092(.O (g23299), .I (I22400));
INVX1 gate9093(.O (g9974), .I (g2518));
INVX1 gate9094(.O (I32067), .I (g33661));
INVX1 gate9095(.O (g17188), .I (I18224));
INVX1 gate9096(.O (I11721), .I (g4145));
INVX1 gate9097(.O (g17124), .I (g14051));
INVX1 gate9098(.O (g17678), .I (I18653));
INVX1 gate9099(.O (g34787), .I (I32991));
INVX1 gate9100(.O (g26803), .I (g25389));
INVX1 gate9101(.O (g12487), .I (g9340));
INVX1 gate9102(.O (g20526), .I (g15171));
INVX1 gate9103(.O (I22576), .I (g21282));
INVX1 gate9104(.O (I28185), .I (g28803));
INVX1 gate9105(.O (I18835), .I (g6365));
INVX1 gate9106(.O (I13054), .I (g6744));
INVX1 gate9107(.O (g24526), .I (g22942));
INVX1 gate9108(.O (g19542), .I (g16349));
INVX1 gate9109(.O (g30302), .I (g28924));
INVX1 gate9110(.O (g7752), .I (g1542));
INVX1 gate9111(.O (I16181), .I (g3672));
INVX1 gate9112(.O (g18102), .I (I18912));
INVX1 gate9113(.O (g8439), .I (g3129));
INVX1 gate9114(.O (g9073), .I (g150));
INVX1 gate9115(.O (g32629), .I (g31376));
INVX1 gate9116(.O (g34302), .I (I32305));
INVX1 gate9117(.O (I26989), .I (g27277));
INVX1 gate9118(.O (I32150), .I (g33923));
INVX1 gate9119(.O (g30105), .I (I28336));
INVX1 gate9120(.O (g6836), .I (g1322));
INVX1 gate9121(.O (g7917), .I (g1157));
INVX1 gate9122(.O (I14630), .I (g7717));
INVX1 gate9123(.O (g27279), .I (g26330));
INVX1 gate9124(.O (g32472), .I (g30825));
INVX1 gate9125(.O (g10159), .I (g4477));
INVX1 gate9126(.O (g34827), .I (I33041));
INVX1 gate9127(.O (g10532), .I (g10233));
INVX1 gate9128(.O (g32628), .I (g31542));
INVX1 gate9129(.O (g17093), .I (I18165));
INVX1 gate9130(.O (g6918), .I (g3639));
INVX1 gate9131(.O (g32911), .I (g31376));
INVX1 gate9132(.O (g14125), .I (I16345));
INVX1 gate9133(.O (g15344), .I (g14851));
INVX1 gate9134(.O (g10158), .I (g2461));
INVX1 gate9135(.O (g11403), .I (g7595));
INVX1 gate9136(.O (g11547), .I (I14505));
INVX1 gate9137(.O (g13895), .I (I16193));
INVX1 gate9138(.O (g20917), .I (g15224));
INVX1 gate9139(.O (I33140), .I (g34884));
INVX1 gate9140(.O (I28883), .I (g30105));
INVX1 gate9141(.O (g23232), .I (I22331));
INVX1 gate9142(.O (g24866), .I (I24038));
INVX1 gate9143(.O (g19905), .I (g15885));
INVX1 gate9144(.O (I12790), .I (g4340));
INVX1 gate9145(.O (I17609), .I (g13510));
INVX1 gate9146(.O (g34769), .I (I32953));
INVX1 gate9147(.O (I11655), .I (g1246));
INVX1 gate9148(.O (g18876), .I (g15373));
INVX1 gate9149(.O (g18885), .I (g15979));
INVX1 gate9150(.O (g10353), .I (g6803));
INVX1 gate9151(.O (g25046), .I (g23729));
INVX1 gate9152(.O (g6993), .I (g4859));
INVX1 gate9153(.O (g10295), .I (I13723));
INVX1 gate9154(.O (g8919), .I (I12896));
INVX1 gate9155(.O (g21697), .I (I21258));
INVX1 gate9156(.O (g29013), .I (I27368));
INVX1 gate9157(.O (I29981), .I (g31591));
INVX1 gate9158(.O (g34768), .I (I32950));
INVX1 gate9159(.O (g12039), .I (I14899));
INVX1 gate9160(.O (g13715), .I (g10573));
INVX1 gate9161(.O (I22745), .I (g19458));
INVX1 gate9162(.O (g29214), .I (I27558));
INVX1 gate9163(.O (g27038), .I (g25932));
INVX1 gate9164(.O (g9206), .I (g5164));
INVX1 gate9165(.O (g32591), .I (g30614));
INVX1 gate9166(.O (I15572), .I (g10499));
INVX1 gate9167(.O (g23995), .I (g19277));
INVX1 gate9168(.O (g32776), .I (g31672));
INVX1 gate9169(.O (g32785), .I (g31710));
INVX1 gate9170(.O (I30989), .I (g32441));
INVX1 gate9171(.O (g19565), .I (g16000));
INVX1 gate9172(.O (g24077), .I (g20720));
INVX1 gate9173(.O (g20706), .I (g18008));
INVX1 gate9174(.O (I11734), .I (g4473));
INVX1 gate9175(.O (g23880), .I (g19210));
INVX1 gate9176(.O (g12038), .I (I14896));
INVX1 gate9177(.O (g20597), .I (g17847));
INVX1 gate9178(.O (I21042), .I (g15824));
INVX1 gate9179(.O (g32754), .I (g30825));
INVX1 gate9180(.O (I14570), .I (g7932));
INVX1 gate9181(.O (g33435), .I (I30959));
INVX1 gate9182(.O (g25282), .I (g22763));
INVX1 gate9183(.O (I21189), .I (g17475));
INVX1 gate9184(.O (g14336), .I (I16498));
INVX1 gate9185(.O (g27187), .I (I25882));
INVX1 gate9186(.O (g7296), .I (g5313));
INVX1 gate9187(.O (g23512), .I (g20248));
INVX1 gate9188(.O (g8616), .I (g2803));
INVX1 gate9189(.O (g28752), .I (I27232));
INVX1 gate9190(.O (g20923), .I (g15277));
INVX1 gate9191(.O (g27975), .I (g26694));
INVX1 gate9192(.O (g32859), .I (g30614));
INVX1 gate9193(.O (g32825), .I (g30735));
INVX1 gate9194(.O (g32950), .I (g31672));
INVX1 gate9195(.O (g28954), .I (g27830));
INVX1 gate9196(.O (g26710), .I (g25349));
INVX1 gate9197(.O (g18660), .I (I19484));
INVX1 gate9198(.O (g20624), .I (g18065));
INVX1 gate9199(.O (g22455), .I (g19801));
INVX1 gate9200(.O (g12975), .I (g12752));
INVX1 gate9201(.O (g7532), .I (g1157));
INVX1 gate9202(.O (I13694), .I (g117));
INVX1 gate9203(.O (I16024), .I (g11171));
INVX1 gate9204(.O (g32858), .I (g31327));
INVX1 gate9205(.O (g33744), .I (I31604));
INVX1 gate9206(.O (g7553), .I (g1274));
INVX1 gate9207(.O (g8404), .I (g5005));
INVX1 gate9208(.O (g15506), .I (I17131));
INVX1 gate9209(.O (g31849), .I (g29385));
INVX1 gate9210(.O (g8647), .I (g3416));
INVX1 gate9211(.O (g14631), .I (g12239));
INVX1 gate9212(.O (g10364), .I (g6869));
INVX1 gate9213(.O (g19409), .I (g16431));
INVX1 gate9214(.O (I14567), .I (g9708));
INVX1 gate9215(.O (g12143), .I (I14999));
INVX1 gate9216(.O (g20102), .I (g17533));
INVX1 gate9217(.O (g16767), .I (I17989));
INVX1 gate9218(.O (g20157), .I (g16886));
INVX1 gate9219(.O (g25640), .I (I24781));
INVX1 gate9220(.O (g12937), .I (g12419));
INVX1 gate9221(.O (g28669), .I (g27705));
INVX1 gate9222(.O (g26081), .I (g24619));
INVX1 gate9223(.O (g8764), .I (g4826));
INVX1 gate9224(.O (g22201), .I (g19277));
INVX1 gate9225(.O (g24102), .I (g21143));
INVX1 gate9226(.O (g23445), .I (I22564));
INVX1 gate9227(.O (g31848), .I (g29385));
INVX1 gate9228(.O (g18916), .I (g16053));
INVX1 gate9229(.O (g24157), .I (I23315));
INVX1 gate9230(.O (g32844), .I (g30937));
INVX1 gate9231(.O (g9898), .I (g6444));
AN2X1 gate9232(.O (g33848), .I1 (g33261), .I2 (g20384));
AN2X1 gate9233(.O (g28260), .I1 (g27703), .I2 (g26518));
AN2X1 gate9234(.O (g17617), .I1 (g7885), .I2 (g13326));
AN2X1 gate9235(.O (g18550), .I1 (g2819), .I2 (g15277));
AN2X1 gate9236(.O (g25768), .I1 (g2912), .I2 (g24560));
AN2X1 gate9237(.O (g25803), .I1 (g24798), .I2 (g21024));
AN2X1 gate9238(.O (g31141), .I1 (g12224), .I2 (g30038));
AN3X1 gate9239(.O (I26960), .I1 (g24995), .I2 (g26424), .I3 (g22698));
AN2X1 gate9240(.O (g22075), .I1 (g6247), .I2 (g19210));
AN2X1 gate9241(.O (g18314), .I1 (g1585), .I2 (g16931));
AN2X1 gate9242(.O (g33652), .I1 (g33393), .I2 (g18889));
AN2X1 gate9243(.O (g18287), .I1 (g1442), .I2 (g16449));
AN2X1 gate9244(.O (g27410), .I1 (g26549), .I2 (g17527));
AN2X1 gate9245(.O (g16633), .I1 (g5196), .I2 (g14921));
AN2X1 gate9246(.O (g30248), .I1 (g28743), .I2 (g23938));
AN2X1 gate9247(.O (g34482), .I1 (g34405), .I2 (g18917));
AN2X1 gate9248(.O (g23498), .I1 (g20234), .I2 (g12998));
AN2X1 gate9249(.O (g28489), .I1 (g27010), .I2 (g12417));
AN2X1 gate9250(.O (g26356), .I1 (g15581), .I2 (g25523));
AN2X1 gate9251(.O (g18307), .I1 (g1559), .I2 (g16931));
AN2X1 gate9252(.O (g29771), .I1 (g28322), .I2 (g23242));
AN2X1 gate9253(.O (g30003), .I1 (g28149), .I2 (g9021));
AN2X1 gate9254(.O (g34710), .I1 (g34553), .I2 (g20903));
AN2X1 gate9255(.O (g16191), .I1 (g5475), .I2 (g14262));
AN2X1 gate9256(.O (g22623), .I1 (g19337), .I2 (g19470));
AN2X1 gate9257(.O (g21989), .I1 (g5587), .I2 (g19074));
AN2X1 gate9258(.O (g30204), .I1 (g28670), .I2 (g23868));
AN2X1 gate9259(.O (g13671), .I1 (g4498), .I2 (g10532));
AN2X1 gate9260(.O (g26826), .I1 (g24907), .I2 (g15747));
AN2X1 gate9261(.O (g27666), .I1 (g26865), .I2 (g23521));
AN4X1 gate9262(.O (I31246), .I1 (g31672), .I2 (g31839), .I3 (g32810), .I4 (g32811));
AN2X1 gate9263(.O (g18721), .I1 (g15138), .I2 (g16077));
AN2X1 gate9264(.O (g22037), .I1 (g5941), .I2 (g19147));
AN2X1 gate9265(.O (g25881), .I1 (g3821), .I2 (g24685));
AN2X1 gate9266(.O (g26380), .I1 (g19572), .I2 (g25547));
AN2X1 gate9267(.O (g33263), .I1 (g32393), .I2 (g25481));
AN2X1 gate9268(.O (g18596), .I1 (g2941), .I2 (g16349));
AN2X1 gate9269(.O (g32420), .I1 (g31127), .I2 (g19533));
AN2X1 gate9270(.O (g28488), .I1 (g27969), .I2 (g17713));
AN2X1 gate9271(.O (g27363), .I1 (g10231), .I2 (g26812));
AN2X1 gate9272(.O (g23056), .I1 (g16052), .I2 (g19860));
AN3X1 gate9273(.O (g27217), .I1 (g26236), .I2 (g8418), .I3 (g2610));
AN2X1 gate9274(.O (g29683), .I1 (g1821), .I2 (g29046));
AN2X1 gate9275(.O (g18243), .I1 (g1189), .I2 (g16431));
AN2X1 gate9276(.O (g33332), .I1 (g32217), .I2 (g20608));
AN3X1 gate9277(.O (I17692), .I1 (g14988), .I2 (g11450), .I3 (g6756));
AN2X1 gate9278(.O (g21988), .I1 (g5583), .I2 (g19074));
AN2X1 gate9279(.O (g26090), .I1 (g1624), .I2 (g25081));
AN2X1 gate9280(.O (g21924), .I1 (g5057), .I2 (g21468));
AN2X1 gate9281(.O (g28558), .I1 (g7301), .I2 (g27046));
AN2X1 gate9282(.O (g18431), .I1 (g2185), .I2 (g18008));
AN2X1 gate9283(.O (g26233), .I1 (g2279), .I2 (g25309));
AN4X1 gate9284(.O (I31071), .I1 (g31170), .I2 (g31808), .I3 (g32557), .I4 (g32558));
AN2X1 gate9285(.O (g26182), .I1 (g9978), .I2 (g25317));
AN2X1 gate9286(.O (g26651), .I1 (g22707), .I2 (g24425));
AN2X1 gate9287(.O (g12015), .I1 (g1002), .I2 (g7567));
AN2X1 gate9288(.O (g34081), .I1 (g33706), .I2 (g19552));
AN2X1 gate9289(.O (g27486), .I1 (g26519), .I2 (g17645));
AN2X1 gate9290(.O (g31962), .I1 (g8033), .I2 (g31013));
AN2X1 gate9291(.O (g24763), .I1 (g17569), .I2 (g22457));
AN2X1 gate9292(.O (g33406), .I1 (g32355), .I2 (g21399));
AN2X1 gate9293(.O (g18269), .I1 (g15069), .I2 (g16031));
AN2X1 gate9294(.O (g33361), .I1 (g32257), .I2 (g20911));
AN2X1 gate9295(.O (g15903), .I1 (g13796), .I2 (g13223));
AN2X1 gate9296(.O (g18773), .I1 (g5694), .I2 (g15615));
AN4X1 gate9297(.O (I31147), .I1 (g32668), .I2 (g32669), .I3 (g32670), .I4 (g32671));
AN2X1 gate9298(.O (g18341), .I1 (g1648), .I2 (g17873));
AN2X1 gate9299(.O (g29515), .I1 (g28888), .I2 (g22342));
AN2X1 gate9300(.O (g29882), .I1 (g2361), .I2 (g29151));
AN2X1 gate9301(.O (g18268), .I1 (g1280), .I2 (g16000));
AN2X1 gate9302(.O (g29991), .I1 (g29179), .I2 (g12922));
AN2X1 gate9303(.O (g21753), .I1 (g3179), .I2 (g20785));
AN2X1 gate9304(.O (g31500), .I1 (g29802), .I2 (g23449));
AN2X1 gate9305(.O (g18156), .I1 (g572), .I2 (g17533));
AN2X1 gate9306(.O (g18655), .I1 (g15106), .I2 (g14454));
AN3X1 gate9307(.O (g33500), .I1 (g32744), .I2 (I31196), .I3 (I31197));
AN2X1 gate9308(.O (g24660), .I1 (g22648), .I2 (g19737));
AN2X1 gate9309(.O (g33833), .I1 (g33093), .I2 (g25852));
AN2X1 gate9310(.O (g32203), .I1 (g4249), .I2 (g31327));
AN2X1 gate9311(.O (g18180), .I1 (g767), .I2 (g17328));
AN2X1 gate9312(.O (g26513), .I1 (g19501), .I2 (g24365));
AN2X1 gate9313(.O (g17418), .I1 (g9618), .I2 (g14407));
AN3X1 gate9314(.O (I27409), .I1 (g25556), .I2 (g26424), .I3 (g22698));
AN2X1 gate9315(.O (g34999), .I1 (g34998), .I2 (g23085));
AN2X1 gate9316(.O (g18670), .I1 (g4621), .I2 (g15758));
AN2X1 gate9317(.O (g34380), .I1 (g34158), .I2 (g20571));
AN3X1 gate9318(.O (g25482), .I1 (g5752), .I2 (g23816), .I3 (I24597));
AN2X1 gate9319(.O (g32044), .I1 (g31483), .I2 (g20085));
AN4X1 gate9320(.O (I24684), .I1 (g20014), .I2 (g24033), .I3 (g24034), .I4 (g24035));
AN2X1 gate9321(.O (g16612), .I1 (g5603), .I2 (g14927));
AN2X1 gate9322(.O (g21736), .I1 (g3065), .I2 (g20330));
AN2X1 gate9323(.O (g11546), .I1 (g7289), .I2 (g4375));
AN2X1 gate9324(.O (g21887), .I1 (g15101), .I2 (g19801));
AN2X1 gate9325(.O (g30233), .I1 (g28720), .I2 (g23913));
AN2X1 gate9326(.O (g18734), .I1 (g4966), .I2 (g16826));
AN4X1 gate9327(.O (I31151), .I1 (g30825), .I2 (g31822), .I3 (g32673), .I4 (g32674));
AN2X1 gate9328(.O (g16324), .I1 (g13657), .I2 (g182));
AN4X1 gate9329(.O (I31172), .I1 (g32703), .I2 (g32704), .I3 (g32705), .I4 (g32706));
AN2X1 gate9330(.O (g18335), .I1 (g1687), .I2 (g17873));
AN2X1 gate9331(.O (g16701), .I1 (g5547), .I2 (g14845));
AN2X1 gate9332(.O (g22589), .I1 (g19267), .I2 (g19451));
AN2X1 gate9333(.O (g32281), .I1 (g31257), .I2 (g20500));
AN2X1 gate9334(.O (g34182), .I1 (g33691), .I2 (g24384));
AN2X1 gate9335(.O (g28255), .I1 (g8515), .I2 (g27983));
AN2X1 gate9336(.O (g16534), .I1 (g5575), .I2 (g14665));
AN2X1 gate9337(.O (g28679), .I1 (g27572), .I2 (g20638));
AN2X1 gate9338(.O (g11024), .I1 (g5436), .I2 (g9070));
AN2X1 gate9339(.O (g16098), .I1 (g5148), .I2 (g14238));
AN3X1 gate9340(.O (I13937), .I1 (g7340), .I2 (g7293), .I3 (g7261));
AN2X1 gate9341(.O (g18993), .I1 (g11224), .I2 (g16172));
AN2X1 gate9342(.O (g24550), .I1 (g3684), .I2 (g23308));
AN2X1 gate9343(.O (g32301), .I1 (g31276), .I2 (g20547));
AN2X1 gate9344(.O (g14643), .I1 (g11998), .I2 (g12023));
AN2X1 gate9345(.O (g24314), .I1 (g4515), .I2 (g22228));
AN2X1 gate9346(.O (g22588), .I1 (g79), .I2 (g20078));
AN2X1 gate9347(.O (g21843), .I1 (g3869), .I2 (g21070));
AN2X1 gate9348(.O (g32120), .I1 (g31639), .I2 (g29941));
AN2X1 gate9349(.O (g24287), .I1 (g4401), .I2 (g22550));
AN2X1 gate9350(.O (g28124), .I1 (g27368), .I2 (g22842));
AN2X1 gate9351(.O (g15794), .I1 (g3239), .I2 (g14008));
AN2X1 gate9352(.O (g18667), .I1 (g4601), .I2 (g17367));
AN2X1 gate9353(.O (g18694), .I1 (g4722), .I2 (g16053));
AN2X1 gate9354(.O (g12179), .I1 (g9745), .I2 (g10027));
AN2X1 gate9355(.O (g24307), .I1 (g4486), .I2 (g22228));
AN2X1 gate9356(.O (g29584), .I1 (g1706), .I2 (g29018));
AN2X1 gate9357(.O (g27178), .I1 (g25997), .I2 (g16652));
AN2X1 gate9358(.O (g21764), .I1 (g3227), .I2 (g20785));
AN2X1 gate9359(.O (g11497), .I1 (g6398), .I2 (g7192));
AN2X1 gate9360(.O (g18131), .I1 (g482), .I2 (g16971));
AN3X1 gate9361(.O (g29206), .I1 (g24124), .I2 (I27528), .I3 (I27529));
AN2X1 gate9362(.O (g13497), .I1 (g2724), .I2 (g12155));
AN2X1 gate9363(.O (g28686), .I1 (g27574), .I2 (g20650));
AN2X1 gate9364(.O (g32146), .I1 (g31624), .I2 (g29978));
AN4X1 gate9365(.O (g28939), .I1 (g17321), .I2 (g25184), .I3 (g26424), .I4 (g27421));
AN2X1 gate9366(.O (g24721), .I1 (g17488), .I2 (g22369));
AN2X1 gate9367(.O (g22119), .I1 (g6581), .I2 (g19277));
AN2X1 gate9368(.O (g21869), .I1 (g4087), .I2 (g19801));
AN3X1 gate9369(.O (g27186), .I1 (g26195), .I2 (g8316), .I3 (g2342));
AN2X1 gate9370(.O (g31273), .I1 (g30143), .I2 (g27779));
AN2X1 gate9371(.O (g34513), .I1 (g9003), .I2 (g34346));
AN2X1 gate9372(.O (g21960), .I1 (g5421), .I2 (g21514));
AN2X1 gate9373(.O (g27676), .I1 (g26377), .I2 (g20627));
AN2X1 gate9374(.O (g27685), .I1 (g13032), .I2 (g25895));
AN2X1 gate9375(.O (g15633), .I1 (g3841), .I2 (g13584));
AN2X1 gate9376(.O (g33106), .I1 (g32408), .I2 (g18990));
AN2X1 gate9377(.O (g18487), .I1 (g2441), .I2 (g15426));
AN2X1 gate9378(.O (g27373), .I1 (g26488), .I2 (g17477));
AN2X1 gate9379(.O (g29759), .I1 (g28308), .I2 (g23226));
AN2X1 gate9380(.O (g22118), .I1 (g6605), .I2 (g19277));
AN2X1 gate9381(.O (g32290), .I1 (g31267), .I2 (g20525));
AN2X1 gate9382(.O (g11126), .I1 (g6035), .I2 (g10185));
AN2X1 gate9383(.O (g12186), .I1 (g1178), .I2 (g7519));
AN3X1 gate9384(.O (g28267), .I1 (g7328), .I2 (g2227), .I3 (g27421));
AN2X1 gate9385(.O (g17401), .I1 (g1083), .I2 (g13143));
AN2X1 gate9386(.O (g21868), .I1 (g4076), .I2 (g19801));
AN2X1 gate9387(.O (g18619), .I1 (g3466), .I2 (g17062));
AN2X1 gate9388(.O (g18502), .I1 (g2567), .I2 (g15509));
AN2X1 gate9389(.O (g22022), .I1 (g5873), .I2 (g19147));
AN2X1 gate9390(.O (g34961), .I1 (g34944), .I2 (g23019));
AN2X1 gate9391(.O (g12953), .I1 (g411), .I2 (g11048));
AN2X1 gate9392(.O (g18557), .I1 (g2771), .I2 (g15277));
AN3X1 gate9393(.O (g33812), .I1 (g23088), .I2 (g33187), .I3 (g9104));
AN2X1 gate9394(.O (g18210), .I1 (g936), .I2 (g15938));
AN2X1 gate9395(.O (g29758), .I1 (g28306), .I2 (g23222));
AN2X1 gate9396(.O (g17119), .I1 (g5272), .I2 (g14800));
AN3X1 gate9397(.O (g33463), .I1 (g32477), .I2 (I31011), .I3 (I31012));
AN4X1 gate9398(.O (I31227), .I1 (g32784), .I2 (g32785), .I3 (g32786), .I4 (g32787));
AN2X1 gate9399(.O (g18618), .I1 (g3457), .I2 (g17062));
AN2X1 gate9400(.O (g18443), .I1 (g2265), .I2 (g18008));
AN2X1 gate9401(.O (g24773), .I1 (g22832), .I2 (g19872));
AN2X1 gate9402(.O (g21709), .I1 (g283), .I2 (g20283));
AN2X1 gate9403(.O (g18279), .I1 (g1361), .I2 (g16136));
AN2X1 gate9404(.O (g30026), .I1 (g28476), .I2 (g25064));
AN2X1 gate9405(.O (g33371), .I1 (g32280), .I2 (g21155));
AN2X1 gate9406(.O (g30212), .I1 (g28687), .I2 (g23879));
AN2X1 gate9407(.O (g16766), .I1 (g6649), .I2 (g12915));
AN2X1 gate9408(.O (g26387), .I1 (g24813), .I2 (g20231));
AN2X1 gate9409(.O (g27334), .I1 (g12539), .I2 (g26769));
AN2X1 gate9410(.O (g34212), .I1 (g33761), .I2 (g22689));
AN2X1 gate9411(.O (g28219), .I1 (g9316), .I2 (g27573));
AN2X1 gate9412(.O (g21708), .I1 (g15049), .I2 (g20283));
AN2X1 gate9413(.O (g18278), .I1 (g1345), .I2 (g16136));
AN3X1 gate9414(.O (I16111), .I1 (g8691), .I2 (g11409), .I3 (g11381));
AN4X1 gate9415(.O (g26148), .I1 (g25357), .I2 (g11724), .I3 (g11709), .I4 (g11686));
AN2X1 gate9416(.O (g23708), .I1 (g19050), .I2 (g9104));
AN2X1 gate9417(.O (g16871), .I1 (g6597), .I2 (g14908));
AN2X1 gate9418(.O (g29345), .I1 (g4749), .I2 (g28376));
AN2X1 gate9419(.O (g22053), .I1 (g6116), .I2 (g21611));
AN2X1 gate9420(.O (g23471), .I1 (g20148), .I2 (g20523));
AN2X1 gate9421(.O (g26097), .I1 (g5821), .I2 (g25092));
AN2X1 gate9422(.O (g18469), .I1 (g2399), .I2 (g15224));
AN2X1 gate9423(.O (g24670), .I1 (g5138), .I2 (g23590));
AN2X1 gate9424(.O (g33795), .I1 (g33138), .I2 (g20782));
AN2X1 gate9425(.O (g28218), .I1 (g27768), .I2 (g26645));
AN2X1 gate9426(.O (g29940), .I1 (g1740), .I2 (g28758));
AN2X1 gate9427(.O (g26104), .I1 (g2250), .I2 (g25101));
AN2X1 gate9428(.O (g18286), .I1 (g1404), .I2 (g16164));
AN2X1 gate9429(.O (g22900), .I1 (g17137), .I2 (g19697));
AN4X1 gate9430(.O (g27762), .I1 (g22472), .I2 (g25226), .I3 (g26424), .I4 (g26218));
AN2X1 gate9431(.O (g15861), .I1 (g3957), .I2 (g14170));
AN2X1 gate9432(.O (g8690), .I1 (g2941), .I2 (g2936));
AN2X1 gate9433(.O (g27964), .I1 (g25956), .I2 (g22492));
AN2X1 gate9434(.O (g18468), .I1 (g2393), .I2 (g15224));
AN3X1 gate9435(.O (g25331), .I1 (g5366), .I2 (g22194), .I3 (I24508));
AN2X1 gate9436(.O (g18306), .I1 (g15074), .I2 (g16931));
AN2X1 gate9437(.O (g12762), .I1 (g4358), .I2 (g8977));
AN2X1 gate9438(.O (g22036), .I1 (g5937), .I2 (g19147));
AN2X1 gate9439(.O (g25449), .I1 (g6946), .I2 (g22496));
AN2X1 gate9440(.O (g13060), .I1 (g8587), .I2 (g11110));
AN2X1 gate9441(.O (g31514), .I1 (g20041), .I2 (g29956));
AN2X1 gate9442(.O (g32403), .I1 (g31117), .I2 (g15842));
AN2X1 gate9443(.O (g27216), .I1 (g26055), .I2 (g16725));
AN3X1 gate9444(.O (g33514), .I1 (g32844), .I2 (I31266), .I3 (I31267));
AN2X1 gate9445(.O (g22101), .I1 (g6474), .I2 (g18833));
AN2X1 gate9446(.O (g24930), .I1 (g4826), .I2 (g23948));
AN2X1 gate9447(.O (g29652), .I1 (g2667), .I2 (g29157));
AN2X1 gate9448(.O (g29804), .I1 (g1592), .I2 (g29014));
AN2X1 gate9449(.O (g17809), .I1 (g7873), .I2 (g13125));
AN4X1 gate9450(.O (I31281), .I1 (g30735), .I2 (g31845), .I3 (g32861), .I4 (g32862));
AN2X1 gate9451(.O (g28160), .I1 (g26309), .I2 (g27463));
AN2X1 gate9452(.O (g15612), .I1 (g3143), .I2 (g13530));
AN2X1 gate9453(.O (g25448), .I1 (g11202), .I2 (g22680));
AN2X1 gate9454(.O (g18815), .I1 (g6523), .I2 (g15483));
AN2X1 gate9455(.O (g30149), .I1 (g28605), .I2 (g21248));
AN2X1 gate9456(.O (g25961), .I1 (g25199), .I2 (g20682));
AN3X1 gate9457(.O (I27381), .I1 (g25549), .I2 (g26424), .I3 (g22698));
AN3X1 gate9458(.O (g33507), .I1 (g32795), .I2 (I31231), .I3 (I31232));
AN4X1 gate9459(.O (I31301), .I1 (g31327), .I2 (g31849), .I3 (g32889), .I4 (g32890));
AN2X1 gate9460(.O (g20131), .I1 (g15170), .I2 (g14309));
AN2X1 gate9461(.O (g15701), .I1 (g3821), .I2 (g13584));
AN3X1 gate9462(.O (g10705), .I1 (g6850), .I2 (g10219), .I3 (g2689));
AN2X1 gate9463(.O (g18601), .I1 (g3106), .I2 (g16987));
AN2X1 gate9464(.O (g13411), .I1 (g4955), .I2 (g11834));
AN2X1 gate9465(.O (g18187), .I1 (g794), .I2 (g17328));
AN2X1 gate9466(.O (g18677), .I1 (g4639), .I2 (g15758));
AN2X1 gate9467(.O (g14610), .I1 (g1484), .I2 (g10935));
AN2X1 gate9468(.O (g28455), .I1 (g27289), .I2 (g20103));
AN2X1 gate9469(.O (g33421), .I1 (g32374), .I2 (g21455));
AN2X1 gate9470(.O (g21810), .I1 (g3578), .I2 (g20924));
AN2X1 gate9471(.O (g17177), .I1 (g6657), .I2 (g14984));
AN2X1 gate9472(.O (g21774), .I1 (g3361), .I2 (g20391));
AN2X1 gate9473(.O (g29332), .I1 (g29107), .I2 (g22170));
AN2X1 gate9474(.O (g23657), .I1 (g19401), .I2 (g11941));
AN2X1 gate9475(.O (g28617), .I1 (g27533), .I2 (g20552));
AN3X1 gate9476(.O (g34097), .I1 (g33772), .I2 (g9104), .I3 (g18957));
AN2X1 gate9477(.O (g21955), .I1 (g5385), .I2 (g21514));
AN2X1 gate9478(.O (g23774), .I1 (g14867), .I2 (g21252));
AN2X1 gate9479(.O (g22064), .I1 (g15162), .I2 (g19210));
AN3X1 gate9480(.O (I24600), .I1 (g6077), .I2 (g6082), .I3 (g9946));
AN4X1 gate9481(.O (I31146), .I1 (g30735), .I2 (g31821), .I3 (g32666), .I4 (g32667));
AN2X1 gate9482(.O (g25026), .I1 (g22929), .I2 (g10503));
AN2X1 gate9483(.O (g34104), .I1 (g33916), .I2 (g23639));
AN2X1 gate9484(.O (g27117), .I1 (g26055), .I2 (g16528));
AN2X1 gate9485(.O (g21879), .I1 (g4132), .I2 (g19801));
AN2X1 gate9486(.O (g34811), .I1 (g14165), .I2 (g34766));
AN2X1 gate9487(.O (g21970), .I1 (g5401), .I2 (g21514));
AN2X1 gate9488(.O (g18143), .I1 (g586), .I2 (g17533));
AN2X1 gate9489(.O (g24502), .I1 (g23428), .I2 (g13223));
AN2X1 gate9490(.O (g28201), .I1 (g27499), .I2 (g16720));
AN2X1 gate9491(.O (g19536), .I1 (g518), .I2 (g16768));
AN2X1 gate9492(.O (g19948), .I1 (g17515), .I2 (g16320));
AN2X1 gate9493(.O (g29962), .I1 (g23616), .I2 (g28959));
AN2X1 gate9494(.O (g21878), .I1 (g4129), .I2 (g19801));
AN3X1 gate9495(.O (I16695), .I1 (g10207), .I2 (g12523), .I3 (g12463));
AN2X1 gate9496(.O (g32127), .I1 (g31624), .I2 (g29950));
AN2X1 gate9497(.O (g31541), .I1 (g22536), .I2 (g29348));
AN2X1 gate9498(.O (g24618), .I1 (g22625), .I2 (g19672));
AN2X1 gate9499(.O (g26229), .I1 (g1724), .I2 (g25275));
AN3X1 gate9500(.O (g33473), .I1 (g32549), .I2 (I31061), .I3 (I31062));
AN2X1 gate9501(.O (g18169), .I1 (g676), .I2 (g17433));
AN2X1 gate9502(.O (g21886), .I1 (g4153), .I2 (g19801));
AN2X1 gate9503(.O (g27568), .I1 (g26576), .I2 (g17791));
AN2X1 gate9504(.O (g18791), .I1 (g6044), .I2 (g15634));
AN2X1 gate9505(.O (g31789), .I1 (g30201), .I2 (g24013));
AN2X1 gate9506(.O (g28467), .I1 (g26993), .I2 (g12295));
AN2X1 gate9507(.O (g28494), .I1 (g27973), .I2 (g17741));
AN2X1 gate9508(.O (g33789), .I1 (g33159), .I2 (g23022));
AN2X1 gate9509(.O (g21792), .I1 (g3396), .I2 (g20391));
AN2X1 gate9510(.O (g16591), .I1 (g5256), .I2 (g14879));
AN2X1 gate9511(.O (g22009), .I1 (g5782), .I2 (g21562));
AN2X1 gate9512(.O (g22665), .I1 (g17174), .I2 (g20905));
AN2X1 gate9513(.O (g18168), .I1 (g681), .I2 (g17433));
AN2X1 gate9514(.O (g18410), .I1 (g2079), .I2 (g15373));
AN2X1 gate9515(.O (g21967), .I1 (g5456), .I2 (g21514));
AN2X1 gate9516(.O (g21994), .I1 (g5607), .I2 (g19074));
AN2X1 gate9517(.O (g31788), .I1 (g21352), .I2 (g29385));
AN2X1 gate9518(.O (g33724), .I1 (g14145), .I2 (g33258));
AN2X1 gate9519(.O (g32376), .I1 (g2689), .I2 (g31710));
AN2X1 gate9520(.O (g19564), .I1 (g17175), .I2 (g13976));
AN2X1 gate9521(.O (g33359), .I1 (g32252), .I2 (g20853));
AN2X1 gate9522(.O (g25149), .I1 (g14030), .I2 (g23546));
AN2X1 gate9523(.O (g17693), .I1 (g1306), .I2 (g13291));
AN2X1 gate9524(.O (g22008), .I1 (g5774), .I2 (g21562));
AN2X1 gate9525(.O (g32103), .I1 (g31609), .I2 (g29905));
AN2X1 gate9526(.O (g24286), .I1 (g4405), .I2 (g22550));
AN2X1 gate9527(.O (g18479), .I1 (g2449), .I2 (g15426));
AN2X1 gate9528(.O (g18666), .I1 (g4593), .I2 (g17367));
AN2X1 gate9529(.O (g33829), .I1 (g33240), .I2 (g20164));
AN2X1 gate9530(.O (g18363), .I1 (g1840), .I2 (g17955));
AN2X1 gate9531(.O (g32095), .I1 (g7619), .I2 (g30825));
AN2X1 gate9532(.O (g18217), .I1 (g15063), .I2 (g16100));
AN2X1 gate9533(.O (g33434), .I1 (g32239), .I2 (g29702));
AN2X1 gate9534(.O (g24306), .I1 (g4483), .I2 (g22228));
AN2X1 gate9535(.O (g33358), .I1 (g32249), .I2 (g20778));
AN2X1 gate9536(.O (g25148), .I1 (g16867), .I2 (g23545));
AN2X1 gate9537(.O (g11496), .I1 (g4382), .I2 (g7495));
AN2X1 gate9538(.O (g15871), .I1 (g3203), .I2 (g13951));
AN2X1 gate9539(.O (g18478), .I1 (g2445), .I2 (g15426));
AN2X1 gate9540(.O (g30133), .I1 (g28591), .I2 (g21179));
AN2X1 gate9541(.O (g33828), .I1 (g33090), .I2 (g24411));
AN2X1 gate9542(.O (g28352), .I1 (g10014), .I2 (g27705));
AN4X1 gate9543(.O (g11111), .I1 (g5297), .I2 (g7004), .I3 (g5283), .I4 (g9780));
AN2X1 gate9544(.O (g14875), .I1 (g1495), .I2 (g10939));
AN2X1 gate9545(.O (g34133), .I1 (g33845), .I2 (g23958));
AN2X1 gate9546(.O (g21919), .I1 (g15144), .I2 (g21468));
AN2X1 gate9547(.O (g30229), .I1 (g28716), .I2 (g23904));
AN2X1 gate9548(.O (g25104), .I1 (g16800), .I2 (g23504));
AN2X1 gate9549(.O (g11978), .I1 (g2629), .I2 (g7462));
AN2X1 gate9550(.O (g26310), .I1 (g2102), .I2 (g25389));
AN2X1 gate9551(.O (g23919), .I1 (g4122), .I2 (g19546));
AN2X1 gate9552(.O (g32181), .I1 (g31020), .I2 (g19912));
AN2X1 gate9553(.O (g33121), .I1 (g8748), .I2 (g32212));
AN2X1 gate9554(.O (g18486), .I1 (g2485), .I2 (g15426));
AN2X1 gate9555(.O (g27230), .I1 (g25906), .I2 (g19558));
AN2X1 gate9556(.O (g27293), .I1 (g9972), .I2 (g26655));
AN2X1 gate9557(.O (g29613), .I1 (g28208), .I2 (g19763));
AN2X1 gate9558(.O (g28266), .I1 (g23748), .I2 (g27714));
AN2X1 gate9559(.O (g19062), .I1 (g446), .I2 (g16180));
AN2X1 gate9560(.O (g33344), .I1 (g32228), .I2 (g20670));
AN2X1 gate9561(.O (g14218), .I1 (g875), .I2 (g10632));
AN2X1 gate9562(.O (g21918), .I1 (g5097), .I2 (g21468));
AN2X1 gate9563(.O (g30228), .I1 (g28715), .I2 (g23903));
AN2X1 gate9564(.O (g26379), .I1 (g19904), .I2 (g25546));
AN2X1 gate9565(.O (g18556), .I1 (g2823), .I2 (g15277));
AN2X1 gate9566(.O (g25971), .I1 (g1917), .I2 (g24992));
AN2X1 gate9567(.O (g24187), .I1 (g305), .I2 (g22722));
AN2X1 gate9568(.O (g34228), .I1 (g33750), .I2 (g22942));
AN2X1 gate9569(.O (g30011), .I1 (g29183), .I2 (g12930));
AN2X1 gate9570(.O (g27265), .I1 (g26785), .I2 (g26759));
AN4X1 gate9571(.O (I31226), .I1 (g29385), .I2 (g32781), .I3 (g32782), .I4 (g32783));
AN2X1 gate9572(.O (g16844), .I1 (g7212), .I2 (g13000));
AN2X1 gate9573(.O (g18580), .I1 (g2907), .I2 (g16349));
AN2X1 gate9574(.O (g26050), .I1 (g9630), .I2 (g25047));
AN4X1 gate9575(.O (g27416), .I1 (g8046), .I2 (g26314), .I3 (g9187), .I4 (g504));
AN2X1 gate9576(.O (g26378), .I1 (g19576), .I2 (g25544));
AN2X1 gate9577(.O (g13384), .I1 (g4944), .I2 (g11804));
AN2X1 gate9578(.O (g29605), .I1 (g2445), .I2 (g28973));
AN2X1 gate9579(.O (g18223), .I1 (g1030), .I2 (g16100));
AN2X1 gate9580(.O (g23599), .I1 (g19050), .I2 (g9104));
AN2X1 gate9581(.O (g27992), .I1 (g26800), .I2 (g23964));
AN2X1 gate9582(.O (g22074), .I1 (g6239), .I2 (g19210));
AN2X1 gate9583(.O (g27391), .I1 (g26549), .I2 (g17505));
AN2X1 gate9584(.O (g24143), .I1 (g17694), .I2 (g21659));
AN2X1 gate9585(.O (g25368), .I1 (g6946), .I2 (g22408));
AN2X1 gate9586(.O (g27510), .I1 (g26576), .I2 (g17687));
AN2X1 gate9587(.O (g34582), .I1 (g7764), .I2 (g34313));
AN2X1 gate9588(.O (g32190), .I1 (g142), .I2 (g31233));
AN2X1 gate9589(.O (g26096), .I1 (g9733), .I2 (g25268));
AN2X1 gate9590(.O (g29951), .I1 (g1874), .I2 (g28786));
AN2X1 gate9591(.O (g18110), .I1 (g441), .I2 (g17015));
AN2X1 gate9592(.O (g34310), .I1 (g14003), .I2 (g34162));
AN2X1 gate9593(.O (g25850), .I1 (g3502), .I2 (g24636));
AN2X1 gate9594(.O (g15911), .I1 (g3111), .I2 (g13530));
AN2X1 gate9595(.O (g28588), .I1 (g27489), .I2 (g20499));
AN2X1 gate9596(.O (g28524), .I1 (g6821), .I2 (g27084));
AN4X1 gate9597(.O (I31127), .I1 (g32638), .I2 (g32639), .I3 (g32640), .I4 (g32641));
AN2X1 gate9598(.O (g18321), .I1 (g1620), .I2 (g17873));
AN3X1 gate9599(.O (g24884), .I1 (g3401), .I2 (g23555), .I3 (I24051));
AN2X1 gate9600(.O (g30925), .I1 (g29908), .I2 (g23309));
AN2X1 gate9601(.O (g21817), .I1 (g3606), .I2 (g20924));
AN2X1 gate9602(.O (g11019), .I1 (g5092), .I2 (g9036));
AN2X1 gate9603(.O (g18179), .I1 (g763), .I2 (g17328));
AN2X1 gate9604(.O (g13019), .I1 (g194), .I2 (g11737));
AN2X1 gate9605(.O (g18531), .I1 (g2719), .I2 (g15277));
AN2X1 gate9606(.O (g30112), .I1 (g28566), .I2 (g20919));
AN2X1 gate9607(.O (g28477), .I1 (g27966), .I2 (g17676));
AN2X1 gate9608(.O (g33760), .I1 (g33143), .I2 (g20328));
AN2X1 gate9609(.O (g24410), .I1 (g3817), .I2 (g23139));
AN2X1 gate9610(.O (g32089), .I1 (g27261), .I2 (g31021));
AN2X1 gate9611(.O (g25229), .I1 (g7636), .I2 (g22654));
AN2X1 gate9612(.O (g30050), .I1 (g22545), .I2 (g28126));
AN2X1 gate9613(.O (g29795), .I1 (g28344), .I2 (g23257));
AN3X1 gate9614(.O (g34112), .I1 (g22957), .I2 (g9104), .I3 (g33778));
AN3X1 gate9615(.O (g11018), .I1 (g7655), .I2 (g7643), .I3 (g7627));
AN2X1 gate9616(.O (g18178), .I1 (g758), .I2 (g17328));
AN2X1 gate9617(.O (g18740), .I1 (g4572), .I2 (g17384));
AN2X1 gate9618(.O (g26857), .I1 (g25062), .I2 (g25049));
AN2X1 gate9619(.O (g34050), .I1 (g33772), .I2 (g22942));
AN2X1 gate9620(.O (g21977), .I1 (g5535), .I2 (g19074));
AN2X1 gate9621(.O (g22092), .I1 (g6419), .I2 (g18833));
AN2X1 gate9622(.O (g23532), .I1 (g19400), .I2 (g11852));
AN2X1 gate9623(.O (g23901), .I1 (g19606), .I2 (g7963));
AN2X1 gate9624(.O (g34378), .I1 (g13095), .I2 (g34053));
AN2X1 gate9625(.O (g16025), .I1 (g446), .I2 (g14063));
AN3X1 gate9626(.O (g33506), .I1 (g32788), .I2 (I31226), .I3 (I31227));
AN3X1 gate9627(.O (I24530), .I1 (g9501), .I2 (g9733), .I3 (g5747));
AN2X1 gate9628(.O (g32088), .I1 (g27241), .I2 (g31070));
AN2X1 gate9629(.O (g24666), .I1 (g11753), .I2 (g22975));
AN2X1 gate9630(.O (g22518), .I1 (g12982), .I2 (g19398));
AN2X1 gate9631(.O (g21783), .I1 (g3419), .I2 (g20391));
AN4X1 gate9632(.O (I31297), .I1 (g32884), .I2 (g32885), .I3 (g32886), .I4 (g32887));
AN2X1 gate9633(.O (g24217), .I1 (g18200), .I2 (g22594));
AN2X1 gate9634(.O (g18186), .I1 (g753), .I2 (g17328));
AN2X1 gate9635(.O (g15785), .I1 (g3558), .I2 (g14107));
AN2X1 gate9636(.O (g18676), .I1 (g4358), .I2 (g15758));
AN2X1 gate9637(.O (g18685), .I1 (g4688), .I2 (g15885));
AN2X1 gate9638(.O (g34386), .I1 (g10800), .I2 (g34060));
AN2X1 gate9639(.O (g18373), .I1 (g1890), .I2 (g15171));
AN2X1 gate9640(.O (g29514), .I1 (g1608), .I2 (g28780));
AN2X1 gate9641(.O (g24015), .I1 (g19540), .I2 (g10951));
AN2X1 gate9642(.O (g30096), .I1 (g28546), .I2 (g20770));
AN2X1 gate9643(.O (g22637), .I1 (g19363), .I2 (g19489));
AN2X1 gate9644(.O (g17176), .I1 (g8616), .I2 (g13008));
AN2X1 gate9645(.O (g34742), .I1 (g9000), .I2 (g34698));
AN2X1 gate9646(.O (g28616), .I1 (g27532), .I2 (g20551));
AN3X1 gate9647(.O (g34096), .I1 (g22957), .I2 (g9104), .I3 (g33772));
AN2X1 gate9648(.O (g18654), .I1 (g4146), .I2 (g16249));
AN2X1 gate9649(.O (g16203), .I1 (g5821), .I2 (g14297));
AN2X1 gate9650(.O (g28313), .I1 (g27231), .I2 (g19766));
AN2X1 gate9651(.O (g27116), .I1 (g26026), .I2 (g16527));
AN4X1 gate9652(.O (I27509), .I1 (g24084), .I2 (g24085), .I3 (g24086), .I4 (g24087));
AN2X1 gate9653(.O (g21823), .I1 (g3731), .I2 (g20453));
AN2X1 gate9654(.O (g27615), .I1 (g26789), .I2 (g26770));
AN2X1 gate9655(.O (g18800), .I1 (g6187), .I2 (g15348));
AN2X1 gate9656(.O (g15859), .I1 (g3610), .I2 (g13923));
AN4X1 gate9657(.O (I31181), .I1 (g29385), .I2 (g32716), .I3 (g32717), .I4 (g32718));
AN2X1 gate9658(.O (g18417), .I1 (g2116), .I2 (g15373));
AN2X1 gate9659(.O (g24556), .I1 (g4035), .I2 (g23341));
AN2X1 gate9660(.O (g28285), .I1 (g9657), .I2 (g27717));
AN2X1 gate9661(.O (g34681), .I1 (g34491), .I2 (g19438));
AN4X1 gate9662(.O (I27508), .I1 (g19935), .I2 (g24082), .I3 (g24083), .I4 (g28033));
AN2X1 gate9663(.O (g15858), .I1 (g3542), .I2 (g14045));
AN2X1 gate9664(.O (g27041), .I1 (g8519), .I2 (g26330));
AN2X1 gate9665(.O (g32126), .I1 (g31601), .I2 (g29948));
AN2X1 gate9666(.O (g18334), .I1 (g1696), .I2 (g17873));
AN2X1 gate9667(.O (g27275), .I1 (g25945), .I2 (g19745));
AN2X1 gate9668(.O (g19756), .I1 (g9899), .I2 (g17154));
AN2X1 gate9669(.O (g33927), .I1 (g33094), .I2 (g21412));
AN3X1 gate9670(.O (g28254), .I1 (g7268), .I2 (g1668), .I3 (g27395));
AN2X1 gate9671(.O (g27430), .I1 (g26488), .I2 (g17579));
AN2X1 gate9672(.O (g34857), .I1 (g16540), .I2 (g34813));
AN2X1 gate9673(.O (g10822), .I1 (g4264), .I2 (g8514));
AN2X1 gate9674(.O (g24223), .I1 (g239), .I2 (g22594));
AN2X1 gate9675(.O (g27493), .I1 (g246), .I2 (g26837));
AN2X1 gate9676(.O (g16957), .I1 (g13064), .I2 (g10418));
AN2X1 gate9677(.O (g25959), .I1 (g1648), .I2 (g24963));
AN2X1 gate9678(.O (g30730), .I1 (g26346), .I2 (g29778));
AN2X1 gate9679(.O (g25925), .I1 (g24990), .I2 (g23234));
AN2X1 gate9680(.O (g28466), .I1 (g27960), .I2 (g17637));
AN2X1 gate9681(.O (g25112), .I1 (g10428), .I2 (g23510));
AN2X1 gate9682(.O (g21966), .I1 (g5406), .I2 (g21514));
AN2X1 gate9683(.O (g18762), .I1 (g5475), .I2 (g17929));
AN2X1 gate9684(.O (g25050), .I1 (g13056), .I2 (g22312));
AN2X1 gate9685(.O (g20084), .I1 (g11591), .I2 (g16609));
AN2X1 gate9686(.O (g32339), .I1 (g31474), .I2 (g20672));
AN2X1 gate9687(.O (g31240), .I1 (g14793), .I2 (g30206));
AN2X1 gate9688(.O (g19350), .I1 (g15968), .I2 (g13505));
AN2X1 gate9689(.O (g34765), .I1 (g34692), .I2 (g20057));
AN2X1 gate9690(.O (g27340), .I1 (g10199), .I2 (g26784));
AN2X1 gate9691(.O (g27035), .I1 (g26348), .I2 (g1500));
AN2X1 gate9692(.O (g18423), .I1 (g12851), .I2 (g18008));
AN2X1 gate9693(.O (g29789), .I1 (g28270), .I2 (g10233));
AN2X1 gate9694(.O (g32338), .I1 (g31466), .I2 (g20668));
AN3X1 gate9695(.O (g33491), .I1 (g32679), .I2 (I31151), .I3 (I31152));
AN2X1 gate9696(.O (g33903), .I1 (g33447), .I2 (g19146));
AN2X1 gate9697(.O (g24922), .I1 (g4831), .I2 (g23931));
AN2X1 gate9698(.O (g26129), .I1 (g2384), .I2 (g25121));
AN2X1 gate9699(.O (g18216), .I1 (g967), .I2 (g15979));
AN2X1 gate9700(.O (g24321), .I1 (g4558), .I2 (g22228));
AN2X1 gate9701(.O (g16699), .I1 (g7134), .I2 (g12933));
AN2X1 gate9702(.O (g27684), .I1 (g26386), .I2 (g20657));
AN2X1 gate9703(.O (g28642), .I1 (g27555), .I2 (g20598));
AN2X1 gate9704(.O (g18587), .I1 (g2980), .I2 (g16349));
AN2X1 gate9705(.O (g25096), .I1 (g23778), .I2 (g20560));
AN2X1 gate9706(.O (g29788), .I1 (g28335), .I2 (g23250));
AN2X1 gate9707(.O (g26128), .I1 (g2319), .I2 (g25120));
AN2X1 gate9708(.O (g14589), .I1 (g10586), .I2 (g10569));
AN2X1 gate9709(.O (g29535), .I1 (g2303), .I2 (g28871));
AN4X1 gate9710(.O (I31211), .I1 (g31021), .I2 (g31833), .I3 (g32759), .I4 (g32760));
AN2X1 gate9711(.O (g27517), .I1 (g26400), .I2 (g17707));
AN2X1 gate9712(.O (g10588), .I1 (g7004), .I2 (g5297));
AN2X1 gate9713(.O (g18909), .I1 (g16226), .I2 (g13570));
AN2X1 gate9714(.O (g32197), .I1 (g31144), .I2 (g20088));
AN2X1 gate9715(.O (g18543), .I1 (g2779), .I2 (g15277));
AN2X1 gate9716(.O (g26323), .I1 (g10262), .I2 (g25273));
AN2X1 gate9717(.O (g24186), .I1 (g18102), .I2 (g22722));
AN2X1 gate9718(.O (g14588), .I1 (g11957), .I2 (g11974));
AN2X1 gate9719(.O (g24676), .I1 (g2748), .I2 (g23782));
AN3X1 gate9720(.O (I16721), .I1 (g10224), .I2 (g12589), .I3 (g12525));
AN2X1 gate9721(.O (g18117), .I1 (g464), .I2 (g17015));
AN2X1 gate9722(.O (g16427), .I1 (g5216), .I2 (g14876));
AN2X1 gate9723(.O (g25802), .I1 (g8106), .I2 (g24586));
AN2X1 gate9724(.O (g22083), .I1 (g6287), .I2 (g19210));
AN2X1 gate9725(.O (g32411), .I1 (g31119), .I2 (g13469));
AN2X1 gate9726(.O (g23023), .I1 (g650), .I2 (g20248));
AN2X1 gate9727(.O (g19691), .I1 (g9614), .I2 (g17085));
AN2X1 gate9728(.O (g24654), .I1 (g11735), .I2 (g22922));
AN2X1 gate9729(.O (g28630), .I1 (g27544), .I2 (g20575));
AN2X1 gate9730(.O (g29344), .I1 (g29168), .I2 (g18932));
AN2X1 gate9731(.O (g18569), .I1 (g94), .I2 (g16349));
AN2X1 gate9732(.O (g30002), .I1 (g28481), .I2 (g23487));
AN2X1 gate9733(.O (g27130), .I1 (g26026), .I2 (g16585));
AN2X1 gate9734(.O (g30057), .I1 (g29144), .I2 (g9462));
AN2X1 gate9735(.O (g22622), .I1 (g19336), .I2 (g19469));
AN2X1 gate9736(.O (g18568), .I1 (g37), .I2 (g16349));
AN2X1 gate9737(.O (g18747), .I1 (g5138), .I2 (g17847));
AN2X1 gate9738(.O (g25765), .I1 (g24989), .I2 (g24973));
AN2X1 gate9739(.O (g27362), .I1 (g26080), .I2 (g20036));
AN2X1 gate9740(.O (g31990), .I1 (g31772), .I2 (g18945));
AN2X1 gate9741(.O (g33899), .I1 (g32132), .I2 (g33335));
AN2X1 gate9742(.O (g18242), .I1 (g962), .I2 (g16431));
AN2X1 gate9743(.O (g10616), .I1 (g7998), .I2 (g174));
AN2X1 gate9744(.O (g27523), .I1 (g26549), .I2 (g17718));
AN2X1 gate9745(.O (g30245), .I1 (g28733), .I2 (g23935));
AN4X1 gate9746(.O (I31126), .I1 (g30673), .I2 (g31818), .I3 (g32636), .I4 (g32637));
AN2X1 gate9747(.O (g26232), .I1 (g2193), .I2 (g25396));
AN2X1 gate9748(.O (g33898), .I1 (g33419), .I2 (g15655));
AN2X1 gate9749(.O (g21816), .I1 (g3602), .I2 (g20924));
AN2X1 gate9750(.O (g18123), .I1 (g479), .I2 (g16886));
AN2X1 gate9751(.O (g18814), .I1 (g6519), .I2 (g15483));
AN2X1 gate9752(.O (g33719), .I1 (g33141), .I2 (g19433));
AN2X1 gate9753(.O (g24762), .I1 (g655), .I2 (g23573));
AN3X1 gate9754(.O (g10704), .I1 (g2145), .I2 (g10200), .I3 (g2130));
AN2X1 gate9755(.O (g34533), .I1 (g34318), .I2 (g19731));
AN2X1 gate9756(.O (g18751), .I1 (g5156), .I2 (g17847));
AN2X1 gate9757(.O (g18807), .I1 (g6386), .I2 (g15656));
AN2X1 gate9758(.O (g21976), .I1 (g5527), .I2 (g19074));
AN2X1 gate9759(.O (g21985), .I1 (g5571), .I2 (g19074));
AN2X1 gate9760(.O (g15902), .I1 (g441), .I2 (g13975));
AN2X1 gate9761(.O (g18772), .I1 (g5689), .I2 (g15615));
AN2X1 gate9762(.O (g28555), .I1 (g27429), .I2 (g20373));
AN2X1 gate9763(.O (g33718), .I1 (g33147), .I2 (g19432));
AN2X1 gate9764(.O (g34298), .I1 (g8679), .I2 (g34132));
AN2X1 gate9765(.O (g28454), .I1 (g26976), .I2 (g12233));
AN3X1 gate9766(.O (g33521), .I1 (g32895), .I2 (I31301), .I3 (I31302));
AN2X1 gate9767(.O (g18974), .I1 (g174), .I2 (g16127));
AN4X1 gate9768(.O (g26261), .I1 (g24688), .I2 (g10678), .I3 (g8778), .I4 (g8757));
AN2X1 gate9769(.O (g32315), .I1 (g31306), .I2 (g23517));
AN2X1 gate9770(.O (g24423), .I1 (g4950), .I2 (g22897));
AN2X1 gate9771(.O (g21752), .I1 (g3171), .I2 (g20785));
AN4X1 gate9772(.O (g27727), .I1 (g22432), .I2 (g25211), .I3 (g26424), .I4 (g26195));
AN4X1 gate9773(.O (I31296), .I1 (g30937), .I2 (g31848), .I3 (g32882), .I4 (g32883));
AN2X1 gate9774(.O (g18639), .I1 (g3831), .I2 (g17096));
AN2X1 gate9775(.O (g28570), .I1 (g27456), .I2 (g20434));
AN2X1 gate9776(.O (g28712), .I1 (g27590), .I2 (g20708));
AN2X1 gate9777(.O (g21954), .I1 (g5381), .I2 (g21514));
AN2X1 gate9778(.O (g27222), .I1 (g26055), .I2 (g13932));
AN2X1 gate9779(.O (g29760), .I1 (g28309), .I2 (g23227));
AN2X1 gate9780(.O (g33832), .I1 (g33088), .I2 (g27991));
AN2X1 gate9781(.O (g18230), .I1 (g1111), .I2 (g16326));
AN4X1 gate9782(.O (g29029), .I1 (g14506), .I2 (g25227), .I3 (g26424), .I4 (g27494));
AN2X1 gate9783(.O (g17139), .I1 (g8635), .I2 (g12967));
AN2X1 gate9784(.O (g18293), .I1 (g1484), .I2 (g16449));
AN4X1 gate9785(.O (g17653), .I1 (g11547), .I2 (g11592), .I3 (g6789), .I4 (I18620));
AN2X1 gate9786(.O (g15738), .I1 (g1111), .I2 (g13260));
AN2X1 gate9787(.O (g18638), .I1 (g3827), .I2 (g17096));
AN2X1 gate9788(.O (g27437), .I1 (g26576), .I2 (g17589));
AN2X1 gate9789(.O (g33440), .I1 (g32250), .I2 (g29719));
AN2X1 gate9790(.O (g32055), .I1 (g10999), .I2 (g30825));
AN2X1 gate9791(.O (g17138), .I1 (g255), .I2 (g13239));
AN2X1 gate9792(.O (g18265), .I1 (g1270), .I2 (g16000));
AN2X1 gate9793(.O (g25129), .I1 (g17682), .I2 (g23527));
AN2X1 gate9794(.O (g15699), .I1 (g1437), .I2 (g13861));
AN2X1 gate9795(.O (g30232), .I1 (g28719), .I2 (g23912));
AN2X1 gate9796(.O (g32111), .I1 (g31616), .I2 (g29922));
AN2X1 gate9797(.O (g18416), .I1 (g2112), .I2 (g15373));
AN2X1 gate9798(.O (g25057), .I1 (g23275), .I2 (g20511));
AN2X1 gate9799(.O (g32070), .I1 (g10967), .I2 (g30825));
AN2X1 gate9800(.O (g33861), .I1 (g33271), .I2 (g20502));
AN2X1 gate9801(.O (g28239), .I1 (g27135), .I2 (g19659));
AN2X1 gate9802(.O (g25128), .I1 (g17418), .I2 (g23525));
AN2X1 gate9803(.O (g17636), .I1 (g10829), .I2 (g13463));
AN2X1 gate9804(.O (g11916), .I1 (g2227), .I2 (g7328));
AN2X1 gate9805(.O (g33247), .I1 (g32130), .I2 (g19980));
AN2X1 gate9806(.O (g28567), .I1 (g6832), .I2 (g27101));
AN4X1 gate9807(.O (I31197), .I1 (g32740), .I2 (g32741), .I3 (g32742), .I4 (g32743));
AN2X1 gate9808(.O (g27347), .I1 (g26400), .I2 (g17390));
AN2X1 gate9809(.O (g18992), .I1 (g8341), .I2 (g16171));
AN2X1 gate9810(.O (g18391), .I1 (g1982), .I2 (g15171));
AN3X1 gate9811(.O (g24908), .I1 (g3752), .I2 (g23239), .I3 (I24075));
AN2X1 gate9812(.O (g28238), .I1 (g27133), .I2 (g19658));
AN2X1 gate9813(.O (g21842), .I1 (g3863), .I2 (g21070));
AN2X1 gate9814(.O (g18510), .I1 (g2625), .I2 (g15509));
AN2X1 gate9815(.O (g30261), .I1 (g28772), .I2 (g23961));
AN2X1 gate9816(.O (g23392), .I1 (g7247), .I2 (g21430));
AN2X1 gate9817(.O (g24569), .I1 (g5115), .I2 (g23382));
AN2X1 gate9818(.O (g25323), .I1 (g6888), .I2 (g22359));
AN2X1 gate9819(.O (g31324), .I1 (g30171), .I2 (g27937));
AN2X1 gate9820(.O (g33099), .I1 (g32395), .I2 (g18944));
AN2X1 gate9821(.O (g13287), .I1 (g1221), .I2 (g11472));
AN2X1 gate9822(.O (g27600), .I1 (g26755), .I2 (g26725));
AN4X1 gate9823(.O (g10733), .I1 (g3639), .I2 (g6905), .I3 (g3625), .I4 (g8542));
AN2X1 gate9824(.O (g18579), .I1 (g2984), .I2 (g16349));
AN2X1 gate9825(.O (g31777), .I1 (g21343), .I2 (g29385));
AN2X1 gate9826(.O (g33701), .I1 (g33162), .I2 (g16305));
AN2X1 gate9827(.O (g24747), .I1 (g17510), .I2 (g22417));
AN2X1 gate9828(.O (g32067), .I1 (g4727), .I2 (g30614));
AN2X1 gate9829(.O (g21559), .I1 (g16236), .I2 (g10897));
AN2X1 gate9830(.O (g31272), .I1 (g30117), .I2 (g27742));
AN3X1 gate9831(.O (I16618), .I1 (g10124), .I2 (g12341), .I3 (g12293));
AN2X1 gate9832(.O (g15632), .I1 (g3494), .I2 (g13555));
AN2X1 gate9833(.O (g28185), .I1 (g27026), .I2 (g19435));
AN3X1 gate9834(.O (g10874), .I1 (g7791), .I2 (g6219), .I3 (g6227));
AN2X1 gate9835(.O (g18578), .I1 (g2873), .I2 (g16349));
AN2X1 gate9836(.O (g25775), .I1 (g2922), .I2 (g24568));
AN2X1 gate9837(.O (g23424), .I1 (g7345), .I2 (g21556));
AN2X1 gate9838(.O (g27351), .I1 (g10218), .I2 (g26804));
AN2X1 gate9839(.O (g27372), .I1 (g26488), .I2 (g17476));
AN2X1 gate9840(.O (g19768), .I1 (g2803), .I2 (g15833));
AN2X1 gate9841(.O (g14874), .I1 (g1099), .I2 (g10909));
AN2X1 gate9842(.O (g16671), .I1 (g6275), .I2 (g14817));
AN2X1 gate9843(.O (g21558), .I1 (g15904), .I2 (g13729));
AN2X1 gate9844(.O (g27821), .I1 (g7680), .I2 (g25892));
AN2X1 gate9845(.O (g32150), .I1 (g31624), .I2 (g29995));
AN2X1 gate9846(.O (g28154), .I1 (g8492), .I2 (g27306));
AN2X1 gate9847(.O (g18586), .I1 (g2886), .I2 (g16349));
AN2X1 gate9848(.O (g29649), .I1 (g2241), .I2 (g28678));
AN3X1 gate9849(.O (g33462), .I1 (g32470), .I2 (I31006), .I3 (I31007));
AN2X1 gate9850(.O (g21830), .I1 (g3774), .I2 (g20453));
AN2X1 gate9851(.O (g26611), .I1 (g24935), .I2 (g20580));
AN2X1 gate9852(.O (g20751), .I1 (g16260), .I2 (g4836));
AN2X1 gate9853(.O (g10665), .I1 (g209), .I2 (g8292));
AN2X1 gate9854(.O (g28637), .I1 (g22399), .I2 (g27011));
AN2X1 gate9855(.O (g18442), .I1 (g2259), .I2 (g18008));
AN2X1 gate9856(.O (g32019), .I1 (g30579), .I2 (g22358));
AN2X1 gate9857(.O (g24772), .I1 (g16287), .I2 (g23061));
AN2X1 gate9858(.O (g29648), .I1 (g2112), .I2 (g29121));
AN2X1 gate9859(.O (g27264), .I1 (g25941), .I2 (g19714));
AN2X1 gate9860(.O (g22115), .I1 (g6573), .I2 (g19277));
AN2X1 gate9861(.O (g27137), .I1 (g26026), .I2 (g16606));
AN2X1 gate9862(.O (g21865), .I1 (g3965), .I2 (g21070));
AN2X1 gate9863(.O (g31140), .I1 (g2102), .I2 (g30037));
AN2X1 gate9864(.O (g32196), .I1 (g27587), .I2 (g31376));
AN2X1 gate9865(.O (g13942), .I1 (g5897), .I2 (g12512));
AN2X1 gate9866(.O (g24639), .I1 (g6181), .I2 (g23699));
AN2X1 gate9867(.O (g32018), .I1 (g4146), .I2 (g30937));
AN2X1 gate9868(.O (g26271), .I1 (g1992), .I2 (g25341));
AN2X1 gate9869(.O (g29604), .I1 (g2315), .I2 (g28966));
AN3X1 gate9870(.O (g30316), .I1 (g29199), .I2 (g7097), .I3 (g6682));
AN2X1 gate9871(.O (g21713), .I1 (g298), .I2 (g20283));
AN2X1 gate9872(.O (g34499), .I1 (g31288), .I2 (g34339));
AN2X1 gate9873(.O (g24230), .I1 (g901), .I2 (g22594));
AN3X1 gate9874(.O (g13156), .I1 (g10816), .I2 (g10812), .I3 (g10805));
AN2X1 gate9875(.O (g18116), .I1 (g168), .I2 (g17015));
AN2X1 gate9876(.O (g24293), .I1 (g4438), .I2 (g22550));
AN2X1 gate9877(.O (g18615), .I1 (g3347), .I2 (g17200));
AN2X1 gate9878(.O (g22052), .I1 (g6113), .I2 (g21611));
AN3X1 gate9879(.O (g10476), .I1 (g7244), .I2 (g7259), .I3 (I13862));
AN2X1 gate9880(.O (g24638), .I1 (g22763), .I2 (g19690));
AN2X1 gate9881(.O (g29770), .I1 (g28320), .I2 (g23238));
AN2X1 gate9882(.O (g16190), .I1 (g14626), .I2 (g11810));
AN2X1 gate9883(.O (g29563), .I1 (g1616), .I2 (g28853));
AN4X1 gate9884(.O (I31202), .I1 (g32747), .I2 (g32748), .I3 (g32749), .I4 (g32750));
AN2X1 gate9885(.O (g34498), .I1 (g13888), .I2 (g34336));
AN2X1 gate9886(.O (g18720), .I1 (g15137), .I2 (g16795));
AN2X1 gate9887(.O (g26753), .I1 (g16024), .I2 (g24452));
AN4X1 gate9888(.O (I31257), .I1 (g32826), .I2 (g32827), .I3 (g32828), .I4 (g32829));
AN2X1 gate9889(.O (g25880), .I1 (g8443), .I2 (g24814));
AN4X1 gate9890(.O (g14555), .I1 (g12521), .I2 (g12356), .I3 (g12307), .I4 (I16671));
AN2X1 gate9891(.O (g24416), .I1 (g4939), .I2 (g22870));
AN2X1 gate9892(.O (g16520), .I1 (g5909), .I2 (g14965));
AN2X1 gate9893(.O (g21705), .I1 (g209), .I2 (g20283));
AN2X1 gate9894(.O (g30056), .I1 (g29165), .I2 (g12659));
AN2X1 gate9895(.O (g18275), .I1 (g15070), .I2 (g16136));
AN2X1 gate9896(.O (g26145), .I1 (g11962), .I2 (g25131));
AN4X1 gate9897(.O (I31111), .I1 (g31070), .I2 (g31815), .I3 (g32615), .I4 (g32616));
AN2X1 gate9898(.O (g18430), .I1 (g2204), .I2 (g18008));
AN2X1 gate9899(.O (g18746), .I1 (g5134), .I2 (g17847));
AN3X1 gate9900(.O (g27209), .I1 (g26213), .I2 (g8365), .I3 (g2051));
AN2X1 gate9901(.O (g32402), .I1 (g4888), .I2 (g30990));
AN2X1 gate9902(.O (g18493), .I1 (g2514), .I2 (g15426));
AN2X1 gate9903(.O (g33871), .I1 (g33281), .I2 (g20546));
AN2X1 gate9904(.O (g30080), .I1 (g28121), .I2 (g20674));
AN2X1 gate9905(.O (g28215), .I1 (g9264), .I2 (g27565));
AN2X1 gate9906(.O (g26650), .I1 (g10796), .I2 (g24424));
AN3X1 gate9907(.O (g34080), .I1 (g22957), .I2 (g9104), .I3 (g33750));
AN2X1 gate9908(.O (g16211), .I1 (g5445), .I2 (g14215));
AN2X1 gate9909(.O (g27208), .I1 (g9037), .I2 (g26598));
AN2X1 gate9910(.O (g18465), .I1 (g2384), .I2 (g15224));
AN2X1 gate9911(.O (g29767), .I1 (g28317), .I2 (g23236));
AN2X1 gate9912(.O (g29794), .I1 (g28342), .I2 (g23256));
AN2X1 gate9913(.O (g21188), .I1 (g7666), .I2 (g15705));
AN2X1 gate9914(.O (g33360), .I1 (g32253), .I2 (g20869));
AN2X1 gate9915(.O (g18237), .I1 (g1146), .I2 (g16326));
AN2X1 gate9916(.O (g29845), .I1 (g28375), .I2 (g23291));
AN2X1 gate9917(.O (g23188), .I1 (g13994), .I2 (g20025));
AN3X1 gate9918(.O (I16143), .I1 (g8751), .I2 (g11491), .I3 (g11445));
AN2X1 gate9919(.O (g28439), .I1 (g27273), .I2 (g10233));
AN2X1 gate9920(.O (g18340), .I1 (g1720), .I2 (g17873));
AN2X1 gate9921(.O (g29899), .I1 (g28428), .I2 (g23375));
AN2X1 gate9922(.O (g29990), .I1 (g29007), .I2 (g9239));
AN2X1 gate9923(.O (g21939), .I1 (g5224), .I2 (g18997));
AN2X1 gate9924(.O (g25831), .I1 (g3151), .I2 (g24623));
AN2X1 gate9925(.O (g15784), .I1 (g3235), .I2 (g13977));
AN2X1 gate9926(.O (g18806), .I1 (g6381), .I2 (g15656));
AN2X1 gate9927(.O (g18684), .I1 (g4681), .I2 (g15885));
AN2X1 gate9928(.O (g26393), .I1 (g19467), .I2 (g25558));
AN2X1 gate9929(.O (g14567), .I1 (g10568), .I2 (g10552));
AN2X1 gate9930(.O (g24835), .I1 (g8720), .I2 (g23233));
AN2X1 gate9931(.O (g29633), .I1 (g1978), .I2 (g29085));
AN4X1 gate9932(.O (I31067), .I1 (g32552), .I2 (g32553), .I3 (g32554), .I4 (g32555));
AN2X1 gate9933(.O (g24014), .I1 (g7933), .I2 (g19063));
AN2X1 gate9934(.O (g15103), .I1 (g4180), .I2 (g14454));
AN2X1 gate9935(.O (g34753), .I1 (g34676), .I2 (g19586));
AN2X1 gate9936(.O (g21938), .I1 (g5216), .I2 (g18997));
AN2X1 gate9937(.O (g18142), .I1 (g577), .I2 (g17533));
AN2X1 gate9938(.O (g34342), .I1 (g34103), .I2 (g19998));
AN2X1 gate9939(.O (g30145), .I1 (g28603), .I2 (g21247));
AN2X1 gate9940(.O (g30031), .I1 (g29071), .I2 (g10540));
AN2X1 gate9941(.O (g27614), .I1 (g26785), .I2 (g26759));
AN2X1 gate9942(.O (g32256), .I1 (g31249), .I2 (g20382));
AN2X1 gate9943(.O (g18517), .I1 (g2652), .I2 (g15509));
AN2X1 gate9944(.O (g27436), .I1 (g26576), .I2 (g17588));
AN2X1 gate9945(.O (g30199), .I1 (g28664), .I2 (g23861));
AN2X1 gate9946(.O (g29718), .I1 (g28512), .I2 (g11136));
AN2X1 gate9947(.O (g29521), .I1 (g1744), .I2 (g28824));
AN2X1 gate9948(.O (g16700), .I1 (g5208), .I2 (g14838));
AN2X1 gate9949(.O (g31220), .I1 (g30273), .I2 (g25202));
AN3X1 gate9950(.O (g33472), .I1 (g32542), .I2 (I31056), .I3 (I31057));
AN2X1 gate9951(.O (g16126), .I1 (g5495), .I2 (g14262));
AN2X1 gate9952(.O (g28284), .I1 (g11398), .I2 (g27994));
AN2X1 gate9953(.O (g10675), .I1 (g3436), .I2 (g8500));
AN2X1 gate9954(.O (g25989), .I1 (g25258), .I2 (g21012));
AN4X1 gate9955(.O (g27073), .I1 (g7121), .I2 (g3873), .I3 (g3881), .I4 (g26281));
AN2X1 gate9956(.O (g30198), .I1 (g28662), .I2 (g23860));
AN2X1 gate9957(.O (g32300), .I1 (g31274), .I2 (g20544));
AN2X1 gate9958(.O (g14185), .I1 (g8686), .I2 (g11744));
AN2X1 gate9959(.O (g25056), .I1 (g12779), .I2 (g23456));
AN2X1 gate9960(.O (g28304), .I1 (g27226), .I2 (g19753));
AN2X1 gate9961(.O (g33911), .I1 (g33137), .I2 (g10725));
AN2X1 gate9962(.O (g34198), .I1 (g33688), .I2 (g24491));
AN2X1 gate9963(.O (g26161), .I1 (g2518), .I2 (g25139));
AN2X1 gate9964(.O (g34529), .I1 (g34306), .I2 (g19634));
AN2X1 gate9965(.O (g21875), .I1 (g4116), .I2 (g19801));
AN2X1 gate9966(.O (g25988), .I1 (g9510), .I2 (g25016));
AN4X1 gate9967(.O (I31196), .I1 (g30825), .I2 (g31830), .I3 (g32738), .I4 (g32739));
AN2X1 gate9968(.O (g25924), .I1 (g24976), .I2 (g16846));
AN2X1 gate9969(.O (g27346), .I1 (g26400), .I2 (g17389));
AN2X1 gate9970(.O (g34528), .I1 (g34305), .I2 (g19617));
AN2X1 gate9971(.O (g17692), .I1 (g1124), .I2 (g13307));
AN2X1 gate9972(.O (g18130), .I1 (g528), .I2 (g16971));
AN2X1 gate9973(.O (g34696), .I1 (g34531), .I2 (g20004));
AN2X1 gate9974(.O (g18193), .I1 (g837), .I2 (g17821));
AN2X1 gate9975(.O (g22013), .I1 (g5802), .I2 (g21562));
AN2X1 gate9976(.O (g32157), .I1 (g31646), .I2 (g30021));
AN2X1 gate9977(.O (g34393), .I1 (g34189), .I2 (g21304));
AN2X1 gate9978(.O (g26259), .I1 (g24430), .I2 (g25232));
AN3X1 gate9979(.O (I24508), .I1 (g9434), .I2 (g9672), .I3 (g5401));
AN2X1 gate9980(.O (g18362), .I1 (g1834), .I2 (g17955));
AN2X1 gate9981(.O (g23218), .I1 (g20200), .I2 (g16530));
AN2X1 gate9982(.O (g29861), .I1 (g28390), .I2 (g23313));
AN2X1 gate9983(.O (g29573), .I1 (g1752), .I2 (g28892));
AN2X1 gate9984(.O (g33071), .I1 (g31591), .I2 (g32404));
AN2X1 gate9985(.O (g21837), .I1 (g3719), .I2 (g20453));
AN2X1 gate9986(.O (g34764), .I1 (g34691), .I2 (g20009));
AN2X1 gate9987(.O (g22329), .I1 (g11940), .I2 (g20329));
AN2X1 gate9988(.O (g10883), .I1 (g3355), .I2 (g9061));
AN2X1 gate9989(.O (g18165), .I1 (g650), .I2 (g17433));
AN2X1 gate9990(.O (g23837), .I1 (g21160), .I2 (g10804));
AN2X1 gate9991(.O (g18523), .I1 (g2675), .I2 (g15509));
AN2X1 gate9992(.O (g26087), .I1 (g5475), .I2 (g25072));
AN2X1 gate9993(.O (g27034), .I1 (g26328), .I2 (g8609));
AN2X1 gate9994(.O (g13306), .I1 (g441), .I2 (g11048));
AN2X1 gate9995(.O (g31776), .I1 (g21329), .I2 (g29385));
AN2X1 gate9996(.O (g34365), .I1 (g34149), .I2 (g20451));
AN2X1 gate9997(.O (g26258), .I1 (g12875), .I2 (g25231));
AN2X1 gate9998(.O (g19651), .I1 (g1111), .I2 (g16119));
AN2X1 gate9999(.O (g33785), .I1 (g33100), .I2 (g20550));
AN2X1 gate10000(.O (g29926), .I1 (g1604), .I2 (g28736));
AN2X1 gate10001(.O (g34869), .I1 (g34816), .I2 (g19869));
AN2X1 gate10002(.O (g28139), .I1 (g27337), .I2 (g26054));
AN2X1 gate10003(.O (g22005), .I1 (g5759), .I2 (g21562));
AN2X1 gate10004(.O (g31147), .I1 (g12286), .I2 (g30054));
AN2X1 gate10005(.O (g28653), .I1 (g7544), .I2 (g27014));
AN2X1 gate10006(.O (g13038), .I1 (g8509), .I2 (g11034));
AN2X1 gate10007(.O (g27292), .I1 (g1714), .I2 (g26654));
AN2X1 gate10008(.O (g29612), .I1 (g27875), .I2 (g28633));
AN2X1 gate10009(.O (g24465), .I1 (g3827), .I2 (g23139));
AN3X1 gate10010(.O (g12641), .I1 (g10295), .I2 (g3171), .I3 (g3179));
AN2X1 gate10011(.O (g22538), .I1 (g14035), .I2 (g20248));
AN2X1 gate10012(.O (g27153), .I1 (g26055), .I2 (g16629));
AN2X1 gate10013(.O (g33355), .I1 (g32243), .I2 (g20769));
AN2X1 gate10014(.O (g29324), .I1 (g29078), .I2 (g18883));
AN2X1 gate10015(.O (g34868), .I1 (g34813), .I2 (g19866));
AN2X1 gate10016(.O (g7396), .I1 (g392), .I2 (g441));
AN2X1 gate10017(.O (g25031), .I1 (g20675), .I2 (g23432));
AN2X1 gate10018(.O (g30161), .I1 (g28614), .I2 (g21275));
AN2X1 gate10019(.O (g18475), .I1 (g12853), .I2 (g15426));
AN2X1 gate10020(.O (g33859), .I1 (g33426), .I2 (g10531));
AN4X1 gate10021(.O (g26244), .I1 (g24688), .I2 (g8812), .I3 (g10658), .I4 (g8757));
AN2X1 gate10022(.O (g29534), .I1 (g28965), .I2 (g22457));
AN2X1 gate10023(.O (g33370), .I1 (g32279), .I2 (g21139));
AN2X1 gate10024(.O (g24983), .I1 (g23217), .I2 (g20238));
AN2X1 gate10025(.O (g27409), .I1 (g26519), .I2 (g17524));
AN2X1 gate10026(.O (g16855), .I1 (g4392), .I2 (g13107));
AN2X1 gate10027(.O (g18727), .I1 (g4931), .I2 (g16077));
AN2X1 gate10028(.O (g28415), .I1 (g27250), .I2 (g19963));
AN2X1 gate10029(.O (g24684), .I1 (g11769), .I2 (g22989));
AN2X1 gate10030(.O (g28333), .I1 (g27239), .I2 (g19787));
AN2X1 gate10031(.O (g33858), .I1 (g33268), .I2 (g20448));
AN2X1 gate10032(.O (g34709), .I1 (g34549), .I2 (g17242));
AN2X1 gate10033(.O (g18222), .I1 (g1024), .I2 (g16100));
AN2X1 gate10034(.O (g10501), .I1 (g1233), .I2 (g9007));
AN2X1 gate10035(.O (g16870), .I1 (g6625), .I2 (g14905));
AN2X1 gate10036(.O (g27136), .I1 (g26026), .I2 (g16605));
AN2X1 gate10037(.O (g27408), .I1 (g26519), .I2 (g17523));
AN4X1 gate10038(.O (g27635), .I1 (g23032), .I2 (g26281), .I3 (g26424), .I4 (g24996));
AN2X1 gate10039(.O (g21915), .I1 (g5080), .I2 (g21468));
AN2X1 gate10040(.O (g30225), .I1 (g28705), .I2 (g23897));
AN2X1 gate10041(.O (g31151), .I1 (g10037), .I2 (g30065));
AN2X1 gate10042(.O (g18437), .I1 (g2241), .I2 (g18008));
AN2X1 gate10043(.O (g24142), .I1 (g17700), .I2 (g21657));
AN4X1 gate10044(.O (I31001), .I1 (g29385), .I2 (g32456), .I3 (g32457), .I4 (g32458));
AN2X1 gate10045(.O (g31996), .I1 (g31779), .I2 (g18979));
AN2X1 gate10046(.O (g34225), .I1 (g33744), .I2 (g22942));
AN4X1 gate10047(.O (I31077), .I1 (g32566), .I2 (g32567), .I3 (g32568), .I4 (g32569));
AN2X1 gate10048(.O (g26602), .I1 (g7487), .I2 (g24453));
AN2X1 gate10049(.O (g30258), .I1 (g28751), .I2 (g23953));
AN2X1 gate10050(.O (g11937), .I1 (g1936), .I2 (g7362));
AN2X1 gate10051(.O (g15860), .I1 (g3889), .I2 (g14160));
AN3X1 gate10052(.O (g34087), .I1 (g33766), .I2 (g9104), .I3 (g18957));
AN2X1 gate10053(.O (g23201), .I1 (g14027), .I2 (g20040));
AN2X1 gate10054(.O (g33844), .I1 (g33257), .I2 (g20327));
AN2X1 gate10055(.O (g33367), .I1 (g32271), .I2 (g21053));
AN4X1 gate10056(.O (I31256), .I1 (g31021), .I2 (g31841), .I3 (g32824), .I4 (g32825));
AN2X1 gate10057(.O (g18703), .I1 (g4776), .I2 (g16782));
AN2X1 gate10058(.O (g22100), .I1 (g6466), .I2 (g18833));
AN2X1 gate10059(.O (g18347), .I1 (g1756), .I2 (g17955));
AN2X1 gate10060(.O (g19717), .I1 (g6527), .I2 (g17122));
AN2X1 gate10061(.O (g14438), .I1 (g1087), .I2 (g10726));
AN2X1 gate10062(.O (g30043), .I1 (g29106), .I2 (g9392));
AN2X1 gate10063(.O (g18253), .I1 (g1211), .I2 (g16897));
AN2X1 gate10064(.O (g25132), .I1 (g10497), .I2 (g23528));
AN2X1 gate10065(.O (g30244), .I1 (g28732), .I2 (g23930));
AN4X1 gate10066(.O (g26171), .I1 (g25357), .I2 (g6856), .I3 (g11709), .I4 (g11686));
AN2X1 gate10067(.O (g15700), .I1 (g3089), .I2 (g13483));
AN3X1 gate10068(.O (I24051), .I1 (g3380), .I2 (g3385), .I3 (g8492));
AN2X1 gate10069(.O (g18600), .I1 (g3111), .I2 (g16987));
AN2X1 gate10070(.O (g20193), .I1 (g15578), .I2 (g17264));
AN2X1 gate10071(.O (g18781), .I1 (g5831), .I2 (g18065));
AN2X1 gate10072(.O (g28585), .I1 (g27063), .I2 (g10530));
AN2X1 gate10073(.O (g24193), .I1 (g336), .I2 (g22722));
AN4X1 gate10074(.O (g28484), .I1 (g27187), .I2 (g10290), .I3 (g21163), .I4 (I26972));
AN2X1 gate10075(.O (g33420), .I1 (g32373), .I2 (g21454));
AN2X1 gate10076(.O (g30069), .I1 (g29175), .I2 (g12708));
AN2X1 gate10077(.O (g29766), .I1 (g28316), .I2 (g23235));
AN2X1 gate10078(.O (g18236), .I1 (g15065), .I2 (g16326));
AN2X1 gate10079(.O (g21782), .I1 (g3416), .I2 (g20391));
AN2X1 gate10080(.O (g17771), .I1 (g13288), .I2 (g13190));
AN2X1 gate10081(.O (g20165), .I1 (g5156), .I2 (g17733));
AN2X1 gate10082(.O (g34069), .I1 (g8774), .I2 (g33797));
AN2X1 gate10083(.O (g21984), .I1 (g5563), .I2 (g19074));
AN4X1 gate10084(.O (I31102), .I1 (g32603), .I2 (g32604), .I3 (g32605), .I4 (g32606));
AN4X1 gate10085(.O (g26994), .I1 (g23032), .I2 (g26226), .I3 (g26424), .I4 (g25557));
AN4X1 gate10086(.O (g27474), .I1 (g8038), .I2 (g26314), .I3 (g518), .I4 (g504));
AN2X1 gate10087(.O (g28554), .I1 (g27426), .I2 (g20372));
AN4X1 gate10088(.O (I31157), .I1 (g32682), .I2 (g32683), .I3 (g32684), .I4 (g32685));
AN2X1 gate10089(.O (g18351), .I1 (g1760), .I2 (g17955));
AN2X1 gate10090(.O (g18372), .I1 (g1886), .I2 (g15171));
AN2X1 gate10091(.O (g24523), .I1 (g22318), .I2 (g19468));
AN2X1 gate10092(.O (g32314), .I1 (g31304), .I2 (g23516));
AN2X1 gate10093(.O (g29871), .I1 (g28400), .I2 (g23332));
AN2X1 gate10094(.O (g33446), .I1 (g32385), .I2 (g21607));
AN4X1 gate10095(.O (g27711), .I1 (g22369), .I2 (g25193), .I3 (g26424), .I4 (g26166));
AN2X1 gate10096(.O (g16707), .I1 (g6641), .I2 (g15033));
AN2X1 gate10097(.O (g21419), .I1 (g16681), .I2 (g13595));
AN2X1 gate10098(.O (g32287), .I1 (g2823), .I2 (g30578));
AN2X1 gate10099(.O (g34774), .I1 (g34695), .I2 (g20180));
AN2X1 gate10100(.O (g18175), .I1 (g744), .I2 (g17328));
AN2X1 gate10101(.O (g18821), .I1 (g15168), .I2 (g15680));
AN2X1 gate10102(.O (g34955), .I1 (g34931), .I2 (g34320));
AN2X1 gate10103(.O (g27327), .I1 (g2116), .I2 (g26732));
AN2X1 gate10104(.O (g34375), .I1 (g13077), .I2 (g34049));
AN2X1 gate10105(.O (g16202), .I1 (g86), .I2 (g14197));
AN2X1 gate10106(.O (g28312), .I1 (g27828), .I2 (g26608));
AN2X1 gate10107(.O (g28200), .I1 (g27652), .I2 (g11383));
AN2X1 gate10108(.O (g32307), .I1 (g31291), .I2 (g23500));
AN2X1 gate10109(.O (g14566), .I1 (g10566), .I2 (g10551));
AN2X1 gate10110(.O (g32085), .I1 (g27253), .I2 (g31021));
AN4X1 gate10111(.O (I31066), .I1 (g31070), .I2 (g31807), .I3 (g32550), .I4 (g32551));
AN2X1 gate10112(.O (g29360), .I1 (g27364), .I2 (g28294));
AN2X1 gate10113(.O (g21822), .I1 (g3727), .I2 (g20453));
AN2X1 gate10114(.O (g22515), .I1 (g12981), .I2 (g19395));
AN4X1 gate10115(.O (I31231), .I1 (g31376), .I2 (g31836), .I3 (g32789), .I4 (g32790));
AN2X1 gate10116(.O (g22991), .I1 (g645), .I2 (g20248));
AN2X1 gate10117(.O (g27537), .I1 (g26549), .I2 (g17742));
AN2X1 gate10118(.O (g28115), .I1 (g27354), .I2 (g22759));
AN2X1 gate10119(.O (g31540), .I1 (g29904), .I2 (g23548));
AN2X1 gate10120(.O (g25087), .I1 (g17307), .I2 (g23489));
AN2X1 gate10121(.O (g32054), .I1 (g10890), .I2 (g30735));
AN2X1 gate10122(.O (g24475), .I1 (g3831), .I2 (g23139));
AN2X1 gate10123(.O (g7685), .I1 (g4382), .I2 (g4375));
AN2X1 gate10124(.O (g18264), .I1 (g1263), .I2 (g16000));
AN2X1 gate10125(.O (g18790), .I1 (g6040), .I2 (g15634));
AN2X1 gate10126(.O (g18137), .I1 (g538), .I2 (g17249));
AN4X1 gate10127(.O (I27513), .I1 (g19984), .I2 (g24089), .I3 (g24090), .I4 (g28034));
AN2X1 gate10128(.O (g18516), .I1 (g2638), .I2 (g15509));
AN2X1 gate10129(.O (g34337), .I1 (g34095), .I2 (g19881));
AN2X1 gate10130(.O (g24727), .I1 (g13300), .I2 (g23016));
AN2X1 gate10131(.O (g34171), .I1 (g33925), .I2 (g24360));
AN2X1 gate10132(.O (g16590), .I1 (g5236), .I2 (g14683));
AN2X1 gate10133(.O (g24222), .I1 (g262), .I2 (g22594));
AN2X1 gate10134(.O (g16986), .I1 (g246), .I2 (g13142));
AN2X1 gate10135(.O (g27303), .I1 (g11996), .I2 (g26681));
AN2X1 gate10136(.O (g11223), .I1 (g8281), .I2 (g8505));
AN2X1 gate10137(.O (g25043), .I1 (g20733), .I2 (g23447));
AN2X1 gate10138(.O (g32269), .I1 (g31253), .I2 (g20443));
AN2X1 gate10139(.O (g21853), .I1 (g3917), .I2 (g21070));
AN4X1 gate10140(.O (g28799), .I1 (g21434), .I2 (g26424), .I3 (g25348), .I4 (g27445));
AN2X1 gate10141(.O (g26079), .I1 (g6199), .I2 (g25060));
AN2X1 gate10142(.O (g34967), .I1 (g34951), .I2 (g23189));
AN2X1 gate10143(.O (g28813), .I1 (g4104), .I2 (g27038));
AN2X1 gate10144(.O (g29629), .I1 (g28211), .I2 (g19779));
AN2X1 gate10145(.O (g32341), .I1 (g31472), .I2 (g23610));
AN2X1 gate10146(.O (g31281), .I1 (g30106), .I2 (g27742));
AN2X1 gate10147(.O (g15870), .I1 (g3231), .I2 (g13948));
AN2X1 gate10148(.O (g26078), .I1 (g5128), .I2 (g25055));
AN2X1 gate10149(.O (g32156), .I1 (g31639), .I2 (g30018));
AN2X1 gate10150(.O (g25069), .I1 (g23296), .I2 (g20535));
AN2X1 gate10151(.O (g24703), .I1 (g17592), .I2 (g22369));
AN2X1 gate10152(.O (g31301), .I1 (g30170), .I2 (g27907));
AN2X1 gate10153(.O (g18209), .I1 (g921), .I2 (g15938));
AN2X1 gate10154(.O (g29628), .I1 (g27924), .I2 (g28648));
AN2X1 gate10155(.O (g33902), .I1 (g33085), .I2 (g13202));
AN2X1 gate10156(.O (g21836), .I1 (g3805), .I2 (g20453));
AN2X1 gate10157(.O (g31120), .I1 (g1700), .I2 (g29976));
AN2X1 gate10158(.O (g32180), .I1 (g2791), .I2 (g31638));
AN2X1 gate10159(.O (g23836), .I1 (g4129), .I2 (g19495));
AN2X1 gate10160(.O (g26086), .I1 (g9672), .I2 (g25255));
AN2X1 gate10161(.O (g28674), .I1 (g27569), .I2 (g20629));
AN2X1 gate10162(.O (g13321), .I1 (g847), .I2 (g11048));
AN2X1 gate10163(.O (g25068), .I1 (g17574), .I2 (g23477));
AN2X1 gate10164(.O (g25955), .I1 (g24720), .I2 (g19580));
AN2X1 gate10165(.O (g30919), .I1 (g29898), .I2 (g23286));
AN2X1 gate10166(.O (g18208), .I1 (g930), .I2 (g15938));
AN2X1 gate10167(.O (g16801), .I1 (g5120), .I2 (g14238));
AN2X1 gate10168(.O (g16735), .I1 (g6235), .I2 (g15027));
AN2X1 gate10169(.O (g23401), .I1 (g7262), .I2 (g21460));
AN2X1 gate10170(.O (g25879), .I1 (g11135), .I2 (g24683));
AN2X1 gate10171(.O (g24600), .I1 (g22591), .I2 (g19652));
AN2X1 gate10172(.O (g25970), .I1 (g1792), .I2 (g24991));
AN2X1 gate10173(.O (g31146), .I1 (g12285), .I2 (g30053));
AN2X1 gate10174(.O (g30010), .I1 (g29035), .I2 (g9274));
AN2X1 gate10175(.O (g30918), .I1 (g8681), .I2 (g29707));
AN2X1 gate10176(.O (g32335), .I1 (g6199), .I2 (g31566));
AN4X1 gate10177(.O (g11178), .I1 (g6682), .I2 (g7097), .I3 (g6668), .I4 (g10061));
AN2X1 gate10178(.O (g11740), .I1 (g8769), .I2 (g703));
AN2X1 gate10179(.O (g18542), .I1 (g2787), .I2 (g15277));
AN3X1 gate10180(.O (I18803), .I1 (g13156), .I2 (g11450), .I3 (g6756));
AN2X1 gate10181(.O (g18453), .I1 (g2315), .I2 (g15224));
AN2X1 gate10182(.O (g29591), .I1 (g28552), .I2 (g11346));
AN2X1 gate10183(.O (g29785), .I1 (g28332), .I2 (g23248));
AN2X1 gate10184(.O (g31290), .I1 (g29734), .I2 (g23335));
AN2X1 gate10185(.O (g22114), .I1 (g6565), .I2 (g19277));
AN2X1 gate10186(.O (g26159), .I1 (g2370), .I2 (g25137));
AN2X1 gate10187(.O (g26125), .I1 (g1894), .I2 (g25117));
AN2X1 gate10188(.O (g21864), .I1 (g3961), .I2 (g21070));
AN2X1 gate10189(.O (g34079), .I1 (g33703), .I2 (g19532));
AN2X1 gate10190(.O (g22082), .I1 (g6283), .I2 (g19210));
AN2X1 gate10191(.O (g27390), .I1 (g26549), .I2 (g17504));
AN2X1 gate10192(.O (g18726), .I1 (g4927), .I2 (g16077));
AN4X1 gate10193(.O (g26977), .I1 (g23032), .I2 (g26261), .I3 (g26424), .I4 (g25550));
AN2X1 gate10194(.O (g30599), .I1 (g18911), .I2 (g29863));
AN2X1 gate10195(.O (g22107), .I1 (g6411), .I2 (g18833));
AN2X1 gate10196(.O (g30078), .I1 (g28526), .I2 (g20667));
AN2X1 gate10197(.O (g21749), .I1 (g3155), .I2 (g20785));
AN2X1 gate10198(.O (g26158), .I1 (g2255), .I2 (g25432));
AN4X1 gate10199(.O (g17725), .I1 (g11547), .I2 (g11592), .I3 (g6789), .I4 (I18716));
AN2X1 gate10200(.O (g26783), .I1 (g25037), .I2 (g21048));
AN4X1 gate10201(.O (I31287), .I1 (g32870), .I2 (g32871), .I3 (g32872), .I4 (g32873));
AN2X1 gate10202(.O (g18614), .I1 (g3343), .I2 (g17200));
AN2X1 gate10203(.O (g28692), .I1 (g27578), .I2 (g20661));
AN4X1 gate10204(.O (g28761), .I1 (g21434), .I2 (g26424), .I3 (g25299), .I4 (g27416));
AN2X1 gate10205(.O (g34078), .I1 (g33699), .I2 (g19531));
AN2X1 gate10206(.O (g18436), .I1 (g2227), .I2 (g18008));
AN2X1 gate10207(.O (g25967), .I1 (g9373), .I2 (g24986));
AN2X1 gate10208(.O (g30598), .I1 (g18898), .I2 (g29862));
AN2X1 gate10209(.O (g14585), .I1 (g1141), .I2 (g10905));
AN2X1 gate10210(.O (g29859), .I1 (g28388), .I2 (g23307));
AN4X1 gate10211(.O (I31307), .I1 (g32898), .I2 (g32899), .I3 (g32900), .I4 (g32901));
AN4X1 gate10212(.O (I31076), .I1 (g30614), .I2 (g31809), .I3 (g32564), .I4 (g32565));
AN2X1 gate10213(.O (g30086), .I1 (g28536), .I2 (g20704));
AN2X1 gate10214(.O (g21748), .I1 (g15089), .I2 (g20785));
AN2X1 gate10215(.O (g15707), .I1 (g4082), .I2 (g13506));
AN2X1 gate10216(.O (g15819), .I1 (g3251), .I2 (g14101));
AN2X1 gate10217(.O (g18607), .I1 (g3139), .I2 (g16987));
AN3X1 gate10218(.O (g34086), .I1 (g20114), .I2 (g33766), .I3 (g9104));
AN2X1 gate10219(.O (g18320), .I1 (g1616), .I2 (g17873));
AN2X1 gate10220(.O (g24790), .I1 (g7074), .I2 (g23681));
AN2X1 gate10221(.O (g21276), .I1 (g10157), .I2 (g17625));
AN2X1 gate10222(.O (g21285), .I1 (g7857), .I2 (g16027));
AN2X1 gate10223(.O (g26295), .I1 (g13070), .I2 (g25266));
AN2X1 gate10224(.O (g29858), .I1 (g28387), .I2 (g23306));
AN2X1 gate10225(.O (g21704), .I1 (g164), .I2 (g20283));
AN2X1 gate10226(.O (g18274), .I1 (g1311), .I2 (g16031));
AN2X1 gate10227(.O (g22849), .I1 (g1227), .I2 (g19653));
AN2X1 gate10228(.O (g33366), .I1 (g32268), .I2 (g21010));
AN2X1 gate10229(.O (g27522), .I1 (g26549), .I2 (g17717));
AN2X1 gate10230(.O (g26823), .I1 (g24401), .I2 (g13106));
AN2X1 gate10231(.O (g15818), .I1 (g3941), .I2 (g14082));
AN2X1 gate10232(.O (g18530), .I1 (g2715), .I2 (g15277));
AN3X1 gate10233(.O (g25459), .I1 (g6058), .I2 (g23844), .I3 (I24582));
AN2X1 gate10234(.O (g18593), .I1 (g2999), .I2 (g16349));
AN2X1 gate10235(.O (g18346), .I1 (g1752), .I2 (g17955));
AN2X1 gate10236(.O (g19716), .I1 (g12100), .I2 (g17121));
AN2X1 gate10237(.O (g21809), .I1 (g3574), .I2 (g20924));
AN2X1 gate10238(.O (g23254), .I1 (g20056), .I2 (g20110));
AN2X1 gate10239(.O (g28214), .I1 (g27731), .I2 (g26625));
AN2X1 gate10240(.O (g15111), .I1 (g4281), .I2 (g14454));
AN2X1 gate10241(.O (g22848), .I1 (g19449), .I2 (g19649));
AN2X1 gate10242(.O (g18122), .I1 (g15052), .I2 (g17015));
AN2X1 gate10243(.O (g23900), .I1 (g1129), .I2 (g19408));
AN2X1 gate10244(.O (g34322), .I1 (g14188), .I2 (g34174));
AN4X1 gate10245(.O (g14608), .I1 (g12638), .I2 (g12476), .I3 (g12429), .I4 (I16721));
AN2X1 gate10246(.O (g15978), .I1 (g246), .I2 (g14032));
AN2X1 gate10247(.O (g18565), .I1 (g2852), .I2 (g16349));
AN2X1 gate10248(.O (g26336), .I1 (g10307), .I2 (g25480));
AN2X1 gate10249(.O (g30125), .I1 (g28581), .I2 (g21056));
AN2X1 gate10250(.O (g18464), .I1 (g2370), .I2 (g15224));
AN2X1 gate10251(.O (g21808), .I1 (g3570), .I2 (g20924));
AN2X1 gate10252(.O (g29844), .I1 (g28374), .I2 (g23290));
AN2X1 gate10253(.O (g34532), .I1 (g34314), .I2 (g19710));
AN2X1 gate10254(.O (g15590), .I1 (g3139), .I2 (g13530));
AN2X1 gate10255(.O (g29367), .I1 (g8575), .I2 (g28325));
AN2X1 gate10256(.O (g28539), .I1 (g27187), .I2 (g12762));
AN2X1 gate10257(.O (g10921), .I1 (g1548), .I2 (g8685));
AN2X1 gate10258(.O (g27483), .I1 (g26488), .I2 (g17642));
AN2X1 gate10259(.O (g30158), .I1 (g28613), .I2 (g21274));
AN2X1 gate10260(.O (g33403), .I1 (g32352), .I2 (g21396));
AN2X1 gate10261(.O (g24422), .I1 (g4771), .I2 (g22896));
AN4X1 gate10262(.O (I31341), .I1 (g31710), .I2 (g31856), .I3 (g32947), .I4 (g32948));
AN2X1 gate10263(.O (g32278), .I1 (g2811), .I2 (g30572));
AN2X1 gate10264(.O (g27553), .I1 (g26293), .I2 (g23353));
AN2X1 gate10265(.O (g18641), .I1 (g3841), .I2 (g17096));
AN2X1 gate10266(.O (g18797), .I1 (g6173), .I2 (g15348));
AN2X1 gate10267(.O (g25079), .I1 (g21011), .I2 (g23483));
AN4X1 gate10268(.O (I31156), .I1 (g31070), .I2 (g31823), .I3 (g32680), .I4 (g32681));
AN2X1 gate10269(.O (g18292), .I1 (g1472), .I2 (g16449));
AN2X1 gate10270(.O (g16706), .I1 (g6621), .I2 (g14868));
AN2X1 gate10271(.O (g31226), .I1 (g30282), .I2 (g25218));
AN2X1 gate10272(.O (g32286), .I1 (g31658), .I2 (g29312));
AN2X1 gate10273(.O (g34561), .I1 (g34368), .I2 (g17410));
AN2X1 gate10274(.O (g16597), .I1 (g6263), .I2 (g15021));
AN2X1 gate10275(.O (g18153), .I1 (g626), .I2 (g17533));
AN2X1 gate10276(.O (g27326), .I1 (g12048), .I2 (g26731));
AN2X1 gate10277(.O (g25078), .I1 (g23298), .I2 (g20538));
AN2X1 gate10278(.O (g31481), .I1 (g29768), .I2 (g23417));
AN2X1 gate10279(.O (g32039), .I1 (g31476), .I2 (g20070));
AN2X1 gate10280(.O (g33715), .I1 (g33135), .I2 (g19416));
AN2X1 gate10281(.O (g32306), .I1 (g31289), .I2 (g23499));
AN2X1 gate10282(.O (g34295), .I1 (g34057), .I2 (g19370));
AN3X1 gate10283(.O (g33481), .I1 (g32607), .I2 (I31101), .I3 (I31102));
AN2X1 gate10284(.O (g22135), .I1 (g6657), .I2 (g19277));
AN2X1 gate10285(.O (g27536), .I1 (g26519), .I2 (g17738));
AN2X1 gate10286(.O (g18409), .I1 (g2084), .I2 (g15373));
AN4X1 gate10287(.O (g27040), .I1 (g7812), .I2 (g6565), .I3 (g6573), .I4 (g26226));
AN2X1 gate10288(.O (g25086), .I1 (g13941), .I2 (g23488));
AN2X1 gate10289(.O (g21733), .I1 (g3034), .I2 (g20330));
AN3X1 gate10290(.O (g10674), .I1 (g6841), .I2 (g10200), .I3 (g2130));
AN2X1 gate10291(.O (g18136), .I1 (g550), .I2 (g17249));
AN2X1 gate10292(.O (g18408), .I1 (g2070), .I2 (g15373));
AN2X1 gate10293(.O (g18635), .I1 (g3808), .I2 (g17096));
AN2X1 gate10294(.O (g24726), .I1 (g15965), .I2 (g23015));
AN2X1 gate10295(.O (g27252), .I1 (g26733), .I2 (g26703));
AN2X1 gate10296(.O (g24913), .I1 (g4821), .I2 (g23908));
AN2X1 gate10297(.O (g21874), .I1 (g4112), .I2 (g19801));
AN2X1 gate10298(.O (g25817), .I1 (g24807), .I2 (g21163));
AN2X1 gate10299(.O (g32187), .I1 (g30672), .I2 (g25287));
AN2X1 gate10300(.O (g26289), .I1 (g2551), .I2 (g25400));
AN2X1 gate10301(.O (g24436), .I1 (g3125), .I2 (g23067));
AN2X1 gate10302(.O (g25159), .I1 (g4907), .I2 (g22908));
AN3X1 gate10303(.O (g10732), .I1 (g6850), .I2 (g2697), .I3 (g2689));
AN2X1 gate10304(.O (g22049), .I1 (g6082), .I2 (g21611));
AN2X1 gate10305(.O (g25125), .I1 (g20187), .I2 (g23520));
AN2X1 gate10306(.O (g27564), .I1 (g26305), .I2 (g23378));
AN2X1 gate10307(.O (g25901), .I1 (g24853), .I2 (g16290));
AN2X1 gate10308(.O (g26023), .I1 (g9528), .I2 (g25036));
AN4X1 gate10309(.O (I31131), .I1 (g31542), .I2 (g31819), .I3 (g32643), .I4 (g32644));
AN2X1 gate10310(.O (g34966), .I1 (g34950), .I2 (g23170));
AN2X1 gate10311(.O (g31490), .I1 (g29786), .I2 (g23429));
AN2X1 gate10312(.O (g10934), .I1 (g9197), .I2 (g7918));
AN2X1 gate10313(.O (g24607), .I1 (g5817), .I2 (g23666));
AN2X1 gate10314(.O (g25977), .I1 (g25236), .I2 (g20875));
AN2X1 gate10315(.O (g26288), .I1 (g2259), .I2 (g25309));
AN3X1 gate10316(.O (g33490), .I1 (g32672), .I2 (I31146), .I3 (I31147));
AN2X1 gate10317(.O (g19681), .I1 (g5835), .I2 (g17014));
AN2X1 gate10318(.O (g24320), .I1 (g6973), .I2 (g22228));
AN2X1 gate10319(.O (g28235), .I1 (g9467), .I2 (g27592));
AN2X1 gate10320(.O (g26571), .I1 (g10472), .I2 (g24386));
AN2X1 gate10321(.O (g23166), .I1 (g13959), .I2 (g19979));
AN2X1 gate10322(.O (g23009), .I1 (g20196), .I2 (g14219));
AN2X1 gate10323(.O (g22048), .I1 (g6052), .I2 (g21611));
AN2X1 gate10324(.O (g26308), .I1 (g6961), .I2 (g25289));
AN3X1 gate10325(.O (g29203), .I1 (g24095), .I2 (I27513), .I3 (I27514));
AN2X1 gate10326(.O (g18164), .I1 (g699), .I2 (g17433));
AN2X1 gate10327(.O (g28683), .I1 (g27876), .I2 (g20649));
AN2X1 gate10328(.O (g32143), .I1 (g31646), .I2 (g29967));
AN2X1 gate10329(.O (g31784), .I1 (g30176), .I2 (g24003));
AN2X1 gate10330(.O (g34364), .I1 (g34048), .I2 (g24366));
AN2X1 gate10331(.O (g33784), .I1 (g33107), .I2 (g20531));
AN2X1 gate10332(.O (g31376), .I1 (g24952), .I2 (g29814));
AN2X1 gate10333(.O (g31297), .I1 (g30144), .I2 (g27837));
AN2X1 gate10334(.O (g27183), .I1 (g26055), .I2 (g16658));
AN2X1 gate10335(.O (g33376), .I1 (g32294), .I2 (g21268));
AN2X1 gate10336(.O (g27673), .I1 (g25769), .I2 (g23541));
AN2X1 gate10337(.O (g22004), .I1 (g5742), .I2 (g21562));
AN2X1 gate10338(.O (g23008), .I1 (g1570), .I2 (g19783));
AN2X1 gate10339(.O (g33889), .I1 (g33303), .I2 (g20641));
AN4X1 gate10340(.O (g11123), .I1 (g5644), .I2 (g7028), .I3 (g5630), .I4 (g9864));
AN2X1 gate10341(.O (g24464), .I1 (g3480), .I2 (g23112));
AN3X1 gate10342(.O (I24027), .I1 (g3029), .I2 (g3034), .I3 (g8426));
AN2X1 gate10343(.O (g16885), .I1 (g6605), .I2 (g14950));
AN2X1 gate10344(.O (g32169), .I1 (g31014), .I2 (g23046));
AN2X1 gate10345(.O (g18575), .I1 (g2878), .I2 (g16349));
AN2X1 gate10346(.O (g18474), .I1 (g2287), .I2 (g15224));
AN2X1 gate10347(.O (g29902), .I1 (g28430), .I2 (g23377));
AN2X1 gate10348(.O (g30289), .I1 (g28884), .I2 (g24000));
AN2X1 gate10349(.O (g29377), .I1 (g28132), .I2 (g19387));
AN2X1 gate10350(.O (g13807), .I1 (g4504), .I2 (g10606));
AN2X1 gate10351(.O (g18711), .I1 (g15136), .I2 (g15915));
AN2X1 gate10352(.O (g32168), .I1 (g30597), .I2 (g25185));
AN2X1 gate10353(.O (g32410), .I1 (g4933), .I2 (g30997));
AN4X1 gate10354(.O (g28991), .I1 (g14438), .I2 (g25209), .I3 (g26424), .I4 (g27469));
AN2X1 gate10355(.O (g13974), .I1 (g6243), .I2 (g12578));
AN2X1 gate10356(.O (g18327), .I1 (g1636), .I2 (g17873));
AN2X1 gate10357(.O (g24797), .I1 (g22872), .I2 (g19960));
AN2X1 gate10358(.O (g30023), .I1 (g28508), .I2 (g20570));
AN2X1 gate10359(.O (g21712), .I1 (g294), .I2 (g20283));
AN3X1 gate10360(.O (I24482), .I1 (g9364), .I2 (g9607), .I3 (g5057));
AN2X1 gate10361(.O (g18109), .I1 (g437), .I2 (g17015));
AN2X1 gate10362(.O (g27508), .I1 (g26549), .I2 (g17684));
AN2X1 gate10363(.O (g16763), .I1 (g6239), .I2 (g14937));
AN2X1 gate10364(.O (g27634), .I1 (g26805), .I2 (g26793));
AN2X1 gate10365(.O (g34309), .I1 (g13947), .I2 (g34147));
AN2X1 gate10366(.O (g21914), .I1 (g5077), .I2 (g21468));
AN2X1 gate10367(.O (g24292), .I1 (g4443), .I2 (g22550));
AN2X1 gate10368(.O (g30224), .I1 (g28704), .I2 (g23896));
AN2X1 gate10369(.O (g18537), .I1 (g6856), .I2 (g15277));
AN4X1 gate10370(.O (I24710), .I1 (g24071), .I2 (g24072), .I3 (g24073), .I4 (g24074));
AN2X1 gate10371(.O (g34224), .I1 (g33736), .I2 (g22670));
AN3X1 gate10372(.O (g30308), .I1 (g29178), .I2 (g7004), .I3 (g5297));
AN2X1 gate10373(.O (g22106), .I1 (g6497), .I2 (g18833));
AN3X1 gate10374(.O (I24552), .I1 (g9733), .I2 (g9316), .I3 (g5747));
AN2X1 gate10375(.O (g29645), .I1 (g1714), .I2 (g29018));
AN3X1 gate10376(.O (I24003), .I1 (g8097), .I2 (g8334), .I3 (g3045));
AN4X1 gate10377(.O (g17613), .I1 (g11547), .I2 (g11592), .I3 (g11640), .I4 (I18568));
AN2X1 gate10378(.O (g34571), .I1 (g27225), .I2 (g34299));
AN2X1 gate10379(.O (g18108), .I1 (g433), .I2 (g17015));
AN2X1 gate10380(.O (g14207), .I1 (g8639), .I2 (g11793));
AN2X1 gate10381(.O (g21907), .I1 (g5033), .I2 (g21468));
AN4X1 gate10382(.O (I31286), .I1 (g30825), .I2 (g31846), .I3 (g32868), .I4 (g32869));
AN3X1 gate10383(.O (I13862), .I1 (g7232), .I2 (g7219), .I3 (g7258));
AN2X1 gate10384(.O (g15077), .I1 (g2138), .I2 (g12955));
AN2X1 gate10385(.O (g24409), .I1 (g3484), .I2 (g23112));
AN2X1 gate10386(.O (g25966), .I1 (g9364), .I2 (g24985));
AN4X1 gate10387(.O (I31306), .I1 (g30614), .I2 (g31850), .I3 (g32896), .I4 (g32897));
AN2X1 gate10388(.O (g13265), .I1 (g9018), .I2 (g11493));
AN2X1 gate10389(.O (g18283), .I1 (g1384), .I2 (g16136));
AN2X1 gate10390(.O (g15706), .I1 (g13296), .I2 (g13484));
AN2X1 gate10391(.O (g18606), .I1 (g3133), .I2 (g16987));
AN2X1 gate10392(.O (g18492), .I1 (g2523), .I2 (g15426));
AN2X1 gate10393(.O (g18303), .I1 (g1536), .I2 (g16489));
AN2X1 gate10394(.O (g24408), .I1 (g23989), .I2 (g18946));
AN2X1 gate10395(.O (g24635), .I1 (g19874), .I2 (g22883));
AN2X1 gate10396(.O (g34495), .I1 (g34274), .I2 (g19365));
AN2X1 gate10397(.O (g22033), .I1 (g5925), .I2 (g19147));
AN2X1 gate10398(.O (g27213), .I1 (g26026), .I2 (g16721));
AN2X1 gate10399(.O (g18750), .I1 (g15145), .I2 (g17847));
AN2X1 gate10400(.O (g31520), .I1 (g29879), .I2 (g23507));
AN4X1 gate10401(.O (I31187), .I1 (g32726), .I2 (g32727), .I3 (g32728), .I4 (g32729));
AN3X1 gate10402(.O (g33520), .I1 (g32888), .I2 (I31296), .I3 (I31297));
AN2X1 gate10403(.O (g18982), .I1 (g3835), .I2 (g16159));
AN2X1 gate10404(.O (g18381), .I1 (g1882), .I2 (g15171));
AN2X1 gate10405(.O (g34687), .I1 (g14181), .I2 (g34543));
AN2X1 gate10406(.O (g21941), .I1 (g5232), .I2 (g18997));
AN2X1 gate10407(.O (g26842), .I1 (g2894), .I2 (g24522));
AN3X1 gate10408(.O (I27429), .I1 (g25562), .I2 (g26424), .I3 (g22698));
AN2X1 gate10409(.O (g27452), .I1 (g26400), .I2 (g17600));
AN2X1 gate10410(.O (g21382), .I1 (g10086), .I2 (g17625));
AN2X1 gate10411(.O (g29632), .I1 (g28899), .I2 (g22417));
AN2X1 gate10412(.O (g31211), .I1 (g10156), .I2 (g30102));
AN4X1 gate10413(.O (g26195), .I1 (g25357), .I2 (g6856), .I3 (g11709), .I4 (g7558));
AN2X1 gate10414(.O (g34752), .I1 (g34675), .I2 (g19544));
AN2X1 gate10415(.O (g23675), .I1 (g19050), .I2 (g9104));
AN2X1 gate10416(.O (g18174), .I1 (g739), .I2 (g17328));
AN2X1 gate10417(.O (g27311), .I1 (g12431), .I2 (g26693));
AN2X1 gate10418(.O (g18796), .I1 (g6167), .I2 (g15348));
AN2X1 gate10419(.O (g28725), .I1 (g27596), .I2 (g20779));
AN2X1 gate10420(.O (g32084), .I1 (g10948), .I2 (g30825));
AN2X1 gate10421(.O (g32110), .I1 (g31639), .I2 (g29921));
AN2X1 gate10422(.O (g16596), .I1 (g5941), .I2 (g14892));
AN2X1 gate10423(.O (g28114), .I1 (g25869), .I2 (g27051));
AN2X1 gate10424(.O (g25571), .I1 (I24694), .I2 (I24695));
AN2X1 gate10425(.O (g33860), .I1 (g33270), .I2 (g20501));
AN2X1 gate10426(.O (g32321), .I1 (g27613), .I2 (g31376));
AN2X1 gate10427(.O (g16243), .I1 (g6483), .I2 (g14275));
AN2X1 gate10428(.O (g29661), .I1 (g1687), .I2 (g29015));
AN2X1 gate10429(.O (g29547), .I1 (g1748), .I2 (g28857));
AN2X1 gate10430(.O (g29895), .I1 (g2495), .I2 (g29170));
AN2X1 gate10431(.O (g28107), .I1 (g27970), .I2 (g18874));
AN2X1 gate10432(.O (g10683), .I1 (g7289), .I2 (g4438));
AN2X1 gate10433(.O (g32179), .I1 (g31748), .I2 (g27907));
AN2X1 gate10434(.O (g21935), .I1 (g5196), .I2 (g18997));
AN2X1 gate10435(.O (g18390), .I1 (g1978), .I2 (g15171));
AN2X1 gate10436(.O (g31497), .I1 (g20041), .I2 (g29930));
AN3X1 gate10437(.O (g33497), .I1 (g32723), .I2 (I31181), .I3 (I31182));
AN2X1 gate10438(.O (g20109), .I1 (g17954), .I2 (g17616));
AN2X1 gate10439(.O (g24327), .I1 (g4549), .I2 (g22228));
AN2X1 gate10440(.O (g21883), .I1 (g4141), .I2 (g19801));
AN2X1 gate10441(.O (g32178), .I1 (g31747), .I2 (g27886));
AN2X1 gate10442(.O (g15876), .I1 (g13512), .I2 (g13223));
AN2X1 gate10443(.O (g24537), .I1 (g22626), .I2 (g10851));
AN2X1 gate10444(.O (g11116), .I1 (g9960), .I2 (g6466));
AN2X1 gate10445(.O (g20108), .I1 (g15508), .I2 (g11048));
AN2X1 gate10446(.O (g34842), .I1 (g34762), .I2 (g20168));
AN2X1 gate10447(.O (g18192), .I1 (g817), .I2 (g17821));
AN2X1 gate10448(.O (g22012), .I1 (g5752), .I2 (g21562));
AN2X1 gate10449(.O (g26544), .I1 (g7446), .I2 (g24357));
AN4X1 gate10450(.O (I27504), .I1 (g24077), .I2 (g24078), .I3 (g24079), .I4 (g24080));
AN3X1 gate10451(.O (I18620), .I1 (g13156), .I2 (g11450), .I3 (g11498));
AN2X1 gate10452(.O (g25816), .I1 (g8164), .I2 (g24604));
AN2X1 gate10453(.O (g33700), .I1 (g33148), .I2 (g11012));
AN2X1 gate10454(.O (g33126), .I1 (g9044), .I2 (g32201));
AN2X1 gate10455(.O (g31987), .I1 (g31767), .I2 (g22198));
AN2X1 gate10456(.O (g29551), .I1 (g2173), .I2 (g28867));
AN2X1 gate10457(.O (g29572), .I1 (g1620), .I2 (g28885));
AN2X1 gate10458(.O (g26713), .I1 (g25447), .I2 (g20714));
AN4X1 gate10459(.O (I31217), .I1 (g32768), .I2 (g32769), .I3 (g32770), .I4 (g32771));
AN2X1 gate10460(.O (g34489), .I1 (g34421), .I2 (g19068));
AN2X1 gate10461(.O (g24283), .I1 (g4411), .I2 (g22550));
AN2X1 gate10462(.O (g18522), .I1 (g2671), .I2 (g15509));
AN2X1 gate10463(.O (g27350), .I1 (g10217), .I2 (g26803));
AN2X1 gate10464(.O (g18663), .I1 (g4311), .I2 (g17367));
AN2X1 gate10465(.O (g24606), .I1 (g5489), .I2 (g23630));
AN2X1 gate10466(.O (g25976), .I1 (g9443), .I2 (g25000));
AN2X1 gate10467(.O (g24303), .I1 (g4369), .I2 (g22228));
AN2X1 gate10468(.O (g16670), .I1 (g5953), .I2 (g14999));
AN2X1 gate10469(.O (g27820), .I1 (g7670), .I2 (g25932));
AN2X1 gate10470(.O (g34525), .I1 (g34297), .I2 (g19528));
AN4X1 gate10471(.O (g28141), .I1 (g10831), .I2 (g11797), .I3 (g11261), .I4 (g27163));
AN2X1 gate10472(.O (g34488), .I1 (g34417), .I2 (g18988));
AN2X1 gate10473(.O (g28652), .I1 (g27282), .I2 (g10288));
AN2X1 gate10474(.O (g13493), .I1 (g9880), .I2 (g11866));
AN3X1 gate10475(.O (g25374), .I1 (g5366), .I2 (g23789), .I3 (I24527));
AN2X1 gate10476(.O (g31943), .I1 (g4717), .I2 (g30614));
AN3X1 gate10477(.O (I24505), .I1 (g9607), .I2 (g9229), .I3 (g5057));
AN2X1 gate10478(.O (g21729), .I1 (g3021), .I2 (g20330));
AN2X1 gate10479(.O (g26610), .I1 (g14198), .I2 (g24405));
AN2X1 gate10480(.O (g33339), .I1 (g32221), .I2 (g20634));
AN2X1 gate10481(.O (g33943), .I1 (g33384), .I2 (g21609));
AN2X1 gate10482(.O (g31296), .I1 (g30119), .I2 (g27779));
AN2X1 gate10483(.O (g34558), .I1 (g34353), .I2 (g20578));
AN2X1 gate10484(.O (g16734), .I1 (g5961), .I2 (g14735));
AN2X1 gate10485(.O (g23577), .I1 (g19444), .I2 (g13033));
AN2X1 gate10486(.O (g18483), .I1 (g2453), .I2 (g15426));
AN2X1 gate10487(.O (g24750), .I1 (g17662), .I2 (g22472));
AN2X1 gate10488(.O (g32334), .I1 (g31375), .I2 (g23568));
AN2X1 gate10489(.O (g21728), .I1 (g3010), .I2 (g20330));
AN2X1 gate10490(.O (g33338), .I1 (g32220), .I2 (g20633));
AN2X1 gate10491(.O (g28263), .I1 (g23747), .I2 (g27711));
AN2X1 gate10492(.O (g16930), .I1 (g239), .I2 (g13132));
AN2X1 gate10493(.O (g23439), .I1 (g13771), .I2 (g20452));
AN2X1 gate10494(.O (g11035), .I1 (g5441), .I2 (g9800));
AN2X1 gate10495(.O (g18553), .I1 (g2827), .I2 (g15277));
AN2X1 gate10496(.O (g13035), .I1 (g8497), .I2 (g11033));
AN2X1 gate10497(.O (g26270), .I1 (g1700), .I2 (g25275));
AN2X1 gate10498(.O (g31969), .I1 (g31189), .I2 (g22139));
AN2X1 gate10499(.O (g29784), .I1 (g28331), .I2 (g23247));
AN2X1 gate10500(.O (g26124), .I1 (g1811), .I2 (g25116));
AN2X1 gate10501(.O (g22920), .I1 (g19764), .I2 (g19719));
AN2X1 gate10502(.O (g16667), .I1 (g5268), .I2 (g14659));
AN2X1 gate10503(.O (g20174), .I1 (g5503), .I2 (g17754));
AN2X1 gate10504(.O (g29376), .I1 (g14002), .I2 (g28504));
AN2X1 gate10505(.O (g27413), .I1 (g26576), .I2 (g17530));
AN2X1 gate10506(.O (g34865), .I1 (g16540), .I2 (g34836));
AN2X1 gate10507(.O (g16965), .I1 (g269), .I2 (g13140));
AN2X1 gate10508(.O (g18949), .I1 (g10183), .I2 (g17625));
AN2X1 gate10509(.O (g31968), .I1 (g31757), .I2 (g22168));
AN2X1 gate10510(.O (g18326), .I1 (g1664), .I2 (g17873));
AN2X1 gate10511(.O (g24796), .I1 (g7097), .I2 (g23714));
AN2X1 gate10512(.O (g11142), .I1 (g6381), .I2 (g10207));
AN2X1 gate10513(.O (g27691), .I1 (g25778), .I2 (g23609));
AN4X1 gate10514(.O (g17724), .I1 (g11547), .I2 (g11592), .I3 (g11640), .I4 (I18713));
AN2X1 gate10515(.O (g29354), .I1 (g4961), .I2 (g28421));
AN4X1 gate10516(.O (I27533), .I1 (g21143), .I2 (g24125), .I3 (g24126), .I4 (g24127));
AN2X1 gate10517(.O (g18536), .I1 (g2748), .I2 (g15277));
AN2X1 gate10518(.O (g23349), .I1 (g13662), .I2 (g20182));
AN2X1 gate10519(.O (g22121), .I1 (g6593), .I2 (g19277));
AN2X1 gate10520(.O (g29888), .I1 (g28418), .I2 (g23352));
AN2X1 gate10521(.O (g33855), .I1 (g33265), .I2 (g20441));
AN2X1 gate10522(.O (g14206), .I1 (g8655), .I2 (g11790));
AN2X1 gate10523(.O (g21906), .I1 (g5022), .I2 (g21468));
AN2X1 gate10524(.O (g18702), .I1 (g15133), .I2 (g16856));
AN2X1 gate10525(.O (g21348), .I1 (g10121), .I2 (g17625));
AN2X1 gate10526(.O (g18757), .I1 (g5352), .I2 (g15595));
AN2X1 gate10527(.O (g31527), .I1 (g7553), .I2 (g29343));
AN2X1 gate10528(.O (g23083), .I1 (g16076), .I2 (g19878));
AN2X1 gate10529(.O (g23348), .I1 (g15570), .I2 (g21393));
AN2X1 gate10530(.O (g15076), .I1 (g2130), .I2 (g12955));
AN2X1 gate10531(.O (g33870), .I1 (g33280), .I2 (g20545));
AN2X1 gate10532(.O (g33411), .I1 (g32361), .I2 (g21410));
AN3X1 gate10533(.O (g33527), .I1 (g32939), .I2 (I31331), .I3 (I31332));
AN2X1 gate10534(.O (g26294), .I1 (g4245), .I2 (g25230));
AN4X1 gate10535(.O (I31321), .I1 (g31376), .I2 (g31852), .I3 (g32919), .I4 (g32920));
AN2X1 gate10536(.O (g16619), .I1 (g6629), .I2 (g14947));
AN2X1 gate10537(.O (g30042), .I1 (g29142), .I2 (g12601));
AN2X1 gate10538(.O (g18252), .I1 (g990), .I2 (g16897));
AN2X1 gate10539(.O (g18621), .I1 (g3476), .I2 (g17062));
AN2X1 gate10540(.O (g25559), .I1 (g13004), .I2 (g22649));
AN2X1 gate10541(.O (g30255), .I1 (g28748), .I2 (g23946));
AN3X1 gate10542(.O (g25488), .I1 (g6404), .I2 (g23865), .I3 (I24603));
AN4X1 gate10543(.O (g28833), .I1 (g21434), .I2 (g26424), .I3 (g25388), .I4 (g27469));
AN2X1 gate10544(.O (g16618), .I1 (g6609), .I2 (g15039));
AN2X1 gate10545(.O (g34679), .I1 (g14093), .I2 (g34539));
AN2X1 gate10546(.O (g18564), .I1 (g2844), .I2 (g16349));
AN2X1 gate10547(.O (g30188), .I1 (g28644), .I2 (g23841));
AN2X1 gate10548(.O (g24192), .I1 (g311), .I2 (g22722));
AN2X1 gate10549(.O (g30124), .I1 (g28580), .I2 (g21055));
AN2X1 gate10550(.O (g16279), .I1 (g4512), .I2 (g14424));
AN2X1 gate10551(.O (g34678), .I1 (g34490), .I2 (g19431));
AN2X1 gate10552(.O (g27020), .I1 (g4601), .I2 (g25852));
AN2X1 gate10553(.O (g31503), .I1 (g20041), .I2 (g29945));
AN3X1 gate10554(.O (I18716), .I1 (g13156), .I2 (g11450), .I3 (g6756));
AN4X1 gate10555(.O (I31186), .I1 (g31376), .I2 (g31828), .I3 (g32724), .I4 (g32725));
AN3X1 gate10556(.O (g33503), .I1 (g32765), .I2 (I31211), .I3 (I31212));
AN2X1 gate10557(.O (g24663), .I1 (g16621), .I2 (g22974));
AN2X1 gate10558(.O (g33867), .I1 (g33277), .I2 (g20529));
AN2X1 gate10559(.O (g17682), .I1 (g9742), .I2 (g14637));
AN2X1 gate10560(.O (g34686), .I1 (g34494), .I2 (g19494));
AN2X1 gate10561(.O (g13523), .I1 (g7046), .I2 (g12246));
AN2X1 gate10562(.O (g18183), .I1 (g781), .I2 (g17328));
AN2X1 gate10563(.O (g18673), .I1 (g4643), .I2 (g15758));
AN2X1 gate10564(.O (g25865), .I1 (g25545), .I2 (g18991));
AN4X1 gate10565(.O (g26218), .I1 (g25357), .I2 (g6856), .I3 (g7586), .I4 (g11686));
AN2X1 gate10566(.O (g18397), .I1 (g2004), .I2 (g15373));
AN2X1 gate10567(.O (g30030), .I1 (g29198), .I2 (g12347));
AN2X1 gate10568(.O (g30267), .I1 (g28776), .I2 (g23967));
AN3X1 gate10569(.O (g34093), .I1 (g20114), .I2 (g33755), .I3 (g9104));
AN2X1 gate10570(.O (g33450), .I1 (g32266), .I2 (g29737));
AN2X1 gate10571(.O (g22760), .I1 (g9360), .I2 (g20237));
AN2X1 gate10572(.O (g22134), .I1 (g6653), .I2 (g19277));
AN2X1 gate10573(.O (g27113), .I1 (g25997), .I2 (g16522));
AN2X1 gate10574(.O (g32242), .I1 (g31245), .I2 (g20324));
AN2X1 gate10575(.O (g18509), .I1 (g2587), .I2 (g15509));
AN2X1 gate10576(.O (g22029), .I1 (g5901), .I2 (g19147));
AN2X1 gate10577(.O (g31707), .I1 (g30081), .I2 (g23886));
AN2X1 gate10578(.O (g34065), .I1 (g33813), .I2 (g23148));
AN3X1 gate10579(.O (g33819), .I1 (g23088), .I2 (g33176), .I3 (g9104));
AN2X1 gate10580(.O (g33707), .I1 (g33174), .I2 (g13346));
AN2X1 gate10581(.O (g18933), .I1 (g16237), .I2 (g13597));
AN2X1 gate10582(.O (g33910), .I1 (g33134), .I2 (g7836));
AN2X1 gate10583(.O (g24553), .I1 (g22983), .I2 (g19539));
AN2X1 gate10584(.O (g26160), .I1 (g2453), .I2 (g25138));
AN2X1 gate10585(.O (g28273), .I1 (g27927), .I2 (g23729));
AN2X1 gate10586(.O (g7696), .I1 (g2955), .I2 (g2950));
AN2X1 gate10587(.O (g18508), .I1 (g2606), .I2 (g15509));
AN2X1 gate10588(.O (g22028), .I1 (g5893), .I2 (g19147));
AN2X1 gate10589(.O (g27302), .I1 (g1848), .I2 (g26680));
AN2X1 gate10590(.O (g18634), .I1 (g3813), .I2 (g17096));
AN2X1 gate10591(.O (g21333), .I1 (g1300), .I2 (g15740));
AN2X1 gate10592(.O (g23415), .I1 (g20077), .I2 (g20320));
AN2X1 gate10593(.O (g27357), .I1 (g26400), .I2 (g17414));
AN2X1 gate10594(.O (g25042), .I1 (g23262), .I2 (g20496));
AN2X1 gate10595(.O (g31496), .I1 (g2338), .I2 (g30312));
AN2X1 gate10596(.O (g33818), .I1 (g33236), .I2 (g20113));
AN2X1 gate10597(.O (g24949), .I1 (g23796), .I2 (g20751));
AN3X1 gate10598(.O (g33496), .I1 (g32714), .I2 (I31176), .I3 (I31177));
AN2X1 gate10599(.O (g19461), .I1 (g11708), .I2 (g16846));
AN2X1 gate10600(.O (g27105), .I1 (g26026), .I2 (g16511));
AN2X1 gate10601(.O (g24326), .I1 (g4552), .I2 (g22228));
AN2X1 gate10602(.O (g30219), .I1 (g28698), .I2 (g23887));
AN2X1 gate10603(.O (g17134), .I1 (g5619), .I2 (g14851));
AN2X1 gate10604(.O (g21852), .I1 (g3909), .I2 (g21070));
AN2X1 gate10605(.O (g15839), .I1 (g3929), .I2 (g13990));
AN2X1 gate10606(.O (g34875), .I1 (g34836), .I2 (g20073));
AN2X1 gate10607(.O (g28812), .I1 (g26972), .I2 (g13037));
AN2X1 gate10608(.O (g33111), .I1 (g24005), .I2 (g32421));
AN2X1 gate10609(.O (g34219), .I1 (g33736), .I2 (g22942));
AN2X1 gate10610(.O (g31070), .I1 (g29814), .I2 (g25985));
AN2X1 gate10611(.O (g19145), .I1 (g8450), .I2 (g16200));
AN2X1 gate10612(.O (g24536), .I1 (g19516), .I2 (g22635));
AN2X1 gate10613(.O (g29860), .I1 (g28389), .I2 (g23312));
AN2X1 gate10614(.O (g17506), .I1 (g9744), .I2 (g14505));
AN2X1 gate10615(.O (g25124), .I1 (g4917), .I2 (g22908));
AN2X1 gate10616(.O (g15694), .I1 (g457), .I2 (g13437));
AN2X1 gate10617(.O (g15838), .I1 (g3602), .I2 (g14133));
AN2X1 gate10618(.O (g21963), .I1 (g5436), .I2 (g21514));
AN2X1 gate10619(.O (g24702), .I1 (g17464), .I2 (g22342));
AN2X1 gate10620(.O (g34218), .I1 (g33744), .I2 (g22670));
AN2X1 gate10621(.O (g24757), .I1 (g7004), .I2 (g23563));
AN2X1 gate10622(.O (g31986), .I1 (g31766), .I2 (g22197));
AN2X1 gate10623(.O (g19736), .I1 (g12136), .I2 (g17136));
AN2X1 gate10624(.O (g24904), .I1 (g11761), .I2 (g23279));
AN2X1 gate10625(.O (g28234), .I1 (g27877), .I2 (g26686));
AN2X1 gate10626(.O (g32293), .I1 (g2827), .I2 (g30593));
AN4X1 gate10627(.O (I31216), .I1 (g30937), .I2 (g31834), .I3 (g32766), .I4 (g32767));
AN2X1 gate10628(.O (g25939), .I1 (g24583), .I2 (g19490));
AN2X1 gate10629(.O (g26277), .I1 (g2547), .I2 (g25400));
AN2X1 gate10630(.O (g18213), .I1 (g952), .I2 (g15979));
AN2X1 gate10631(.O (g32265), .I1 (g2799), .I2 (g30567));
AN2X1 gate10632(.O (g25030), .I1 (g23251), .I2 (g20432));
AN2X1 gate10633(.O (g25938), .I1 (g8997), .I2 (g24953));
AN2X1 gate10634(.O (g25093), .I1 (g12831), .I2 (g23493));
AN2X1 gate10635(.O (g31067), .I1 (g29484), .I2 (g22868));
AN2X1 gate10636(.O (g24564), .I1 (g23198), .I2 (g21163));
AN2X1 gate10637(.O (g29625), .I1 (g28514), .I2 (g14226));
AN3X1 gate10638(.O (g29987), .I1 (g29197), .I2 (g26424), .I3 (g22763));
AN2X1 gate10639(.O (g19393), .I1 (g691), .I2 (g16325));
AN2X1 gate10640(.O (g16884), .I1 (g6159), .I2 (g14321));
AN2X1 gate10641(.O (g18574), .I1 (g2882), .I2 (g16349));
AN2X1 gate10642(.O (g23484), .I1 (g20160), .I2 (g20541));
AN2X1 gate10643(.O (g18452), .I1 (g2311), .I2 (g15224));
AN2X1 gate10644(.O (g18205), .I1 (g904), .I2 (g15938));
AN2X1 gate10645(.O (g31150), .I1 (g1682), .I2 (g30063));
AN2X1 gate10646(.O (g23554), .I1 (g20390), .I2 (g13024));
AN4X1 gate10647(.O (I31117), .I1 (g32624), .I2 (g32625), .I3 (g32626), .I4 (g32627));
AN2X1 gate10648(.O (g18311), .I1 (g1554), .I2 (g16931));
AN2X1 gate10649(.O (g33801), .I1 (g33437), .I2 (g25327));
AN2X1 gate10650(.O (g24673), .I1 (g22659), .I2 (g19748));
AN2X1 gate10651(.O (g33735), .I1 (g33118), .I2 (g19553));
AN2X1 gate10652(.O (g33877), .I1 (g33287), .I2 (g20563));
AN3X1 gate10653(.O (I24582), .I1 (g9809), .I2 (g9397), .I3 (g6093));
AN2X1 gate10654(.O (g30915), .I1 (g29886), .I2 (g24778));
AN2X1 gate10655(.O (g29943), .I1 (g2165), .I2 (g28765));
AN2X1 gate10656(.O (g34470), .I1 (g7834), .I2 (g34325));
AN2X1 gate10657(.O (g16666), .I1 (g5200), .I2 (g14794));
AN2X1 gate10658(.O (g25875), .I1 (g8390), .I2 (g24809));
AN2X1 gate10659(.O (g31019), .I1 (g29481), .I2 (g22856));
AN3X1 gate10660(.O (I18765), .I1 (g13156), .I2 (g11450), .I3 (g11498));
AN2X1 gate10661(.O (g29644), .I1 (g28216), .I2 (g19794));
AN2X1 gate10662(.O (g29338), .I1 (g29145), .I2 (g22181));
AN2X1 gate10663(.O (g30277), .I1 (g28817), .I2 (g23987));
AN2X1 gate10664(.O (g13063), .I1 (g8567), .I2 (g10808));
AN2X1 gate10665(.O (g31018), .I1 (g29480), .I2 (g22855));
AN2X1 gate10666(.O (g32014), .I1 (g8715), .I2 (g30673));
AN2X1 gate10667(.O (g29969), .I1 (g28121), .I2 (g20509));
AN2X1 gate10668(.O (g30075), .I1 (g28525), .I2 (g20662));
AN2X1 gate10669(.O (g26155), .I1 (g1945), .I2 (g25134));
AN2X1 gate10670(.O (g14221), .I1 (g8686), .I2 (g11823));
AN2X1 gate10671(.O (g21921), .I1 (g5109), .I2 (g21468));
AN2X1 gate10672(.O (g26822), .I1 (g24841), .I2 (g13116));
AN4X1 gate10673(.O (I31242), .I1 (g32805), .I2 (g32806), .I3 (g32807), .I4 (g32808));
AN4X1 gate10674(.O (g16486), .I1 (g6772), .I2 (g11592), .I3 (g6789), .I4 (I17692));
AN2X1 gate10675(.O (g18592), .I1 (g2994), .I2 (g16349));
AN2X1 gate10676(.O (g23921), .I1 (g19379), .I2 (g4146));
AN2X1 gate10677(.O (g18756), .I1 (g5348), .I2 (g15595));
AN2X1 gate10678(.O (g34075), .I1 (g33692), .I2 (g19517));
AN2X1 gate10679(.O (g31526), .I1 (g22521), .I2 (g29342));
AN2X1 gate10680(.O (g24634), .I1 (g22634), .I2 (g19685));
AN2X1 gate10681(.O (g30595), .I1 (g18911), .I2 (g29847));
AN3X1 gate10682(.O (g33526), .I1 (g32932), .I2 (I31326), .I3 (I31327));
AN2X1 gate10683(.O (g24872), .I1 (g23088), .I2 (g9104));
AN2X1 gate10684(.O (g29968), .I1 (g2433), .I2 (g28843));
AN2X1 gate10685(.O (g21745), .I1 (g3017), .I2 (g20330));
AN2X1 gate10686(.O (g18780), .I1 (g5827), .I2 (g18065));
AN2X1 gate10687(.O (g12027), .I1 (g9499), .I2 (g9729));
AN2X1 gate10688(.O (g14613), .I1 (g10602), .I2 (g10585));
AN2X1 gate10689(.O (g27249), .I1 (g25929), .I2 (g19678));
AN2X1 gate10690(.O (g21799), .I1 (g3530), .I2 (g20924));
AN2X1 gate10691(.O (g29855), .I1 (g2287), .I2 (g29093));
AN2X1 gate10692(.O (g17770), .I1 (g7863), .I2 (g13189));
AN2X1 gate10693(.O (g21813), .I1 (g3590), .I2 (g20924));
AN2X1 gate10694(.O (g23799), .I1 (g14911), .I2 (g21279));
AN2X1 gate10695(.O (g27482), .I1 (g26488), .I2 (g17641));
AN2X1 gate10696(.O (g15815), .I1 (g3594), .I2 (g14075));
AN2X1 gate10697(.O (g28541), .I1 (g27403), .I2 (g20274));
AN2X1 gate10698(.O (g10947), .I1 (g9200), .I2 (g1430));
AN2X1 gate10699(.O (g18350), .I1 (g1779), .I2 (g17955));
AN3X1 gate10700(.O (I24603), .I1 (g9892), .I2 (g9467), .I3 (g6439));
AN2X1 gate10701(.O (g33402), .I1 (g32351), .I2 (g21395));
AN2X1 gate10702(.O (g29870), .I1 (g2421), .I2 (g29130));
AN2X1 gate10703(.O (g29527), .I1 (g28945), .I2 (g22432));
AN2X1 gate10704(.O (g27710), .I1 (g26422), .I2 (g20904));
AN2X1 gate10705(.O (g21798), .I1 (g3522), .I2 (g20924));
AN2X1 gate10706(.O (g34782), .I1 (g34711), .I2 (g33888));
AN4X1 gate10707(.O (I27529), .I1 (g28038), .I2 (g24121), .I3 (g24122), .I4 (g24123));
AN2X1 gate10708(.O (g18820), .I1 (g15166), .I2 (g15563));
AN2X1 gate10709(.O (g26853), .I1 (g94), .I2 (g24533));
AN4X1 gate10710(.O (g28789), .I1 (g21434), .I2 (g26424), .I3 (g25340), .I4 (g27440));
AN2X1 gate10711(.O (g21973), .I1 (g5511), .I2 (g19074));
AN2X1 gate10712(.O (g32116), .I1 (g31658), .I2 (g29929));
AN2X1 gate10713(.O (g27204), .I1 (g26026), .I2 (g16689));
AN2X1 gate10714(.O (g33866), .I1 (g33276), .I2 (g20528));
AN2X1 gate10715(.O (g22899), .I1 (g19486), .I2 (g19695));
AN2X1 gate10716(.O (g21805), .I1 (g3550), .I2 (g20924));
AN2X1 gate10717(.O (g22990), .I1 (g19555), .I2 (g19760));
AN4X1 gate10718(.O (I27528), .I1 (g20998), .I2 (g24118), .I3 (g24119), .I4 (g24120));
AN2X1 gate10719(.O (g18152), .I1 (g613), .I2 (g17533));
AN2X1 gate10720(.O (g25915), .I1 (g24926), .I2 (g9602));
AN2X1 gate10721(.O (g32041), .I1 (g13913), .I2 (g31262));
AN2X1 gate10722(.O (g18396), .I1 (g2008), .I2 (g15373));
AN2X1 gate10723(.O (g22633), .I1 (g19359), .I2 (g19479));
AN4X1 gate10724(.O (g17767), .I1 (g6772), .I2 (g11592), .I3 (g6789), .I4 (I18765));
AN2X1 gate10725(.O (g18731), .I1 (g15140), .I2 (g16861));
AN2X1 gate10726(.O (g30266), .I1 (g28775), .I2 (g23966));
AN2X1 gate10727(.O (g28535), .I1 (g11981), .I2 (g27088));
AN2X1 gate10728(.O (g15937), .I1 (g11950), .I2 (g14387));
AN2X1 gate10729(.O (g25201), .I1 (g12346), .I2 (g23665));
AN2X1 gate10730(.O (g22191), .I1 (g8119), .I2 (g19875));
AN2X1 gate10731(.O (g16179), .I1 (g6187), .I2 (g14321));
AN2X1 gate10732(.O (g29867), .I1 (g1996), .I2 (g29117));
AN2X1 gate10733(.O (g29894), .I1 (g2070), .I2 (g29169));
AN2X1 gate10734(.O (g19069), .I1 (g8397), .I2 (g16186));
AN2X1 gate10735(.O (g21732), .I1 (g3004), .I2 (g20330));
AN2X1 gate10736(.O (g16531), .I1 (g5232), .I2 (g14656));
AN2X1 gate10737(.O (g13542), .I1 (g10053), .I2 (g11927));
AN2X1 gate10738(.O (g21934), .I1 (g5220), .I2 (g18997));
AN2X1 gate10739(.O (g18413), .I1 (g2089), .I2 (g15373));
AN2X1 gate10740(.O (g24912), .I1 (g23687), .I2 (g20682));
AN2X1 gate10741(.O (g26119), .I1 (g11944), .I2 (g25109));
AN2X1 gate10742(.O (g24311), .I1 (g4498), .I2 (g22228));
AN2X1 gate10743(.O (g16178), .I1 (g5845), .I2 (g14297));
AN2X1 gate10744(.O (g18691), .I1 (g4727), .I2 (g16053));
AN2X1 gate10745(.O (g15884), .I1 (g3901), .I2 (g14113));
AN2X1 gate10746(.O (g33689), .I1 (g33144), .I2 (g11006));
AN2X1 gate10747(.O (g32340), .I1 (g31468), .I2 (g23585));
AN2X1 gate10748(.O (g29581), .I1 (g28462), .I2 (g11796));
AN2X1 gate10749(.O (g32035), .I1 (g4176), .I2 (g30937));
AN2X1 gate10750(.O (g31280), .I1 (g29717), .I2 (g23305));
AN2X1 gate10751(.O (g17191), .I1 (g1384), .I2 (g13242));
AN2X1 gate10752(.O (g17719), .I1 (g9818), .I2 (g14675));
AN2X1 gate10753(.O (g21761), .I1 (g3215), .I2 (g20785));
AN3X1 gate10754(.O (g29315), .I1 (g29188), .I2 (g7051), .I3 (g5990));
AN4X1 gate10755(.O (g27999), .I1 (g23032), .I2 (g26200), .I3 (g26424), .I4 (g25529));
AN2X1 gate10756(.O (g26864), .I1 (g2907), .I2 (g24548));
AN2X1 gate10757(.O (g26022), .I1 (g25271), .I2 (g20751));
AN2X1 gate10758(.O (g13436), .I1 (g9721), .I2 (g11811));
AN2X1 gate10759(.O (g18405), .I1 (g2040), .I2 (g15373));
AN2X1 gate10760(.O (g31300), .I1 (g30148), .I2 (g27858));
AN2X1 gate10761(.O (g30167), .I1 (g28622), .I2 (g23793));
AN2X1 gate10762(.O (g30194), .I1 (g28651), .I2 (g23849));
AN2X1 gate10763(.O (g30589), .I1 (g18898), .I2 (g29811));
AN4X1 gate10764(.O (I24690), .I1 (g24043), .I2 (g24044), .I3 (g24045), .I4 (g24046));
AN3X1 gate10765(.O (I24549), .I1 (g5385), .I2 (g5390), .I3 (g9792));
AN2X1 gate10766(.O (g26749), .I1 (g24494), .I2 (g23578));
AN2X1 gate10767(.O (g27090), .I1 (g25997), .I2 (g16423));
AN3X1 gate10768(.O (g29202), .I1 (g24088), .I2 (I27508), .I3 (I27509));
AN2X1 gate10769(.O (g25782), .I1 (g2936), .I2 (g24571));
AN2X1 gate10770(.O (g32142), .I1 (g31616), .I2 (g29965));
AN2X1 gate10771(.O (g13320), .I1 (g417), .I2 (g11048));
AN2X1 gate10772(.O (g26313), .I1 (g12645), .I2 (g25326));
AN3X1 gate10773(.O (g28291), .I1 (g7411), .I2 (g2070), .I3 (g27469));
AN2X1 gate10774(.O (g29979), .I1 (g23655), .I2 (g28991));
AN2X1 gate10775(.O (g34588), .I1 (g26082), .I2 (g34323));
AN2X1 gate10776(.O (g22861), .I1 (g19792), .I2 (g19670));
AN2X1 gate10777(.O (g27651), .I1 (g22448), .I2 (g25781));
AN2X1 gate10778(.O (g34524), .I1 (g9083), .I2 (g34359));
AN2X1 gate10779(.O (g33102), .I1 (g32399), .I2 (g18978));
AN4X1 gate10780(.O (I31007), .I1 (g32466), .I2 (g32467), .I3 (g32468), .I4 (g32469));
AN2X1 gate10781(.O (g26276), .I1 (g2461), .I2 (g25476));
AN2X1 gate10782(.O (g26285), .I1 (g1834), .I2 (g25300));
AN2X1 gate10783(.O (g34401), .I1 (g34199), .I2 (g21383));
AN2X1 gate10784(.O (g34477), .I1 (g26344), .I2 (g34328));
AN2X1 gate10785(.O (g22045), .I1 (g6069), .I2 (g21611));
AN2X1 gate10786(.O (g18583), .I1 (g2936), .I2 (g16349));
AN2X1 gate10787(.O (g29590), .I1 (g2625), .I2 (g28615));
AN3X1 gate10788(.O (g34119), .I1 (g20516), .I2 (g9104), .I3 (g33755));
AN2X1 gate10789(.O (g26254), .I1 (g2413), .I2 (g25349));
AN2X1 gate10790(.O (g31066), .I1 (g29483), .I2 (g22865));
AN2X1 gate10791(.O (g31231), .I1 (g30290), .I2 (g25239));
AN2X1 gate10792(.O (g29986), .I1 (g28468), .I2 (g23473));
AN2X1 gate10793(.O (g22099), .I1 (g6462), .I2 (g18833));
AN2X1 gate10794(.O (g27932), .I1 (g25944), .I2 (g19369));
AN2X1 gate10795(.O (g27331), .I1 (g10177), .I2 (g26754));
AN2X1 gate10796(.O (g30118), .I1 (g28574), .I2 (g21050));
AN2X1 gate10797(.O (g24820), .I1 (g13944), .I2 (g23978));
AN2X1 gate10798(.O (g26808), .I1 (g25521), .I2 (g21185));
AN2X1 gate10799(.O (g16762), .I1 (g5901), .I2 (g14930));
AN2X1 gate10800(.O (g20152), .I1 (g11545), .I2 (g16727));
AN2X1 gate10801(.O (g22534), .I1 (g8766), .I2 (g21389));
AN3X1 gate10802(.O (g29384), .I1 (g26424), .I2 (g22763), .I3 (g28179));
AN2X1 gate10803(.O (g22098), .I1 (g6459), .I2 (g18833));
AN2X1 gate10804(.O (g32193), .I1 (g30732), .I2 (g25410));
AN4X1 gate10805(.O (I31116), .I1 (g31154), .I2 (g31816), .I3 (g32622), .I4 (g32623));
AN3X1 gate10806(.O (g24846), .I1 (g3361), .I2 (g23555), .I3 (I24018));
AN2X1 gate10807(.O (g26101), .I1 (g1760), .I2 (g25098));
AN2X1 gate10808(.O (g33876), .I1 (g33286), .I2 (g20562));
AN2X1 gate10809(.O (g33885), .I1 (g33296), .I2 (g20609));
AN2X1 gate10810(.O (g26177), .I1 (g2079), .I2 (g25154));
AN2X1 gate10811(.O (g18113), .I1 (g405), .I2 (g17015));
AN2X1 gate10812(.O (g18787), .I1 (g15158), .I2 (g15634));
AN2X1 gate10813(.O (g32165), .I1 (g31669), .I2 (g27742));
AN2X1 gate10814(.O (g24731), .I1 (g6519), .I2 (g23733));
AN4X1 gate10815(.O (I31041), .I1 (g31566), .I2 (g31803), .I3 (g32513), .I4 (g32514));
AN2X1 gate10816(.O (g18282), .I1 (g1379), .I2 (g16136));
AN2X1 gate10817(.O (g34748), .I1 (g34672), .I2 (g19529));
AN2X1 gate10818(.O (g27505), .I1 (g26519), .I2 (g17681));
AN2X1 gate10819(.O (g27404), .I1 (g26400), .I2 (g17518));
AN2X1 gate10820(.O (g31763), .I1 (g30127), .I2 (g23965));
AN2X1 gate10821(.O (g18302), .I1 (g1514), .I2 (g16489));
AN3X1 gate10822(.O (g33511), .I1 (g32823), .I2 (I31251), .I3 (I31252));
AN2X1 gate10823(.O (g15084), .I1 (g2710), .I2 (g12983));
AN2X1 gate10824(.O (g18357), .I1 (g1816), .I2 (g17955));
AN2X1 gate10825(.O (g19545), .I1 (g3147), .I2 (g16769));
AN2X1 gate10826(.O (g29877), .I1 (g28405), .I2 (g23340));
AN2X1 gate10827(.O (g15110), .I1 (g4245), .I2 (g14454));
AN2X1 gate10828(.O (g18105), .I1 (g417), .I2 (g17015));
AN2X1 gate10829(.O (g10724), .I1 (g3689), .I2 (g8728));
AN2X1 gate10830(.O (g22032), .I1 (g5921), .I2 (g19147));
AN2X1 gate10831(.O (g30254), .I1 (g28747), .I2 (g23944));
AN2X1 gate10832(.O (g18743), .I1 (g5115), .I2 (g17847));
AN2X1 gate10833(.O (g27212), .I1 (g25997), .I2 (g16717));
AN2X1 gate10834(.O (g10829), .I1 (g7289), .I2 (g4375));
AN4X1 gate10835(.O (I31237), .I1 (g32798), .I2 (g32799), .I3 (g32800), .I4 (g32801));
AN2X1 gate10836(.O (g21771), .I1 (g3255), .I2 (g20785));
AN2X1 gate10837(.O (g10828), .I1 (g6888), .I2 (g7640));
AN2X1 gate10838(.O (g18640), .I1 (g3835), .I2 (g17096));
AN2X1 gate10839(.O (g18769), .I1 (g15151), .I2 (g18062));
AN2X1 gate10840(.O (g22061), .I1 (g6065), .I2 (g21611));
AN2X1 gate10841(.O (g30101), .I1 (g28551), .I2 (g20780));
AN2X1 gate10842(.O (g30177), .I1 (g28631), .I2 (g23814));
AN2X1 gate10843(.O (g29526), .I1 (g28938), .I2 (g22384));
AN2X1 gate10844(.O (g17140), .I1 (g8616), .I2 (g12968));
AN2X1 gate10845(.O (g26630), .I1 (g7592), .I2 (g24419));
AN2X1 gate10846(.O (g34560), .I1 (g34366), .I2 (g17366));
AN2X1 gate10847(.O (g18768), .I1 (g5503), .I2 (g17929));
AN2X1 gate10848(.O (g18803), .I1 (g15161), .I2 (g15480));
AN2X1 gate10849(.O (g31480), .I1 (g1644), .I2 (g30296));
AN4X1 gate10850(.O (I31142), .I1 (g32661), .I2 (g32662), .I3 (g32663), .I4 (g32664));
AN3X1 gate10851(.O (g33480), .I1 (g32600), .I2 (I31096), .I3 (I31097));
AN2X1 gate10852(.O (g24929), .I1 (g23751), .I2 (g20875));
AN2X1 gate10853(.O (g22871), .I1 (g9523), .I2 (g20871));
AN4X1 gate10854(.O (g26166), .I1 (g25357), .I2 (g11724), .I3 (g11709), .I4 (g7558));
AN2X1 gate10855(.O (g27723), .I1 (g26512), .I2 (g21049));
AN2X1 gate10856(.O (g15654), .I1 (g3845), .I2 (g13584));
AN2X1 gate10857(.O (g31314), .I1 (g30183), .I2 (g27937));
AN2X1 gate10858(.O (g28240), .I1 (g27356), .I2 (g17239));
AN2X1 gate10859(.O (g27149), .I1 (g25997), .I2 (g16623));
AN2X1 gate10860(.O (g30064), .I1 (g28517), .I2 (g20630));
AN4X1 gate10861(.O (g17766), .I1 (g6772), .I2 (g11592), .I3 (g11640), .I4 (I18762));
AN2X1 gate10862(.O (g27433), .I1 (g26519), .I2 (g17583));
AN2X1 gate10863(.O (g27387), .I1 (g26488), .I2 (g17499));
AN2X1 gate10864(.O (g15936), .I1 (g475), .I2 (g13999));
AN2X1 gate10865(.O (g25285), .I1 (g22152), .I2 (g13061));
AN2X1 gate10866(.O (g29866), .I1 (g1906), .I2 (g29116));
AN2X1 gate10867(.O (g27148), .I1 (g25997), .I2 (g16622));
AN2X1 gate10868(.O (g21882), .I1 (g4057), .I2 (g19801));
AN2X1 gate10869(.O (g21991), .I1 (g5595), .I2 (g19074));
AN2X1 gate10870(.O (g26485), .I1 (g24968), .I2 (g10502));
AN2X1 gate10871(.O (g23991), .I1 (g19209), .I2 (g21428));
AN2X1 gate10872(.O (g27097), .I1 (g25867), .I2 (g22526));
AN2X1 gate10873(.O (g33721), .I1 (g33163), .I2 (g19440));
AN2X1 gate10874(.O (g19656), .I1 (g2807), .I2 (g15844));
AN2X1 gate10875(.O (g27104), .I1 (g25997), .I2 (g16510));
AN2X1 gate10876(.O (g16751), .I1 (g13155), .I2 (g13065));
AN2X1 gate10877(.O (g16807), .I1 (g6585), .I2 (g14978));
AN2X1 gate10878(.O (g27646), .I1 (g13094), .I2 (g25773));
AN2X1 gate10879(.O (g25900), .I1 (g24390), .I2 (g19368));
AN2X1 gate10880(.O (g34874), .I1 (g34833), .I2 (g20060));
AN2X1 gate10881(.O (g23407), .I1 (g9295), .I2 (g20273));
AN2X1 gate10882(.O (g33243), .I1 (g32124), .I2 (g19947));
AN2X1 gate10883(.O (g28563), .I1 (g11981), .I2 (g27100));
AN2X1 gate10884(.O (g25466), .I1 (g23574), .I2 (g21346));
AN2X1 gate10885(.O (g19680), .I1 (g12028), .I2 (g17013));
AN2X1 gate10886(.O (g33431), .I1 (g32364), .I2 (g32377));
AN2X1 gate10887(.O (g16639), .I1 (g6291), .I2 (g14974));
AN2X1 gate10888(.O (g26712), .I1 (g24508), .I2 (g24463));
AN3X1 gate10889(.O (I17741), .I1 (g14988), .I2 (g11450), .I3 (g11498));
AN2X1 gate10890(.O (g18662), .I1 (g15126), .I2 (g17367));
AN2X1 gate10891(.O (g32175), .I1 (g31709), .I2 (g27858));
AN2X1 gate10892(.O (g30166), .I1 (g28621), .I2 (g23792));
AN2X1 gate10893(.O (g30009), .I1 (g29034), .I2 (g10518));
AN2X1 gate10894(.O (g24302), .I1 (g15124), .I2 (g22228));
AN2X1 gate10895(.O (g16638), .I1 (g6271), .I2 (g14773));
AN2X1 gate10896(.O (g33269), .I1 (g31970), .I2 (g15582));
AN2X1 gate10897(.O (g34665), .I1 (g34583), .I2 (g19067));
AN3X1 gate10898(.O (g22472), .I1 (g7753), .I2 (g9285), .I3 (g21289));
AN2X1 gate10899(.O (g18890), .I1 (g10158), .I2 (g17625));
AN2X1 gate10900(.O (g13492), .I1 (g9856), .I2 (g11865));
AN2X1 gate10901(.O (g27369), .I1 (g25894), .I2 (g25324));
AN2X1 gate10902(.O (g24743), .I1 (g22708), .I2 (g19789));
AN2X1 gate10903(.O (g30008), .I1 (g29191), .I2 (g12297));
AN2X1 gate10904(.O (g18249), .I1 (g1216), .I2 (g16897));
AN2X1 gate10905(.O (g33942), .I1 (g33383), .I2 (g21608));
AN2X1 gate10906(.O (g33341), .I1 (g32223), .I2 (g20640));
AN2X1 gate10907(.O (g18482), .I1 (g2472), .I2 (g15426));
AN2X1 gate10908(.O (g14506), .I1 (g1430), .I2 (g10755));
AN2X1 gate10909(.O (g29688), .I1 (g2509), .I2 (g28713));
AN4X1 gate10910(.O (I31006), .I1 (g31376), .I2 (g31796), .I3 (g32464), .I4 (g32465));
AN2X1 gate10911(.O (g29624), .I1 (g28491), .I2 (g8070));
AN2X1 gate10912(.O (g14028), .I1 (g8673), .I2 (g11797));
AN2X1 gate10913(.O (g18248), .I1 (g15067), .I2 (g16897));
AN2X1 gate10914(.O (g16841), .I1 (g5913), .I2 (g14858));
AN2X1 gate10915(.O (g18710), .I1 (g15135), .I2 (g17302));
AN2X1 gate10916(.O (g34476), .I1 (g34399), .I2 (g18891));
AN2X1 gate10917(.O (g34485), .I1 (g34411), .I2 (g18952));
AN2X1 gate10918(.O (g18552), .I1 (g2815), .I2 (g15277));
AN2X1 gate10919(.O (g24640), .I1 (g6509), .I2 (g23733));
AN2X1 gate10920(.O (g24769), .I1 (g19619), .I2 (g23058));
AN2X1 gate10921(.O (g19631), .I1 (g1484), .I2 (g16093));
AN2X1 gate10922(.O (g18204), .I1 (g914), .I2 (g15938));
AN4X1 gate10923(.O (I31222), .I1 (g32775), .I2 (g32776), .I3 (g32777), .I4 (g32778));
AN2X1 gate10924(.O (g27412), .I1 (g26576), .I2 (g17529));
AN2X1 gate10925(.O (g34555), .I1 (g34349), .I2 (g20512));
AN2X1 gate10926(.O (g18779), .I1 (g5821), .I2 (g18065));
AN2X1 gate10927(.O (g22071), .I1 (g6251), .I2 (g19210));
AN2X1 gate10928(.O (g24803), .I1 (g22901), .I2 (g20005));
AN3X1 gate10929(.O (g33734), .I1 (g7806), .I2 (g33136), .I3 (I31593));
AN2X1 gate10930(.O (g30914), .I1 (g29873), .I2 (g20887));
AN2X1 gate10931(.O (g21759), .I1 (g3199), .I2 (g20785));
AN2X1 gate10932(.O (g15117), .I1 (g4300), .I2 (g14454));
AN2X1 gate10933(.O (g23725), .I1 (g14772), .I2 (g21138));
AN2X1 gate10934(.O (g18778), .I1 (g5817), .I2 (g18065));
AN2X1 gate10935(.O (g25874), .I1 (g11118), .I2 (g24665));
AN2X1 gate10936(.O (g27229), .I1 (g26055), .I2 (g16774));
AN2X1 gate10937(.O (g31993), .I1 (g31774), .I2 (g22214));
AN2X1 gate10938(.O (g21758), .I1 (g3191), .I2 (g20785));
AN2X1 gate10939(.O (g26176), .I1 (g1964), .I2 (g25467));
AN2X1 gate10940(.O (g26092), .I1 (g9766), .I2 (g25083));
AN2X1 gate10941(.O (g18786), .I1 (g15156), .I2 (g15345));
AN2X1 gate10942(.O (g27228), .I1 (g26055), .I2 (g16773));
AN3X1 gate10943(.O (g24881), .I1 (g3050), .I2 (g23211), .I3 (I24048));
AN4X1 gate10944(.O (I31347), .I1 (g32956), .I2 (g32957), .I3 (g32958), .I4 (g32959));
AN2X1 gate10945(.O (g22859), .I1 (g9456), .I2 (g20734));
AN2X1 gate10946(.O (g26154), .I1 (g1830), .I2 (g25426));
AN2X1 gate10947(.O (g30239), .I1 (g28728), .I2 (g23923));
AN2X1 gate10948(.O (g17785), .I1 (g13341), .I2 (g10762));
AN2X1 gate10949(.O (g25166), .I1 (g17506), .I2 (g23571));
AN2X1 gate10950(.O (g31131), .I1 (g2393), .I2 (g30020));
AN2X1 gate10951(.O (g18647), .I1 (g4040), .I2 (g17271));
AN2X1 gate10952(.O (g34074), .I1 (g33685), .I2 (g19498));
AN2X1 gate10953(.O (g30594), .I1 (g18898), .I2 (g29846));
AN2X1 gate10954(.O (g18356), .I1 (g1802), .I2 (g17955));
AN2X1 gate10955(.O (g29876), .I1 (g28404), .I2 (g23339));
AN2X1 gate10956(.O (g29885), .I1 (g28416), .I2 (g23350));
AN2X1 gate10957(.O (g21744), .I1 (g3103), .I2 (g20330));
AN2X1 gate10958(.O (g30238), .I1 (g28727), .I2 (g23922));
AN2X1 gate10959(.O (g34567), .I1 (g34377), .I2 (g17491));
AN3X1 gate10960(.O (I31600), .I1 (g31009), .I2 (g8400), .I3 (g7809));
AN2X1 gate10961(.O (g28440), .I1 (g27274), .I2 (g20059));
AN2X1 gate10962(.O (g18826), .I1 (g7097), .I2 (g15680));
AN2X1 gate10963(.O (g18380), .I1 (g1926), .I2 (g15171));
AN2X1 gate10964(.O (g19571), .I1 (g3498), .I2 (g16812));
AN3X1 gate10965(.O (g33487), .I1 (g32649), .I2 (I31131), .I3 (I31132));
AN2X1 gate10966(.O (g22172), .I1 (g8064), .I2 (g19857));
AN2X1 gate10967(.O (g29854), .I1 (g2197), .I2 (g29092));
AN2X1 gate10968(.O (g21849), .I1 (g3889), .I2 (g21070));
AN2X1 gate10969(.O (g21940), .I1 (g5228), .I2 (g18997));
AN4X1 gate10970(.O (I31236), .I1 (g30735), .I2 (g31837), .I3 (g32796), .I4 (g32797));
AN2X1 gate10971(.O (g15814), .I1 (g3574), .I2 (g13920));
AN2X1 gate10972(.O (g31502), .I1 (g2472), .I2 (g29311));
AN2X1 gate10973(.O (g28573), .I1 (g7349), .I2 (g27059));
AN3X1 gate10974(.O (g25485), .I1 (g6098), .I2 (g22220), .I3 (I24600));
AN3X1 gate10975(.O (g33502), .I1 (g32758), .I2 (I31206), .I3 (I31207));
AN2X1 gate10976(.O (g29511), .I1 (g1736), .I2 (g28783));
AN2X1 gate10977(.O (g31210), .I1 (g2509), .I2 (g30100));
AN4X1 gate10978(.O (I31351), .I1 (g30937), .I2 (g31858), .I3 (g32961), .I4 (g32962));
AN2X1 gate10979(.O (g18233), .I1 (g1094), .I2 (g16326));
AN2X1 gate10980(.O (g28247), .I1 (g27147), .I2 (g19675));
AN2X1 gate10981(.O (g21848), .I1 (g3913), .I2 (g21070));
AN2X1 gate10982(.O (g15807), .I1 (g3570), .I2 (g13898));
AN2X1 gate10983(.O (g18182), .I1 (g776), .I2 (g17328));
AN2X1 gate10984(.O (g27310), .I1 (g26574), .I2 (g23059));
AN2X1 gate10985(.O (g18651), .I1 (g15102), .I2 (g16249));
AN2X1 gate10986(.O (g18672), .I1 (g15127), .I2 (g15758));
AN2X1 gate10987(.O (g34382), .I1 (g34167), .I2 (g20618));
AN2X1 gate10988(.O (g30185), .I1 (g28640), .I2 (g23838));
AN2X1 gate10989(.O (g34519), .I1 (g34293), .I2 (g19504));
AN2X1 gate10990(.O (g17151), .I1 (g8659), .I2 (g12996));
AN2X1 gate10991(.O (g21804), .I1 (g3542), .I2 (g20924));
AN2X1 gate10992(.O (g34185), .I1 (g33702), .I2 (g24389));
AN2X1 gate10993(.O (g27627), .I1 (g13266), .I2 (g25790));
AN2X1 gate10994(.O (g25570), .I1 (I24689), .I2 (I24690));
AN2X1 gate10995(.O (g27959), .I1 (g25948), .I2 (g19374));
AN2X1 gate10996(.O (g28612), .I1 (g27524), .I2 (g20539));
AN3X1 gate10997(.O (g34092), .I1 (g33750), .I2 (g9104), .I3 (g18957));
AN2X1 gate10998(.O (g30154), .I1 (g28611), .I2 (g23769));
AN2X1 gate10999(.O (g28324), .I1 (g9875), .I2 (g27687));
AN2X1 gate11000(.O (g24482), .I1 (g6875), .I2 (g23055));
AN2X1 gate11001(.O (g31278), .I1 (g29716), .I2 (g23302));
AN2X1 gate11002(.O (g34518), .I1 (g34292), .I2 (g19503));
AN2X1 gate11003(.O (g32274), .I1 (g31256), .I2 (g20447));
AN2X1 gate11004(.O (g27050), .I1 (g25789), .I2 (g22338));
AN2X1 gate11005(.O (g27958), .I1 (g25950), .I2 (g22449));
AN2X1 gate11006(.O (g25907), .I1 (g24799), .I2 (g22519));
AN2X1 gate11007(.O (g24710), .I1 (g22679), .I2 (g19771));
AN2X1 gate11008(.O (g27378), .I1 (g26089), .I2 (g20052));
AN4X1 gate11009(.O (I31137), .I1 (g32654), .I2 (g32655), .I3 (g32656), .I4 (g32657));
AN2X1 gate11010(.O (g18331), .I1 (g1682), .I2 (g17873));
AN3X1 gate11011(.O (I27364), .I1 (g25541), .I2 (g26424), .I3 (g22698));
AN2X1 gate11012(.O (g24552), .I1 (g22487), .I2 (g19538));
AN3X1 gate11013(.O (g33469), .I1 (g32519), .I2 (I31041), .I3 (I31042));
AN2X1 gate11014(.O (g28251), .I1 (g27826), .I2 (g23662));
AN2X1 gate11015(.O (g30935), .I1 (g8808), .I2 (g29745));
AN2X1 gate11016(.O (g28272), .I1 (g27721), .I2 (g26548));
AN2X1 gate11017(.O (g31286), .I1 (g30159), .I2 (g27858));
AN2X1 gate11018(.O (g32122), .I1 (g31646), .I2 (g29944));
AN2X1 gate11019(.O (g18513), .I1 (g2575), .I2 (g15509));
AN2X1 gate11020(.O (g21332), .I1 (g996), .I2 (g15739));
AN2X1 gate11021(.O (g18449), .I1 (g12852), .I2 (g15224));
AN3X1 gate11022(.O (I26972), .I1 (g25011), .I2 (g26424), .I3 (g22698));
AN2X1 gate11023(.O (g27386), .I1 (g26488), .I2 (g17498));
AN2X1 gate11024(.O (g19752), .I1 (g2771), .I2 (g15864));
AN3X1 gate11025(.O (g33468), .I1 (g32512), .I2 (I31036), .I3 (I31037));
AN2X1 gate11026(.O (g15841), .I1 (g4273), .I2 (g13868));
AN2X1 gate11027(.O (g25567), .I1 (I24674), .I2 (I24675));
AN2X1 gate11028(.O (g27096), .I1 (g26026), .I2 (g16475));
AN2X1 gate11029(.O (g18448), .I1 (g2153), .I2 (g18008));
AN2X1 gate11030(.O (g29550), .I1 (g28990), .I2 (g22457));
AN2X1 gate11031(.O (g32034), .I1 (g14124), .I2 (g31239));
AN2X1 gate11032(.O (g25238), .I1 (g12466), .I2 (g23732));
AN2X1 gate11033(.O (g16806), .I1 (g6247), .I2 (g14971));
AN2X1 gate11034(.O (g29314), .I1 (g29005), .I2 (g22144));
AN2X1 gate11035(.O (g22059), .I1 (g6148), .I2 (g21611));
AN2X1 gate11036(.O (g21962), .I1 (g5428), .I2 (g21514));
AN2X1 gate11037(.O (g18505), .I1 (g2583), .I2 (g15509));
AN2X1 gate11038(.O (g21361), .I1 (g7869), .I2 (g16066));
AN2X1 gate11039(.O (g22025), .I1 (g5905), .I2 (g19147));
AN2X1 gate11040(.O (g18404), .I1 (g2066), .I2 (g15373));
AN2X1 gate11041(.O (g24786), .I1 (g661), .I2 (g23654));
AN2X1 gate11042(.O (g33815), .I1 (g33449), .I2 (g12911));
AN2X1 gate11043(.O (g32292), .I1 (g31269), .I2 (g20530));
AN2X1 gate11044(.O (g10898), .I1 (g3706), .I2 (g9100));
AN2X1 gate11045(.O (g18717), .I1 (g4849), .I2 (g15915));
AN2X1 gate11046(.O (g22058), .I1 (g6098), .I2 (g21611));
AN2X1 gate11047(.O (g31187), .I1 (g10118), .I2 (g30090));
AN2X1 gate11048(.O (g32153), .I1 (g31646), .I2 (g29999));
AN2X1 gate11049(.O (g24647), .I1 (g19903), .I2 (g22907));
AN2X1 gate11050(.O (g33677), .I1 (g33443), .I2 (g31937));
AN2X1 gate11051(.O (g31975), .I1 (g31761), .I2 (g22177));
AN4X1 gate11052(.O (g13252), .I1 (g11561), .I2 (g11511), .I3 (g11469), .I4 (g699));
AN2X1 gate11053(.O (g18212), .I1 (g947), .I2 (g15979));
AN2X1 gate11054(.O (g29596), .I1 (g27823), .I2 (g28620));
AN2X1 gate11055(.O (g24945), .I1 (g23183), .I2 (g20197));
AN3X1 gate11056(.O (g10719), .I1 (g6841), .I2 (g2138), .I3 (g2130));
AN2X1 gate11057(.O (g16517), .I1 (g5248), .I2 (g14797));
AN2X1 gate11058(.O (g21833), .I1 (g15096), .I2 (g20453));
AN2X1 gate11059(.O (g30215), .I1 (g28690), .I2 (g23881));
AN2X1 gate11060(.O (g32409), .I1 (g4754), .I2 (g30996));
AN2X1 gate11061(.O (g14719), .I1 (g4392), .I2 (g10830));
AN2X1 gate11062(.O (g34215), .I1 (g33778), .I2 (g22670));
AN2X1 gate11063(.O (g30577), .I1 (g26267), .I2 (g29679));
AN2X1 gate11064(.O (g34577), .I1 (g24577), .I2 (g34307));
AN3X1 gate11065(.O (g25518), .I1 (g6444), .I2 (g23865), .I3 (I24625));
AN2X1 gate11066(.O (g27428), .I1 (g26400), .I2 (g17576));
AN2X1 gate11067(.O (g13564), .I1 (g4480), .I2 (g12820));
AN2X1 gate11068(.O (g22044), .I1 (g6058), .I2 (g21611));
AN2X1 gate11069(.O (g26304), .I1 (g2697), .I2 (g25246));
AN2X1 gate11070(.O (g31143), .I1 (g29506), .I2 (g22999));
AN4X1 gate11071(.O (I24709), .I1 (g21256), .I2 (g24068), .I3 (g24069), .I4 (g24070));
AN4X1 gate11072(.O (I31021), .I1 (g31070), .I2 (g31799), .I3 (g32485), .I4 (g32486));
AN2X1 gate11073(.O (g24998), .I1 (g17412), .I2 (g23408));
AN2X1 gate11074(.O (g12730), .I1 (g9024), .I2 (g4349));
AN2X1 gate11075(.O (g27765), .I1 (g4146), .I2 (g25886));
AN2X1 gate11076(.O (g24651), .I1 (g2741), .I2 (g23472));
AN2X1 gate11077(.O (g24672), .I1 (g19534), .I2 (g22981));
AN2X1 gate11078(.O (g14832), .I1 (g1489), .I2 (g10939));
AN2X1 gate11079(.O (g29773), .I1 (g28203), .I2 (g10233));
AN2X1 gate11080(.O (g27690), .I1 (g25784), .I2 (g23607));
AN2X1 gate11081(.O (g16193), .I1 (g6533), .I2 (g14348));
AN2X1 gate11082(.O (g27549), .I1 (g26576), .I2 (g14785));
AN2X1 gate11083(.O (g31169), .I1 (g10083), .I2 (g30079));
AN2X1 gate11084(.O (g11397), .I1 (g5360), .I2 (g7139));
AN2X1 gate11085(.O (g18723), .I1 (g4922), .I2 (g16077));
AN2X1 gate11086(.O (g25883), .I1 (g13728), .I2 (g24699));
AN2X1 gate11087(.O (g28360), .I1 (g27401), .I2 (g19861));
AN2X1 gate11088(.O (g22120), .I1 (g6585), .I2 (g19277));
AN2X1 gate11089(.O (g33884), .I1 (g33295), .I2 (g20590));
AN2X1 gate11090(.O (g15116), .I1 (g4297), .I2 (g14454));
AN2X1 gate11091(.O (g18149), .I1 (g608), .I2 (g17533));
AN2X1 gate11092(.O (g27548), .I1 (g26576), .I2 (g17763));
AN2X1 gate11093(.O (g31168), .I1 (g2241), .I2 (g30077));
AN2X1 gate11094(.O (g32164), .I1 (g30733), .I2 (g25171));
AN2X1 gate11095(.O (g18433), .I1 (g2197), .I2 (g18008));
AN2X1 gate11096(.O (g33410), .I1 (g32360), .I2 (g21409));
AN2X1 gate11097(.O (g18387), .I1 (g1955), .I2 (g15171));
AN2X1 gate11098(.O (g24331), .I1 (g6977), .I2 (g22228));
AN2X1 gate11099(.O (g30083), .I1 (g28533), .I2 (g20698));
AN2X1 gate11100(.O (g13509), .I1 (g9951), .I2 (g11889));
AN2X1 gate11101(.O (g27504), .I1 (g26519), .I2 (g17680));
AN2X1 gate11102(.O (g18620), .I1 (g3470), .I2 (g17062));
AN2X1 gate11103(.O (g18148), .I1 (g562), .I2 (g17533));
AN2X1 gate11104(.O (g21947), .I1 (g5256), .I2 (g18997));
AN2X1 gate11105(.O (g30284), .I1 (g28852), .I2 (g23994));
AN2X1 gate11106(.O (g34083), .I1 (g33714), .I2 (g19573));
AN2X1 gate11107(.O (g34348), .I1 (g34125), .I2 (g20128));
AN3X1 gate11108(.O (I31593), .I1 (g31003), .I2 (g8350), .I3 (g7788));
AN3X1 gate11109(.O (g33479), .I1 (g32593), .I2 (I31091), .I3 (I31092));
AN2X1 gate11110(.O (g34284), .I1 (g34046), .I2 (g19351));
AN2X1 gate11111(.O (g21605), .I1 (g13005), .I2 (g15695));
AN4X1 gate11112(.O (I31346), .I1 (g31021), .I2 (g31857), .I3 (g32954), .I4 (g32955));
AN2X1 gate11113(.O (g33363), .I1 (g32262), .I2 (g20918));
AN2X1 gate11114(.O (g13508), .I1 (g9927), .I2 (g11888));
AN2X1 gate11115(.O (g18104), .I1 (g392), .I2 (g17015));
AN2X1 gate11116(.O (g18811), .I1 (g6500), .I2 (g15483));
AN2X1 gate11117(.O (g18646), .I1 (g4031), .I2 (g17271));
AN4X1 gate11118(.O (I31122), .I1 (g32631), .I2 (g32632), .I3 (g32633), .I4 (g32634));
AN2X1 gate11119(.O (g14612), .I1 (g11971), .I2 (g11993));
AN2X1 gate11120(.O (g31478), .I1 (g29764), .I2 (g23410));
AN2X1 gate11121(.O (g8234), .I1 (g4515), .I2 (g4521));
AN2X1 gate11122(.O (g31015), .I1 (g29476), .I2 (g22758));
AN2X1 gate11123(.O (g18343), .I1 (g12847), .I2 (g17955));
AN3X1 gate11124(.O (g24897), .I1 (g3401), .I2 (g23223), .I3 (I24064));
AN2X1 gate11125(.O (g29839), .I1 (g1728), .I2 (g29045));
AN2X1 gate11126(.O (g30566), .I1 (g26247), .I2 (g29507));
AN3X1 gate11127(.O (g33478), .I1 (g32584), .I2 (I31086), .I3 (I31087));
AN2X1 gate11128(.O (g24961), .I1 (g23193), .I2 (g20209));
AN2X1 gate11129(.O (g21812), .I1 (g3586), .I2 (g20924));
AN2X1 gate11130(.O (g17146), .I1 (g5965), .I2 (g14895));
AN2X1 gate11131(.O (g34566), .I1 (g34376), .I2 (g17489));
AN2X1 gate11132(.O (g28451), .I1 (g27283), .I2 (g20090));
AN2X1 gate11133(.O (g16222), .I1 (g6513), .I2 (g14348));
AN2X1 gate11134(.O (g31486), .I1 (g29777), .I2 (g23422));
AN2X1 gate11135(.O (g32327), .I1 (g31319), .I2 (g23544));
AN2X1 gate11136(.O (g29667), .I1 (g2671), .I2 (g29157));
AN2X1 gate11137(.O (g29838), .I1 (g1636), .I2 (g29044));
AN2X1 gate11138(.O (g27129), .I1 (g26026), .I2 (g16584));
AN3X1 gate11139(.O (g33486), .I1 (g32642), .I2 (I31126), .I3 (I31127));
AN2X1 gate11140(.O (g32109), .I1 (g31609), .I2 (g29920));
AN2X1 gate11141(.O (g21951), .I1 (g5272), .I2 (g18997));
AN2X1 gate11142(.O (g26852), .I1 (g24975), .I2 (g24958));
AN2X1 gate11143(.O (g21972), .I1 (g15152), .I2 (g19074));
AN4X1 gate11144(.O (g27057), .I1 (g7791), .I2 (g6219), .I3 (g6227), .I4 (g26261));
AN2X1 gate11145(.O (g19610), .I1 (g1141), .I2 (g16069));
AN2X1 gate11146(.O (g18369), .I1 (g12848), .I2 (g15171));
AN2X1 gate11147(.O (g24717), .I1 (g22684), .I2 (g19777));
AN2X1 gate11148(.O (g27128), .I1 (g25997), .I2 (g16583));
AN2X1 gate11149(.O (g28246), .I1 (g8572), .I2 (g27976));
AN4X1 gate11150(.O (I31292), .I1 (g32877), .I2 (g32878), .I3 (g32879), .I4 (g32880));
AN2X1 gate11151(.O (g32108), .I1 (g31631), .I2 (g29913));
AN2X1 gate11152(.O (g30139), .I1 (g28596), .I2 (g21184));
AN2X1 gate11153(.O (g18368), .I1 (g1728), .I2 (g17955));
AN2X1 gate11154(.O (g34139), .I1 (g33827), .I2 (g23314));
AN2X1 gate11155(.O (g16703), .I1 (g5889), .I2 (g15002));
AN2X1 gate11156(.O (g22632), .I1 (g19356), .I2 (g19476));
AN2X1 gate11157(.O (g31223), .I1 (g20028), .I2 (g29689));
AN2X1 gate11158(.O (g21795), .I1 (g3506), .I2 (g20924));
AN2X1 gate11159(.O (g32283), .I1 (g31259), .I2 (g20506));
AN2X1 gate11160(.O (g27323), .I1 (g26268), .I2 (g23086));
AN2X1 gate11161(.O (g30138), .I1 (g28595), .I2 (g21182));
AN2X1 gate11162(.O (g27299), .I1 (g26546), .I2 (g23028));
AN2X1 gate11163(.O (g29619), .I1 (g2269), .I2 (g29060));
AN2X1 gate11164(.O (g32303), .I1 (g27550), .I2 (g31376));
AN2X1 gate11165(.O (g34138), .I1 (g33929), .I2 (g23828));
AN2X1 gate11166(.O (g11047), .I1 (g6474), .I2 (g9212));
AN2X1 gate11167(.O (g18412), .I1 (g2098), .I2 (g15373));
AN4X1 gate11168(.O (I31136), .I1 (g29385), .I2 (g32651), .I3 (g32652), .I4 (g32653));
AN2X1 gate11169(.O (g11205), .I1 (g8217), .I2 (g8439));
AN2X1 gate11170(.O (g13047), .I1 (g8534), .I2 (g11042));
AN2X1 gate11171(.O (g27298), .I1 (g26573), .I2 (g23026));
AN2X1 gate11172(.O (g29618), .I1 (g28870), .I2 (g22384));
AN2X1 gate11173(.O (g19383), .I1 (g16893), .I2 (g13223));
AN2X1 gate11174(.O (g34415), .I1 (g34207), .I2 (g21458));
AN2X1 gate11175(.O (g18133), .I1 (g15055), .I2 (g17249));
AN2X1 gate11176(.O (g23514), .I1 (g20149), .I2 (g11829));
AN2X1 gate11177(.O (g26484), .I1 (g24946), .I2 (g8841));
AN2X1 gate11178(.O (g33110), .I1 (g32404), .I2 (g32415));
AN2X1 gate11179(.O (g13912), .I1 (g5551), .I2 (g12450));
AN2X1 gate11180(.O (g34333), .I1 (g9984), .I2 (g34192));
AN2X1 gate11181(.O (g24723), .I1 (g17490), .I2 (g22384));
AN2X1 gate11182(.O (g31321), .I1 (g30146), .I2 (g27886));
AN2X1 gate11183(.O (g18229), .I1 (g1099), .I2 (g16326));
AN2X1 gate11184(.O (g33922), .I1 (g33448), .I2 (g7202));
AN2X1 gate11185(.O (g14061), .I1 (g8715), .I2 (g11834));
AN3X1 gate11186(.O (g33531), .I1 (g32967), .I2 (I31351), .I3 (I31352));
AN2X1 gate11187(.O (g18228), .I1 (g1061), .I2 (g16129));
AN2X1 gate11188(.O (g24387), .I1 (g3457), .I2 (g22761));
AN2X1 gate11189(.O (g26312), .I1 (g2704), .I2 (g25264));
AN2X1 gate11190(.O (g34963), .I1 (g34946), .I2 (g23041));
AN4X1 gate11191(.O (g26200), .I1 (g24688), .I2 (g10678), .I3 (g10658), .I4 (g10627));
AN2X1 gate11192(.O (g32174), .I1 (g31708), .I2 (g27837));
AN2X1 gate11193(.O (g21163), .I1 (g16321), .I2 (g4878));
AN2X1 gate11194(.O (g21012), .I1 (g16304), .I2 (g4688));
AN2X1 gate11195(.O (g28151), .I1 (g8426), .I2 (g27295));
AN2X1 gate11196(.O (g18716), .I1 (g4878), .I2 (g15915));
AN2X1 gate11197(.O (g31186), .I1 (g2375), .I2 (g30088));
AN2X1 gate11198(.O (g33186), .I1 (g32037), .I2 (g22830));
AN2X1 gate11199(.O (g24646), .I1 (g22640), .I2 (g19711));
AN2X1 gate11200(.O (g33676), .I1 (g33125), .I2 (g7970));
AN2X1 gate11201(.O (g33373), .I1 (g32288), .I2 (g21205));
AN2X1 gate11202(.O (g16516), .I1 (g5228), .I2 (g14627));
AN2X1 gate11203(.O (g27697), .I1 (g25785), .I2 (g23649));
AN2X1 gate11204(.O (g18582), .I1 (g2922), .I2 (g16349));
AN2X1 gate11205(.O (g27995), .I1 (g26809), .I2 (g23985));
AN2X1 gate11206(.O (g31654), .I1 (g29325), .I2 (g13062));
AN2X1 gate11207(.O (g30576), .I1 (g18898), .I2 (g29800));
AN2X1 gate11208(.O (g22127), .I1 (g6625), .I2 (g19277));
AN2X1 gate11209(.O (g34585), .I1 (g24705), .I2 (g34316));
AN2X1 gate11210(.O (g34484), .I1 (g34407), .I2 (g18939));
AN2X1 gate11211(.O (g18310), .I1 (g1333), .I2 (g16931));
AN2X1 gate11212(.O (g29601), .I1 (g1890), .I2 (g28955));
AN2X1 gate11213(.O (g31936), .I1 (g31213), .I2 (g24005));
AN2X1 gate11214(.O (g33417), .I1 (g32371), .I2 (g21424));
AN4X1 gate11215(.O (I31327), .I1 (g32928), .I2 (g32929), .I3 (g32930), .I4 (g32931));
AN2X1 gate11216(.O (g21789), .I1 (g3451), .I2 (g20391));
AN2X1 gate11217(.O (g26799), .I1 (g25247), .I2 (g21068));
AN2X1 gate11218(.O (g29975), .I1 (g28986), .I2 (g10420));
AN2X1 gate11219(.O (g34554), .I1 (g34347), .I2 (g20495));
AN2X1 gate11220(.O (g18627), .I1 (g15093), .I2 (g17093));
AN2X1 gate11221(.O (g15863), .I1 (g13762), .I2 (g13223));
AN2X1 gate11222(.O (g18379), .I1 (g1906), .I2 (g15171));
AN2X1 gate11223(.O (g30200), .I1 (g28665), .I2 (g23862));
AN2X1 gate11224(.O (g21788), .I1 (g3401), .I2 (g20391));
AN2X1 gate11225(.O (g33334), .I1 (g32219), .I2 (g20613));
AN2X1 gate11226(.O (g18112), .I1 (g182), .I2 (g17015));
AN2X1 gate11227(.O (g16422), .I1 (g8216), .I2 (g13627));
AN2X1 gate11228(.O (g23724), .I1 (g14767), .I2 (g21123));
AN2X1 gate11229(.O (g25852), .I1 (g4593), .I2 (g24411));
AN2X1 gate11230(.O (g18378), .I1 (g1932), .I2 (g15171));
AN2X1 gate11231(.O (g22103), .I1 (g15164), .I2 (g18833));
AN3X1 gate11232(.O (g34115), .I1 (g20516), .I2 (g9104), .I3 (g33750));
AN2X1 gate11233(.O (g21829), .I1 (g3770), .I2 (g20453));
AN2X1 gate11234(.O (g29937), .I1 (g13044), .I2 (g29196));
AN2X1 gate11235(.O (g14220), .I1 (g8612), .I2 (g11820));
AN2X1 gate11236(.O (g21920), .I1 (g5062), .I2 (g21468));
AN2X1 gate11237(.O (g23920), .I1 (g4135), .I2 (g19549));
AN2X1 gate11238(.O (g22095), .I1 (g6428), .I2 (g18833));
AN2X1 gate11239(.O (g16208), .I1 (g3965), .I2 (g14085));
AN2X1 gate11240(.O (g25963), .I1 (g1657), .I2 (g24978));
AN2X1 gate11241(.O (g28318), .I1 (g27233), .I2 (g19770));
AN2X1 gate11242(.O (g18386), .I1 (g1964), .I2 (g15171));
AN2X1 gate11243(.O (g30921), .I1 (g29900), .I2 (g24789));
AN2X1 gate11244(.O (g28227), .I1 (g9397), .I2 (g27583));
AN2X1 gate11245(.O (g21828), .I1 (g3767), .I2 (g20453));
AN2X1 gate11246(.O (g15703), .I1 (g452), .I2 (g13437));
AN2X1 gate11247(.O (g17784), .I1 (g1152), .I2 (g13215));
AN2X1 gate11248(.O (g23828), .I1 (g9104), .I2 (g19128));
AN2X1 gate11249(.O (g18603), .I1 (g3119), .I2 (g16987));
AN2X1 gate11250(.O (g21946), .I1 (g5252), .I2 (g18997));
AN2X1 gate11251(.O (g18742), .I1 (g5120), .I2 (g17847));
AN4X1 gate11252(.O (g27445), .I1 (g8038), .I2 (g26314), .I3 (g9187), .I4 (g504));
AN2X1 gate11253(.O (g33423), .I1 (g32225), .I2 (g29657));
AN2X1 gate11254(.O (g29884), .I1 (g2555), .I2 (g29153));
AN2X1 gate11255(.O (g23121), .I1 (g19128), .I2 (g9104));
AN2X1 gate11256(.O (g24229), .I1 (g896), .I2 (g22594));
AN2X1 gate11257(.O (g34745), .I1 (g34669), .I2 (g19482));
AN2X1 gate11258(.O (g27316), .I1 (g2407), .I2 (g26710));
AN2X1 gate11259(.O (g24228), .I1 (g862), .I2 (g22594));
AN2X1 gate11260(.O (g18681), .I1 (g4653), .I2 (g15885));
AN4X1 gate11261(.O (I31091), .I1 (g29385), .I2 (g32586), .I3 (g32587), .I4 (g32588));
AN2X1 gate11262(.O (g24011), .I1 (g7939), .I2 (g19524));
AN2X1 gate11263(.O (g32326), .I1 (g31317), .I2 (g23539));
AN2X1 gate11264(.O (g29666), .I1 (g28980), .I2 (g22498));
AN2X1 gate11265(.O (g17181), .I1 (g1945), .I2 (g13014));
AN2X1 gate11266(.O (g16614), .I1 (g5945), .I2 (g14933));
AN2X1 gate11267(.O (g17671), .I1 (g7685), .I2 (g13485));
AN2X1 gate11268(.O (g29363), .I1 (g8458), .I2 (g28444));
AN2X1 gate11269(.O (g23682), .I1 (g16970), .I2 (g20874));
AN2X1 gate11270(.O (g18802), .I1 (g6195), .I2 (g15348));
AN2X1 gate11271(.O (g18429), .I1 (g2193), .I2 (g18008));
AN2X1 gate11272(.O (g32040), .I1 (g14122), .I2 (g31243));
AN2X1 gate11273(.O (g24716), .I1 (g15935), .I2 (g23004));
AN4X1 gate11274(.O (I24680), .I1 (g24029), .I2 (g24030), .I3 (g24031), .I4 (g24032));
AN2X1 gate11275(.O (g33909), .I1 (g33131), .I2 (g10708));
AN2X1 gate11276(.O (g34184), .I1 (g33698), .I2 (g24388));
AN2X1 gate11277(.O (g18730), .I1 (g4950), .I2 (g16861));
AN2X1 gate11278(.O (g15821), .I1 (g3598), .I2 (g14110));
AN2X1 gate11279(.O (g27988), .I1 (g26781), .I2 (g23941));
AN2X1 gate11280(.O (g18793), .I1 (g6159), .I2 (g15348));
AN2X1 gate11281(.O (g18428), .I1 (g2169), .I2 (g18008));
AN2X1 gate11282(.O (g24582), .I1 (g5808), .I2 (g23402));
AN2X1 gate11283(.O (g33908), .I1 (g33092), .I2 (g18935));
AN3X1 gate11284(.O (g28281), .I1 (g7362), .I2 (g1936), .I3 (g27440));
AN2X1 gate11285(.O (g16593), .I1 (g5599), .I2 (g14885));
AN2X1 gate11286(.O (g12924), .I1 (g1570), .I2 (g10980));
AN2X1 gate11287(.O (g27432), .I1 (g26519), .I2 (g17582));
AN2X1 gate11288(.O (g13020), .I1 (g401), .I2 (g11048));
AN2X1 gate11289(.O (g18765), .I1 (g5489), .I2 (g17929));
AN2X1 gate11290(.O (g28301), .I1 (g27224), .I2 (g19750));
AN2X1 gate11291(.O (g24310), .I1 (g4495), .I2 (g22228));
AN2X1 gate11292(.O (g16122), .I1 (g9491), .I2 (g14291));
AN2X1 gate11293(.O (g18690), .I1 (g15130), .I2 (g16053));
AN4X1 gate11294(.O (g28739), .I1 (g21434), .I2 (g26424), .I3 (g25274), .I4 (g27395));
AN2X1 gate11295(.O (g18549), .I1 (g2799), .I2 (g15277));
AN2X1 gate11296(.O (g11046), .I1 (g9889), .I2 (g6120));
AN2X1 gate11297(.O (g25921), .I1 (g24936), .I2 (g9664));
AN2X1 gate11298(.O (g13046), .I1 (g6870), .I2 (g11270));
AN2X1 gate11299(.O (g26207), .I1 (g2638), .I2 (g25170));
AN2X1 gate11300(.O (g24627), .I1 (g22763), .I2 (g19679));
AN2X1 gate11301(.O (g29580), .I1 (g28519), .I2 (g14186));
AN2X1 gate11302(.O (g21760), .I1 (g3207), .I2 (g20785));
AN2X1 gate11303(.O (g20112), .I1 (g13540), .I2 (g16661));
AN2X1 gate11304(.O (g31242), .I1 (g29373), .I2 (g25409));
AN2X1 gate11305(.O (g22089), .I1 (g6311), .I2 (g19210));
AN2X1 gate11306(.O (g27461), .I1 (g26576), .I2 (g17611));
AN2X1 gate11307(.O (g33242), .I1 (g32123), .I2 (g19931));
AN2X1 gate11308(.O (g18548), .I1 (g2807), .I2 (g15277));
AN2X1 gate11309(.O (g15873), .I1 (g3550), .I2 (g14072));
AN2X1 gate11310(.O (g28645), .I1 (g27556), .I2 (g20599));
AN4X1 gate11311(.O (I31192), .I1 (g32733), .I2 (g32734), .I3 (g32735), .I4 (g32736));
AN2X1 gate11312(.O (g27342), .I1 (g12592), .I2 (g26792));
AN2X1 gate11313(.O (g24378), .I1 (g3106), .I2 (g22718));
AN2X1 gate11314(.O (g16641), .I1 (g6613), .I2 (g14782));
AN2X1 gate11315(.O (g27145), .I1 (g14121), .I2 (g26382));
AN2X1 gate11316(.O (g22088), .I1 (g6307), .I2 (g19210));
AN2X1 gate11317(.O (g18504), .I1 (g2579), .I2 (g15509));
AN2X1 gate11318(.O (g22024), .I1 (g5897), .I2 (g19147));
AN2X1 gate11319(.O (g31123), .I1 (g1834), .I2 (g29994));
AN2X1 gate11320(.O (g32183), .I1 (g2795), .I2 (g31653));
AN2X1 gate11321(.O (g19266), .I1 (g246), .I2 (g16214));
AN2X1 gate11322(.O (g33814), .I1 (g33098), .I2 (g28144));
AN2X1 gate11323(.O (g28290), .I1 (g23780), .I2 (g27759));
AN2X1 gate11324(.O (g32397), .I1 (g31068), .I2 (g15830));
AN2X1 gate11325(.O (g13282), .I1 (g3546), .I2 (g11480));
AN2X1 gate11326(.O (g27650), .I1 (g26519), .I2 (g15479));
AN4X1 gate11327(.O (g29110), .I1 (g27187), .I2 (g12687), .I3 (g20751), .I4 (I27429));
AN2X1 gate11328(.O (g25973), .I1 (g2342), .I2 (g24994));
AN2X1 gate11329(.O (g18317), .I1 (g12846), .I2 (g17873));
AN2X1 gate11330(.O (g33807), .I1 (g33112), .I2 (g25452));
AN2X1 gate11331(.O (g31974), .I1 (g31760), .I2 (g22176));
AN2X1 gate11332(.O (g29321), .I1 (g29033), .I2 (g22148));
AN2X1 gate11333(.O (g33639), .I1 (g33386), .I2 (g18829));
AN4X1 gate11334(.O (g26241), .I1 (g24688), .I2 (g10678), .I3 (g8778), .I4 (g10627));
AN2X1 gate11335(.O (g34214), .I1 (g33772), .I2 (g22689));
AN2X1 gate11336(.O (g29531), .I1 (g1664), .I2 (g28559));
AN2X1 gate11337(.O (g31230), .I1 (g30285), .I2 (g20751));
AN2X1 gate11338(.O (g18129), .I1 (g518), .I2 (g16971));
AN2X1 gate11339(.O (g30207), .I1 (g28680), .I2 (g23874));
AN2X1 gate11340(.O (g16635), .I1 (g5607), .I2 (g14959));
AN2X1 gate11341(.O (g27696), .I1 (g25800), .I2 (g23647));
AN2X1 gate11342(.O (g34329), .I1 (g14511), .I2 (g34181));
AN2X1 gate11343(.O (g27330), .I1 (g2541), .I2 (g26744));
AN2X1 gate11344(.O (g27393), .I1 (g26099), .I2 (g20066));
AN2X1 gate11345(.O (g28427), .I1 (g27258), .I2 (g20008));
AN2X1 gate11346(.O (g24681), .I1 (g16653), .I2 (g22988));
AN2X1 gate11347(.O (g29178), .I1 (g27163), .I2 (g12687));
AN2X1 gate11348(.O (g29740), .I1 (g2648), .I2 (g29154));
AN2X1 gate11349(.O (g30005), .I1 (g28230), .I2 (g24394));
AN2X1 gate11350(.O (g22126), .I1 (g6621), .I2 (g19277));
AN2X1 gate11351(.O (g18128), .I1 (g504), .I2 (g16971));
AN2X1 gate11352(.O (g21927), .I1 (g5164), .I2 (g18997));
AN2X1 gate11353(.O (g26100), .I1 (g1677), .I2 (g25097));
AN2X1 gate11354(.O (g19588), .I1 (g3849), .I2 (g16853));
AN2X1 gate11355(.O (g33416), .I1 (g32370), .I2 (g21423));
AN2X1 gate11356(.O (g29685), .I1 (g2084), .I2 (g28711));
AN4X1 gate11357(.O (I31326), .I1 (g30735), .I2 (g31853), .I3 (g32926), .I4 (g32927));
AN2X1 gate11358(.O (g18245), .I1 (g1193), .I2 (g16431));
AN2X1 gate11359(.O (g27132), .I1 (g26055), .I2 (g16589));
AN2X1 gate11360(.O (g34538), .I1 (g34330), .I2 (g20054));
AN2X1 gate11361(.O (g18626), .I1 (g3498), .I2 (g17062));
AN2X1 gate11362(.O (g15913), .I1 (g3933), .I2 (g14021));
AN2X1 gate11363(.O (g24730), .I1 (g6177), .I2 (g23699));
AN2X1 gate11364(.O (g31992), .I1 (g31773), .I2 (g22213));
AN2X1 gate11365(.O (g18323), .I1 (g1632), .I2 (g17873));
AN2X1 gate11366(.O (g33841), .I1 (g33254), .I2 (g20268));
AN2X1 gate11367(.O (g18299), .I1 (g1526), .I2 (g16489));
AN2X1 gate11368(.O (g18533), .I1 (g2729), .I2 (g15277));
AN2X1 gate11369(.O (g28547), .I1 (g6821), .I2 (g27091));
AN3X1 gate11370(.O (g33510), .I1 (g32816), .I2 (I31246), .I3 (I31247));
AN2X1 gate11371(.O (g24765), .I1 (g17699), .I2 (g22498));
AN2X1 gate11372(.O (g18298), .I1 (g15073), .I2 (g16489));
AN3X1 gate11373(.O (g27161), .I1 (g26166), .I2 (g8241), .I3 (g1783));
AN2X1 gate11374(.O (g30241), .I1 (g28729), .I2 (g23926));
AN4X1 gate11375(.O (I31252), .I1 (g32819), .I2 (g32820), .I3 (g32821), .I4 (g32822));
AN2X1 gate11376(.O (g31579), .I1 (g19128), .I2 (g29814));
AN2X1 gate11377(.O (g18775), .I1 (g7028), .I2 (g15615));
AN2X1 gate11378(.O (g24549), .I1 (g23162), .I2 (g20887));
AN2X1 gate11379(.O (g28226), .I1 (g27825), .I2 (g26667));
AN2X1 gate11380(.O (g21755), .I1 (g3203), .I2 (g20785));
AN2X1 gate11381(.O (g29334), .I1 (g29148), .I2 (g18908));
AN2X1 gate11382(.O (g16474), .I1 (g8280), .I2 (g13666));
AN2X1 gate11383(.O (g23755), .I1 (g14821), .I2 (g21204));
AN2X1 gate11384(.O (g27259), .I1 (g26755), .I2 (g26725));
AN2X1 gate11385(.O (g19749), .I1 (g732), .I2 (g16646));
AN2X1 gate11386(.O (g32047), .I1 (g27248), .I2 (g31070));
AN2X1 gate11387(.O (g33835), .I1 (g4340), .I2 (g33413));
AN2X1 gate11388(.O (g9968), .I1 (g1339), .I2 (g1500));
AN2X1 gate11389(.O (g21770), .I1 (g3251), .I2 (g20785));
AN2X1 gate11390(.O (g32205), .I1 (g30922), .I2 (g28463));
AN2X1 gate11391(.O (g21981), .I1 (g5543), .I2 (g19074));
AN2X1 gate11392(.O (g22060), .I1 (g6151), .I2 (g21611));
AN2X1 gate11393(.O (g10902), .I1 (g7858), .I2 (g1129));
AN2X1 gate11394(.O (g18737), .I1 (g4975), .I2 (g16826));
AN2X1 gate11395(.O (g27087), .I1 (g13872), .I2 (g26284));
AN2X1 gate11396(.O (g28572), .I1 (g27829), .I2 (g15669));
AN2X1 gate11397(.O (g12259), .I1 (g9480), .I2 (g640));
AN2X1 gate11398(.O (g24504), .I1 (g22226), .I2 (g19410));
AN2X1 gate11399(.O (g32311), .I1 (g31295), .I2 (g20582));
AN2X1 gate11400(.O (g25207), .I1 (g22513), .I2 (g10621));
AN2X1 gate11401(.O (g29762), .I1 (g28298), .I2 (g10233));
AN2X1 gate11402(.O (g18232), .I1 (g1124), .I2 (g16326));
AN2X1 gate11403(.O (g34771), .I1 (g34693), .I2 (g20147));
AN2X1 gate11404(.O (g29964), .I1 (g2008), .I2 (g28830));
AN2X1 gate11405(.O (g16537), .I1 (g5937), .I2 (g14855));
AN2X1 gate11406(.O (g11027), .I1 (g5097), .I2 (g9724));
AN2X1 gate11407(.O (g30235), .I1 (g28723), .I2 (g23915));
AN3X1 gate11408(.O (I18713), .I1 (g13156), .I2 (g6767), .I3 (g6756));
AN3X1 gate11409(.O (g25328), .I1 (g5022), .I2 (g23764), .I3 (I24505));
AN2X1 gate11410(.O (g11890), .I1 (g7499), .I2 (g9155));
AN2X1 gate11411(.O (g24317), .I1 (g4534), .I2 (g22228));
AN2X1 gate11412(.O (g15797), .I1 (g3909), .I2 (g14139));
AN2X1 gate11413(.O (g18697), .I1 (g4749), .I2 (g16777));
AN2X1 gate11414(.O (g27043), .I1 (g26335), .I2 (g8632));
AN2X1 gate11415(.O (g32051), .I1 (g31506), .I2 (g10831));
AN4X1 gate11416(.O (g16283), .I1 (g11547), .I2 (g11592), .I3 (g6789), .I4 (I17606));
AN2X1 gate11417(.O (g29587), .I1 (g2181), .I2 (g28935));
AN4X1 gate11418(.O (I31062), .I1 (g32545), .I2 (g32546), .I3 (g32547), .I4 (g32548));
AN2X1 gate11419(.O (g18261), .I1 (g1256), .I2 (g16000));
AN2X1 gate11420(.O (g21767), .I1 (g3239), .I2 (g20785));
AN2X1 gate11421(.O (g21794), .I1 (g15094), .I2 (g20924));
AN2X1 gate11422(.O (g21845), .I1 (g3881), .I2 (g21070));
AN2X1 gate11423(.O (g12043), .I1 (g1345), .I2 (g7601));
AN2X1 gate11424(.O (g16303), .I1 (g4527), .I2 (g12921));
AN2X1 gate11425(.O (g10290), .I1 (g4358), .I2 (g4349));
AN2X1 gate11426(.O (g24002), .I1 (g19613), .I2 (g10971));
AN2X1 gate11427(.O (g21990), .I1 (g5591), .I2 (g19074));
AN2X1 gate11428(.O (g11003), .I1 (g7880), .I2 (g1300));
AN2X1 gate11429(.O (g18512), .I1 (g2619), .I2 (g15509));
AN2X1 gate11430(.O (g23990), .I1 (g19610), .I2 (g10951));
AN4X1 gate11431(.O (I27524), .I1 (g28037), .I2 (g24114), .I3 (g24115), .I4 (g24116));
AN2X1 gate11432(.O (g33720), .I1 (g33161), .I2 (g19439));
AN3X1 gate11433(.O (g19560), .I1 (g15832), .I2 (g1157), .I3 (g10893));
AN2X1 gate11434(.O (g29909), .I1 (g28435), .I2 (g23388));
AN4X1 gate11435(.O (g27602), .I1 (g23032), .I2 (g26244), .I3 (g26424), .I4 (g24966));
AN2X1 gate11436(.O (g31275), .I1 (g30147), .I2 (g27800));
AN2X1 gate11437(.O (g34515), .I1 (g34288), .I2 (g19491));
AN2X1 gate11438(.O (g34414), .I1 (g34206), .I2 (g21457));
AN4X1 gate11439(.O (g28889), .I1 (g17292), .I2 (g25169), .I3 (g26424), .I4 (g27395));
AN2X1 gate11440(.O (g31746), .I1 (g30093), .I2 (g23905));
AN2X1 gate11441(.O (g27375), .I1 (g26519), .I2 (g17479));
AN2X1 gate11442(.O (g26206), .I1 (g2523), .I2 (g25495));
AN2X1 gate11443(.O (g31493), .I1 (g29791), .I2 (g23434));
AN2X1 gate11444(.O (g32350), .I1 (g2697), .I2 (g31710));
AN2X1 gate11445(.O (g21719), .I1 (g358), .I2 (g21037));
AN3X1 gate11446(.O (g33493), .I1 (g32693), .I2 (I31161), .I3 (I31162));
AN2X1 gate11447(.O (g24323), .I1 (g4546), .I2 (g22228));
AN2X1 gate11448(.O (g24299), .I1 (g4456), .I2 (g22550));
AN2X1 gate11449(.O (g13778), .I1 (g4540), .I2 (g10597));
AN2X1 gate11450(.O (g13081), .I1 (g8626), .I2 (g11122));
AN2X1 gate11451(.O (g29569), .I1 (g29028), .I2 (g22498));
AN2X1 gate11452(.O (g21718), .I1 (g370), .I2 (g21037));
AN3X1 gate11453(.O (g33465), .I1 (g32491), .I2 (I31021), .I3 (I31022));
AN2X1 gate11454(.O (g31237), .I1 (g29366), .I2 (g25325));
AN3X1 gate11455(.O (g10632), .I1 (g7475), .I2 (g7441), .I3 (g890));
AN2X1 gate11456(.O (g24298), .I1 (g4392), .I2 (g22550));
AN2X1 gate11457(.O (g33237), .I1 (g32394), .I2 (g25198));
AN2X1 gate11458(.O (g32152), .I1 (g31631), .I2 (g29998));
AN2X1 gate11459(.O (g18445), .I1 (g2273), .I2 (g18008));
AN2X1 gate11460(.O (g24775), .I1 (g17594), .I2 (g22498));
AN2X1 gate11461(.O (g29568), .I1 (g2571), .I2 (g28950));
AN2X1 gate11462(.O (g29747), .I1 (g28286), .I2 (g23196));
AN2X1 gate11463(.O (g32396), .I1 (g4698), .I2 (g30983));
AN2X1 gate11464(.O (g33340), .I1 (g32222), .I2 (g20639));
AN2X1 gate11465(.O (g21832), .I1 (g3787), .I2 (g20453));
AN2X1 gate11466(.O (g18499), .I1 (g2476), .I2 (g15426));
AN2X1 gate11467(.O (g18316), .I1 (g1564), .I2 (g16931));
AN2X1 gate11468(.O (g33684), .I1 (g33139), .I2 (g13565));
AN2X1 gate11469(.O (g16840), .I1 (g5467), .I2 (g14262));
AN2X1 gate11470(.O (g31142), .I1 (g2527), .I2 (g30039));
AN2X1 gate11471(.O (g22055), .I1 (g6128), .I2 (g21611));
AN2X1 gate11472(.O (g18498), .I1 (g2547), .I2 (g15426));
AN2X1 gate11473(.O (g32413), .I1 (g31121), .I2 (g19518));
AN2X1 gate11474(.O (g19693), .I1 (g6181), .I2 (g17087));
AN2X1 gate11475(.O (g22111), .I1 (g6549), .I2 (g19277));
AN4X1 gate11476(.O (I31047), .I1 (g32524), .I2 (g32525), .I3 (g32526), .I4 (g32527));
AN2X1 gate11477(.O (g21861), .I1 (g3949), .I2 (g21070));
AN2X1 gate11478(.O (g34584), .I1 (g24653), .I2 (g34315));
AN2X1 gate11479(.O (g22070), .I1 (g6243), .I2 (g19210));
AN2X1 gate11480(.O (g13998), .I1 (g6589), .I2 (g12629));
AN2X1 gate11481(.O (g31517), .I1 (g29849), .I2 (g23482));
AN2X1 gate11482(.O (g26345), .I1 (g13051), .I2 (g25505));
AN2X1 gate11483(.O (g28426), .I1 (g27257), .I2 (g20006));
AN3X1 gate11484(.O (g33517), .I1 (g32867), .I2 (I31281), .I3 (I31282));
AN2X1 gate11485(.O (g29751), .I1 (g28297), .I2 (g23216));
AN2X1 gate11486(.O (g29807), .I1 (g28359), .I2 (g23272));
AN4X1 gate11487(.O (I31311), .I1 (g30673), .I2 (g31851), .I3 (g32903), .I4 (g32904));
AN2X1 gate11488(.O (g29772), .I1 (g28323), .I2 (g23243));
AN2X1 gate11489(.O (g22590), .I1 (g19274), .I2 (g19452));
AN2X1 gate11490(.O (g16192), .I1 (g6191), .I2 (g14321));
AN2X1 gate11491(.O (g26849), .I1 (g2994), .I2 (g24527));
AN2X1 gate11492(.O (g29974), .I1 (g29173), .I2 (g12914));
AN2X1 gate11493(.O (g15711), .I1 (g460), .I2 (g13437));
AN2X1 gate11494(.O (g18611), .I1 (g15090), .I2 (g17200));
AN2X1 gate11495(.O (g27459), .I1 (g26549), .I2 (g17609));
AN2X1 gate11496(.O (g21926), .I1 (g15147), .I2 (g18997));
AN2X1 gate11497(.O (g18722), .I1 (g4917), .I2 (g16077));
AN2X1 gate11498(.O (g26399), .I1 (g15572), .I2 (g25566));
AN3X1 gate11499(.O (g25414), .I1 (g5406), .I2 (g22194), .I3 (I24549));
AN2X1 gate11500(.O (g25991), .I1 (g2060), .I2 (g25023));
AN2X1 gate11501(.O (g23389), .I1 (g9072), .I2 (g19757));
AN2X1 gate11502(.O (g29639), .I1 (g28510), .I2 (g11618));
AN2X1 gate11503(.O (g15109), .I1 (g4269), .I2 (g14454));
AN2X1 gate11504(.O (g26848), .I1 (g2950), .I2 (g24526));
AN3X1 gate11505(.O (I16646), .I1 (g10160), .I2 (g12413), .I3 (g12343));
AN2X1 gate11506(.O (g26398), .I1 (g24946), .I2 (g10474));
AN3X1 gate11507(.O (g22384), .I1 (g9354), .I2 (g9285), .I3 (g20784));
AN2X1 gate11508(.O (g18432), .I1 (g2223), .I2 (g18008));
AN4X1 gate11509(.O (I24705), .I1 (g24064), .I2 (g24065), .I3 (g24066), .I4 (g24067));
AN2X1 gate11510(.O (g29638), .I1 (g2583), .I2 (g29025));
AN4X1 gate11511(.O (I31051), .I1 (g31376), .I2 (g31804), .I3 (g32529), .I4 (g32530));
AN2X1 gate11512(.O (g21701), .I1 (g153), .I2 (g20283));
AN4X1 gate11513(.O (I31072), .I1 (g32559), .I2 (g32560), .I3 (g32561), .I4 (g32562));
AN2X1 gate11514(.O (g18271), .I1 (g1296), .I2 (g16031));
AN2X1 gate11515(.O (g30082), .I1 (g29181), .I2 (g12752));
AN2X1 gate11516(.O (g34114), .I1 (g33920), .I2 (g23742));
AN2X1 gate11517(.O (g15108), .I1 (g4264), .I2 (g14454));
AN2X1 gate11518(.O (g21777), .I1 (g3380), .I2 (g20391));
AN2X1 gate11519(.O (g34758), .I1 (g34683), .I2 (g19657));
AN2X1 gate11520(.O (g26652), .I1 (g10799), .I2 (g24426));
AN2X1 gate11521(.O (g31130), .I1 (g12191), .I2 (g30019));
AN2X1 gate11522(.O (g22067), .I1 (g6215), .I2 (g19210));
AN2X1 gate11523(.O (g22094), .I1 (g6398), .I2 (g18833));
AN2X1 gate11524(.O (g34082), .I1 (g33709), .I2 (g19554));
AN2X1 gate11525(.O (g30107), .I1 (g28560), .I2 (g20909));
AN2X1 gate11526(.O (g21251), .I1 (g13969), .I2 (g17470));
AN4X1 gate11527(.O (I24679), .I1 (g19968), .I2 (g24026), .I3 (g24027), .I4 (g24028));
AN2X1 gate11528(.O (g33362), .I1 (g32259), .I2 (g20914));
AN2X1 gate11529(.O (g11449), .I1 (g6052), .I2 (g7175));
AN2X1 gate11530(.O (g27545), .I1 (g26519), .I2 (g17756));
AN2X1 gate11531(.O (g16483), .I1 (g5224), .I2 (g14915));
AN2X1 gate11532(.O (g18753), .I1 (g15148), .I2 (g15595));
AN2X1 gate11533(.O (g18461), .I1 (g2307), .I2 (g15224));
AN2X1 gate11534(.O (g31523), .I1 (g7528), .I2 (g29333));
AN2X1 gate11535(.O (g32020), .I1 (g4157), .I2 (g30937));
AN2X1 gate11536(.O (g18342), .I1 (g1592), .I2 (g17873));
AN3X1 gate11537(.O (g33523), .I1 (g32909), .I2 (I31311), .I3 (I31312));
AN2X1 gate11538(.O (g29841), .I1 (g28371), .I2 (g23283));
AN2X1 gate11539(.O (g19914), .I1 (g2815), .I2 (g15853));
AN2X1 gate11540(.O (g29992), .I1 (g29012), .I2 (g10490));
AN2X1 gate11541(.O (g27599), .I1 (g26337), .I2 (g20033));
AN2X1 gate11542(.O (g34744), .I1 (g34668), .I2 (g19481));
AN2X1 gate11543(.O (g18145), .I1 (g582), .I2 (g17533));
AN2X1 gate11544(.O (g29510), .I1 (g28856), .I2 (g22342));
AN2X1 gate11545(.O (g32046), .I1 (g10925), .I2 (g30735));
AN2X1 gate11546(.O (g18199), .I1 (g832), .I2 (g17821));
AN2X1 gate11547(.O (g22019), .I1 (g5857), .I2 (g19147));
AN2X1 gate11548(.O (g27598), .I1 (g25899), .I2 (g10475));
AN2X1 gate11549(.O (g18650), .I1 (g6928), .I2 (g17271));
AN2X1 gate11550(.O (g18736), .I1 (g4991), .I2 (g16826));
AN2X1 gate11551(.O (g27086), .I1 (g25836), .I2 (g22495));
AN2X1 gate11552(.O (g31475), .I1 (g29756), .I2 (g23406));
AN2X1 gate11553(.O (g29579), .I1 (g28457), .I2 (g7964));
AN2X1 gate11554(.O (g17150), .I1 (g8579), .I2 (g12995));
AN3X1 gate11555(.O (I24030), .I1 (g8390), .I2 (g8016), .I3 (g3396));
AN3X1 gate11556(.O (g33475), .I1 (g32563), .I2 (I31071), .I3 (I31072));
AN2X1 gate11557(.O (g16536), .I1 (g5917), .I2 (g14996));
AN2X1 gate11558(.O (g18198), .I1 (g15059), .I2 (g17821));
AN2X1 gate11559(.O (g22018), .I1 (g15157), .I2 (g19147));
AN2X1 gate11560(.O (g18529), .I1 (g2712), .I2 (g15277));
AN2X1 gate11561(.O (g21997), .I1 (g5619), .I2 (g19074));
AN2X1 gate11562(.O (g32113), .I1 (g31601), .I2 (g29925));
AN2X1 gate11563(.O (g34398), .I1 (g7684), .I2 (g34070));
AN4X1 gate11564(.O (I31152), .I1 (g32675), .I2 (g32676), .I3 (g32677), .I4 (g32678));
AN2X1 gate11565(.O (g33727), .I1 (g33115), .I2 (g19499));
AN2X1 gate11566(.O (g24499), .I1 (g22217), .I2 (g19394));
AN2X1 gate11567(.O (g29578), .I1 (g2491), .I2 (g28606));
AN2X1 gate11568(.O (g33863), .I1 (g33273), .I2 (g20505));
AN2X1 gate11569(.O (g19594), .I1 (g11913), .I2 (g17268));
AN2X1 gate11570(.O (g29835), .I1 (g28326), .I2 (g24866));
AN2X1 gate11571(.O (g34141), .I1 (g33932), .I2 (g23828));
AN2X1 gate11572(.O (g16702), .I1 (g5615), .I2 (g14691));
AN2X1 gate11573(.O (g24316), .I1 (g4527), .I2 (g22228));
AN2X1 gate11574(.O (g31222), .I1 (g2643), .I2 (g30113));
AN2X1 gate11575(.O (g32282), .I1 (g31258), .I2 (g20503));
AN4X1 gate11576(.O (g27817), .I1 (g22498), .I2 (g25245), .I3 (g26424), .I4 (g26236));
AN2X1 gate11577(.O (g15796), .I1 (g3586), .I2 (g14015));
AN2X1 gate11578(.O (g18696), .I1 (g4741), .I2 (g16053));
AN2X1 gate11579(.O (g18330), .I1 (g1668), .I2 (g17873));
AN2X1 gate11580(.O (g32302), .I1 (g31279), .I2 (g23485));
AN2X1 gate11581(.O (g18393), .I1 (g1917), .I2 (g15171));
AN2X1 gate11582(.O (g24498), .I1 (g14036), .I2 (g23850));
AN2X1 gate11583(.O (g29586), .I1 (g1886), .I2 (g28927));
AN2X1 gate11584(.O (g16621), .I1 (g8278), .I2 (g13821));
AN2X1 gate11585(.O (g12817), .I1 (g1351), .I2 (g7601));
AN2X1 gate11586(.O (g21766), .I1 (g3235), .I2 (g20785));
AN2X1 gate11587(.O (g26833), .I1 (g2852), .I2 (g24509));
AN2X1 gate11588(.O (g26049), .I1 (g9621), .I2 (g25046));
AN2X1 gate11589(.O (g30263), .I1 (g28773), .I2 (g23962));
AN2X1 gate11590(.O (g32105), .I1 (g4922), .I2 (g30673));
AN2X1 gate11591(.O (g28658), .I1 (g27563), .I2 (g20611));
AN2X1 gate11592(.O (g18764), .I1 (g5485), .I2 (g17929));
AN4X1 gate11593(.O (g20056), .I1 (g16291), .I2 (g9007), .I3 (g8954), .I4 (g8903));
AN2X1 gate11594(.O (g18365), .I1 (g1848), .I2 (g17955));
AN2X1 gate11595(.O (g27158), .I1 (g26609), .I2 (g16645));
AN2X1 gate11596(.O (g21871), .I1 (g4108), .I2 (g19801));
AN2X1 gate11597(.O (g25107), .I1 (g17643), .I2 (g23508));
AN3X1 gate11598(.O (g22457), .I1 (g7753), .I2 (g7717), .I3 (g21288));
AN2X1 gate11599(.O (g15840), .I1 (g3949), .I2 (g14142));
AN2X1 gate11600(.O (g18132), .I1 (g513), .I2 (g16971));
AN2X1 gate11601(.O (g26048), .I1 (g5853), .I2 (g25044));
AN2X1 gate11602(.O (g28339), .I1 (g9946), .I2 (g27693));
AN2X1 gate11603(.O (g30135), .I1 (g28592), .I2 (g21180));
AN2X1 gate11604(.O (g24722), .I1 (g17618), .I2 (g22417));
AN2X1 gate11605(.O (g34135), .I1 (g33926), .I2 (g23802));
AN3X1 gate11606(.O (I18782), .I1 (g13156), .I2 (g11450), .I3 (g6756));
AN2X1 gate11607(.O (g7948), .I1 (g1548), .I2 (g1430));
AN2X1 gate11608(.O (g29615), .I1 (g1844), .I2 (g29049));
AN2X1 gate11609(.O (g16673), .I1 (g6617), .I2 (g14822));
AN2X1 gate11610(.O (g18161), .I1 (g691), .I2 (g17433));
AN2X1 gate11611(.O (g34962), .I1 (g34945), .I2 (g23020));
AN2X1 gate11612(.O (g19637), .I1 (g5142), .I2 (g16958));
AN2X1 gate11613(.O (g26613), .I1 (g1361), .I2 (g24518));
AN2X1 gate11614(.O (g18709), .I1 (g59), .I2 (g17302));
AN2X1 gate11615(.O (g22001), .I1 (g5731), .I2 (g21562));
AN2X1 gate11616(.O (g22077), .I1 (g6263), .I2 (g19210));
AN2X1 gate11617(.O (g25848), .I1 (g25539), .I2 (g18977));
AN2X1 gate11618(.O (g14190), .I1 (g859), .I2 (g10632));
AN2X1 gate11619(.O (g27336), .I1 (g2675), .I2 (g26777));
AN2X1 gate11620(.O (g30049), .I1 (g13114), .I2 (g28167));
AN2X1 gate11621(.O (g18259), .I1 (g15068), .I2 (g16000));
AN2X1 gate11622(.O (g29746), .I1 (g28279), .I2 (g20037));
AN2X1 gate11623(.O (g34500), .I1 (g34276), .I2 (g30568));
AN2X1 gate11624(.O (g18225), .I1 (g1041), .I2 (g16100));
AN2X1 gate11625(.O (g33351), .I1 (g32236), .I2 (g20707));
AN2X1 gate11626(.O (g33372), .I1 (g32285), .I2 (g21183));
AN2X1 gate11627(.O (g18708), .I1 (g4818), .I2 (g16782));
AN2X1 gate11628(.O (g28197), .I1 (g27647), .I2 (g11344));
AN2X1 gate11629(.O (g25804), .I1 (g8069), .I2 (g24587));
AN2X1 gate11630(.O (g18471), .I1 (g2407), .I2 (g15224));
AN2X1 gate11631(.O (g33821), .I1 (g33238), .I2 (g20153));
AN2X1 gate11632(.O (g26273), .I1 (g2122), .I2 (g25389));
AN2X1 gate11633(.O (g30048), .I1 (g29193), .I2 (g12945));
AN2X1 gate11634(.O (g22689), .I1 (g18918), .I2 (g9104));
AN2X1 gate11635(.O (g18258), .I1 (g1221), .I2 (g16897));
AN2X1 gate11636(.O (g16634), .I1 (g5264), .I2 (g14953));
AN2X1 gate11637(.O (g20887), .I1 (g16282), .I2 (g4864));
AN2X1 gate11638(.O (g23451), .I1 (g13805), .I2 (g20510));
AN2X1 gate11639(.O (g24199), .I1 (g355), .I2 (g22722));
AN2X1 gate11640(.O (g24650), .I1 (g22641), .I2 (g19718));
AN2X1 gate11641(.O (g23220), .I1 (g19417), .I2 (g20067));
AN3X1 gate11642(.O (g24887), .I1 (g3712), .I2 (g23239), .I3 (I24054));
AN2X1 gate11643(.O (g30004), .I1 (g28521), .I2 (g25837));
AN4X1 gate11644(.O (I31046), .I1 (g29385), .I2 (g32521), .I3 (g32522), .I4 (g32523));
AN2X1 gate11645(.O (g22624), .I1 (g19344), .I2 (g19471));
AN2X1 gate11646(.O (g21911), .I1 (g5046), .I2 (g21468));
AN2X1 gate11647(.O (g30221), .I1 (g28700), .I2 (g23893));
AN2X1 gate11648(.O (g31790), .I1 (g21299), .I2 (g29385));
AN2X1 gate11649(.O (g33264), .I1 (g31965), .I2 (g21306));
AN2X1 gate11650(.O (g31516), .I1 (g29848), .I2 (g23476));
AN2X1 gate11651(.O (g24198), .I1 (g351), .I2 (g22722));
AN2X1 gate11652(.O (g33790), .I1 (g33108), .I2 (g20643));
AN3X1 gate11653(.O (g33516), .I1 (g32860), .I2 (I31276), .I3 (I31277));
AN2X1 gate11654(.O (g29806), .I1 (g28358), .I2 (g23271));
AN2X1 gate11655(.O (g29684), .I1 (g1982), .I2 (g29085));
AN2X1 gate11656(.O (g18244), .I1 (g1171), .I2 (g16431));
AN2X1 gate11657(.O (g26234), .I1 (g2657), .I2 (g25514));
AN2X1 gate11658(.O (g22102), .I1 (g6479), .I2 (g18833));
AN3X1 gate11659(.O (g24843), .I1 (g3010), .I2 (g23211), .I3 (I24015));
AN2X1 gate11660(.O (g33873), .I1 (g33291), .I2 (g20549));
AN2X1 gate11661(.O (g24330), .I1 (g18661), .I2 (g22228));
AN2X1 gate11662(.O (g22157), .I1 (g14608), .I2 (g18892));
AN2X1 gate11663(.O (g24393), .I1 (g3808), .I2 (g22844));
AN3X1 gate11664(.O (I24075), .I1 (g3736), .I2 (g3742), .I3 (g8553));
AN4X1 gate11665(.O (I31282), .I1 (g32863), .I2 (g32864), .I3 (g32865), .I4 (g32866));
AN2X1 gate11666(.O (g25962), .I1 (g9258), .I2 (g24971));
AN4X1 gate11667(.O (g16213), .I1 (g6772), .I2 (g6782), .I3 (g11640), .I4 (I17552));
AN2X1 gate11668(.O (g24764), .I1 (g17570), .I2 (g22472));
AN2X1 gate11669(.O (g29517), .I1 (g1870), .I2 (g28827));
AN4X1 gate11670(.O (I31302), .I1 (g32891), .I2 (g32892), .I3 (g32893), .I4 (g32894));
AN4X1 gate11671(.O (I31357), .I1 (g32970), .I2 (g32971), .I3 (g32972), .I4 (g32973));
AN2X1 gate11672(.O (g21776), .I1 (g3376), .I2 (g20391));
AN2X1 gate11673(.O (g21785), .I1 (g3431), .I2 (g20391));
AN4X1 gate11674(.O (I27519), .I1 (g28036), .I2 (g24107), .I3 (g24108), .I4 (g24109));
AN2X1 gate11675(.O (g18602), .I1 (g3115), .I2 (g16987));
AN2X1 gate11676(.O (g18810), .I1 (g6505), .I2 (g15483));
AN2X1 gate11677(.O (g15757), .I1 (g3207), .I2 (g14066));
AN2X1 gate11678(.O (g18657), .I1 (g4308), .I2 (g17128));
AN2X1 gate11679(.O (g22066), .I1 (g6209), .I2 (g19210));
AN2X1 gate11680(.O (g18774), .I1 (g5698), .I2 (g15615));
AN2X1 gate11681(.O (g7918), .I1 (g1205), .I2 (g1087));
AN2X1 gate11682(.O (g18375), .I1 (g1902), .I2 (g15171));
AN2X1 gate11683(.O (g31209), .I1 (g2084), .I2 (g30097));
AN2X1 gate11684(.O (g33422), .I1 (g32375), .I2 (g21456));
AN2X1 gate11685(.O (g34106), .I1 (g33917), .I2 (g23675));
AN2X1 gate11686(.O (g32248), .I1 (g31616), .I2 (g30299));
AN2X1 gate11687(.O (g21754), .I1 (g3195), .I2 (g20785));
AN4X1 gate11688(.O (I27518), .I1 (g20720), .I2 (g24104), .I3 (g24105), .I4 (g24106));
AN2X1 gate11689(.O (g10625), .I1 (g3431), .I2 (g7926));
AN2X1 gate11690(.O (g27309), .I1 (g26603), .I2 (g23057));
AN2X1 gate11691(.O (g23754), .I1 (g14816), .I2 (g21189));
AN2X1 gate11692(.O (g28714), .I1 (g27591), .I2 (g20711));
AN3X1 gate11693(.O (g16047), .I1 (g13322), .I2 (g1500), .I3 (g10699));
AN2X1 gate11694(.O (g25833), .I1 (g8228), .I2 (g24626));
AN2X1 gate11695(.O (g14126), .I1 (g881), .I2 (g10632));
AN4X1 gate11696(.O (g16205), .I1 (g11547), .I2 (g6782), .I3 (g11640), .I4 (I17542));
AN2X1 gate11697(.O (g27288), .I1 (g26515), .I2 (g23013));
AN2X1 gate11698(.O (g28315), .I1 (g27232), .I2 (g19769));
AN2X1 gate11699(.O (g33834), .I1 (g33095), .I2 (g29172));
AN2X1 gate11700(.O (g31208), .I1 (g30262), .I2 (g25188));
AN2X1 gate11701(.O (g32204), .I1 (g4245), .I2 (g31327));
AN2X1 gate11702(.O (g21859), .I1 (g3941), .I2 (g21070));
AN2X1 gate11703(.O (g21825), .I1 (g3736), .I2 (g20453));
AN2X1 gate11704(.O (g21950), .I1 (g5268), .I2 (g18997));
AN2X1 gate11705(.O (g26514), .I1 (g7400), .I2 (g25564));
AN2X1 gate11706(.O (g22876), .I1 (g20136), .I2 (g9104));
AN2X1 gate11707(.O (g18337), .I1 (g1706), .I2 (g17873));
AN2X1 gate11708(.O (g28202), .I1 (g27659), .I2 (g11413));
AN2X1 gate11709(.O (g30033), .I1 (g29189), .I2 (g12937));
AN2X1 gate11710(.O (g28257), .I1 (g27179), .I2 (g19686));
AN2X1 gate11711(.O (g21858), .I1 (g3937), .I2 (g21070));
AN2X1 gate11712(.O (g29362), .I1 (g27379), .I2 (g28307));
AN2X1 gate11713(.O (g18171), .I1 (g728), .I2 (g17433));
AN2X1 gate11714(.O (g30234), .I1 (g28721), .I2 (g23914));
AN2X1 gate11715(.O (g34371), .I1 (g7450), .I2 (g34044));
AN2X1 gate11716(.O (g24709), .I1 (g16690), .I2 (g23000));
AN2X1 gate11717(.O (g31542), .I1 (g19050), .I2 (g29814));
AN2X1 gate11718(.O (g31021), .I1 (g26025), .I2 (g29814));
AN2X1 gate11719(.O (g29523), .I1 (g28930), .I2 (g22417));
AN2X1 gate11720(.O (g23151), .I1 (g18994), .I2 (g7162));
AN2X1 gate11721(.O (g28111), .I1 (g27343), .I2 (g22716));
AN2X1 gate11722(.O (g14296), .I1 (g2638), .I2 (g11897));
AN2X1 gate11723(.O (g21996), .I1 (g5615), .I2 (g19074));
AN2X1 gate11724(.O (g24225), .I1 (g246), .I2 (g22594));
AN2X1 gate11725(.O (g15673), .I1 (g182), .I2 (g13437));
AN2X1 gate11726(.O (g18792), .I1 (g7051), .I2 (g15634));
AN2X1 gate11727(.O (g15847), .I1 (g3191), .I2 (g14005));
AN2X1 gate11728(.O (g23996), .I1 (g19596), .I2 (g10951));
AN2X1 gate11729(.O (g24708), .I1 (g16474), .I2 (g22998));
AN2X1 gate11730(.O (g14644), .I1 (g10610), .I2 (g10605));
AN3X1 gate11731(.O (g33913), .I1 (g23088), .I2 (g33204), .I3 (g9104));
AN2X1 gate11732(.O (g16592), .I1 (g5579), .I2 (g14688));
AN2X1 gate11733(.O (g21844), .I1 (g3873), .I2 (g21070));
AN2X1 gate11734(.O (g21394), .I1 (g13335), .I2 (g15799));
AN2X1 gate11735(.O (g32356), .I1 (g2704), .I2 (g31710));
AN2X1 gate11736(.O (g29475), .I1 (g14033), .I2 (g28500));
AN2X1 gate11737(.O (g18459), .I1 (g2331), .I2 (g15224));
AN2X1 gate11738(.O (g18425), .I1 (g2161), .I2 (g18008));
AN2X1 gate11739(.O (g33905), .I1 (g33089), .I2 (g15574));
AN2X1 gate11740(.O (g33073), .I1 (g32386), .I2 (g18828));
AN2X1 gate11741(.O (g12687), .I1 (g9024), .I2 (g8977));
AN2X1 gate11742(.O (g25106), .I1 (g17391), .I2 (g23506));
AN2X1 gate11743(.O (g26541), .I1 (g319), .I2 (g24375));
AN2X1 gate11744(.O (g34514), .I1 (g34286), .I2 (g19480));
AN2X1 gate11745(.O (g15851), .I1 (g3953), .I2 (g14157));
AN2X1 gate11746(.O (g15872), .I1 (g9095), .I2 (g14234));
AN2X1 gate11747(.O (g18458), .I1 (g2357), .I2 (g15224));
AN2X1 gate11748(.O (g19139), .I1 (g452), .I2 (g16195));
AN2X1 gate11749(.O (g27374), .I1 (g26519), .I2 (g17478));
AN3X1 gate11750(.O (g33530), .I1 (g32960), .I2 (I31346), .I3 (I31347));
AN2X1 gate11751(.O (g21420), .I1 (g16093), .I2 (g13596));
AN2X1 gate11752(.O (g34507), .I1 (g34280), .I2 (g19454));
AN2X1 gate11753(.O (g31122), .I1 (g12144), .I2 (g29993));
AN2X1 gate11754(.O (g32182), .I1 (g31753), .I2 (g27937));
AN4X1 gate11755(.O (g20069), .I1 (g16312), .I2 (g9051), .I3 (g9011), .I4 (g8955));
AN2X1 gate11756(.O (g33122), .I1 (g8859), .I2 (g32192));
AN2X1 gate11757(.O (g8530), .I1 (g2902), .I2 (g2907));
AN4X1 gate11758(.O (I31027), .I1 (g32494), .I2 (g32495), .I3 (g32496), .I4 (g32497));
AN3X1 gate11759(.O (I24524), .I1 (g5041), .I2 (g5046), .I3 (g9716));
AN3X1 gate11760(.O (g33464), .I1 (g32484), .I2 (I31016), .I3 (I31017));
AN3X1 gate11761(.O (I16129), .I1 (g8728), .I2 (g11443), .I3 (g11411));
AN2X1 gate11762(.O (g20602), .I1 (g10803), .I2 (g15580));
AN4X1 gate11763(.O (g28150), .I1 (g10862), .I2 (g11834), .I3 (g11283), .I4 (g27187));
AN3X1 gate11764(.O (g16846), .I1 (g14034), .I2 (g12591), .I3 (g11185));
AN2X1 gate11765(.O (g18545), .I1 (g2783), .I2 (g15277));
AN2X1 gate11766(.O (g25951), .I1 (g24500), .I2 (g19565));
AN2X1 gate11767(.O (g26325), .I1 (g12644), .I2 (g25370));
AN2X1 gate11768(.O (g24602), .I1 (g16507), .I2 (g22854));
AN2X1 gate11769(.O (g25972), .I1 (g2217), .I2 (g24993));
AN2X1 gate11770(.O (g18444), .I1 (g2269), .I2 (g18008));
AN2X1 gate11771(.O (g25033), .I1 (g17500), .I2 (g23433));
AN3X1 gate11772(.O (g25371), .I1 (g5062), .I2 (g22173), .I3 (I24524));
AN2X1 gate11773(.O (g20375), .I1 (g671), .I2 (g16846));
AN2X1 gate11774(.O (g24657), .I1 (g22644), .I2 (g19730));
AN2X1 gate11775(.O (g24774), .I1 (g718), .I2 (g23614));
AN2X1 gate11776(.O (g16731), .I1 (g7153), .I2 (g12941));
AN2X1 gate11777(.O (g26829), .I1 (g2844), .I2 (g24505));
AN2X1 gate11778(.O (g27669), .I1 (g26840), .I2 (g13278));
AN2X1 gate11779(.O (g17480), .I1 (g9683), .I2 (g14433));
AN2X1 gate11780(.O (g19333), .I1 (g464), .I2 (g16223));
AN2X1 gate11781(.O (g29347), .I1 (g29176), .I2 (g22201));
AN2X1 gate11782(.O (g18599), .I1 (g2955), .I2 (g16349));
AN2X1 gate11783(.O (g22307), .I1 (g20027), .I2 (g21163));
AN2X1 gate11784(.O (g22076), .I1 (g6255), .I2 (g19210));
AN2X1 gate11785(.O (g22085), .I1 (g6295), .I2 (g19210));
AN2X1 gate11786(.O (g26358), .I1 (g19522), .I2 (g25528));
AN3X1 gate11787(.O (I27349), .I1 (g25534), .I2 (g26424), .I3 (g22698));
AN2X1 gate11788(.O (g23025), .I1 (g16021), .I2 (g19798));
AN2X1 gate11789(.O (g27260), .I1 (g26766), .I2 (g26737));
AN2X1 gate11790(.O (g32331), .I1 (g31322), .I2 (g20637));
AN2X1 gate11791(.O (g31292), .I1 (g29735), .I2 (g23338));
AN2X1 gate11792(.O (g26828), .I1 (g24919), .I2 (g15756));
AN2X1 gate11793(.O (g27668), .I1 (g1367), .I2 (g25917));
AN2X1 gate11794(.O (g23540), .I1 (g16866), .I2 (g20622));
AN2X1 gate11795(.O (g18598), .I1 (g3003), .I2 (g16349));
AN2X1 gate11796(.O (g22054), .I1 (g6120), .I2 (g21611));
AN2X1 gate11797(.O (g28695), .I1 (g27580), .I2 (g20666));
AN2X1 gate11798(.O (g31153), .I1 (g12336), .I2 (g30068));
AN2X1 gate11799(.O (g27392), .I1 (g26576), .I2 (g17507));
AN2X1 gate11800(.O (g29600), .I1 (g1840), .I2 (g29049));
AN2X1 gate11801(.O (g26121), .I1 (g6167), .I2 (g25111));
AN2X1 gate11802(.O (g20171), .I1 (g16479), .I2 (g10476));
AN2X1 gate11803(.O (g34541), .I1 (g34331), .I2 (g20087));
AN2X1 gate11804(.O (g17307), .I1 (g9498), .I2 (g14343));
AN2X1 gate11805(.O (g15574), .I1 (g4311), .I2 (g13202));
AN2X1 gate11806(.O (g33409), .I1 (g32359), .I2 (g21408));
AN3X1 gate11807(.O (I24616), .I1 (g6082), .I2 (g6088), .I3 (g9946));
AN2X1 gate11808(.O (g29952), .I1 (g23576), .I2 (g28939));
AN2X1 gate11809(.O (g27559), .I1 (g26576), .I2 (g17777));
AN2X1 gate11810(.O (g29351), .I1 (g4771), .I2 (g28406));
AN2X1 gate11811(.O (g27525), .I1 (g26576), .I2 (g17720));
AN2X1 gate11812(.O (g27488), .I1 (g26549), .I2 (g17648));
AN2X1 gate11813(.O (g18817), .I1 (g6533), .I2 (g15483));
AN2X1 gate11814(.O (g15912), .I1 (g3562), .I2 (g14018));
AN4X1 gate11815(.O (g14581), .I1 (g12587), .I2 (g12428), .I3 (g12357), .I4 (I16695));
AN2X1 gate11816(.O (g18322), .I1 (g1608), .I2 (g17873));
AN2X1 gate11817(.O (g33408), .I1 (g32358), .I2 (g21407));
AN4X1 gate11818(.O (I31081), .I1 (g30673), .I2 (g31810), .I3 (g32571), .I4 (g32572));
AN2X1 gate11819(.O (g24967), .I1 (g23197), .I2 (g20213));
AN2X1 gate11820(.O (g10707), .I1 (g3787), .I2 (g8561));
AN2X1 gate11821(.O (g18159), .I1 (g671), .I2 (g17433));
AN2X1 gate11822(.O (g27558), .I1 (g26576), .I2 (g17776));
AN3X1 gate11823(.O (g25507), .I1 (g6098), .I2 (g23844), .I3 (I24616));
AN2X1 gate11824(.O (g22942), .I1 (g9104), .I2 (g20219));
AN2X1 gate11825(.O (g18125), .I1 (g15053), .I2 (g16886));
AN2X1 gate11826(.O (g18532), .I1 (g2724), .I2 (g15277));
AN2X1 gate11827(.O (g26291), .I1 (g2681), .I2 (g25439));
AN2X1 gate11828(.O (g30920), .I1 (g29889), .I2 (g21024));
AN4X1 gate11829(.O (I24704), .I1 (g21193), .I2 (g24061), .I3 (g24062), .I4 (g24063));
AN2X1 gate11830(.O (g19585), .I1 (g17180), .I2 (g14004));
AN2X1 gate11831(.O (g14202), .I1 (g869), .I2 (g10632));
AN2X1 gate11832(.O (g16929), .I1 (g6505), .I2 (g14348));
AN2X1 gate11833(.O (g18158), .I1 (g667), .I2 (g17433));
AN2X1 gate11834(.O (g14257), .I1 (g8612), .I2 (g11878));
AN2X1 gate11835(.O (g21957), .I1 (g5390), .I2 (g21514));
AN2X1 gate11836(.O (g18783), .I1 (g5841), .I2 (g18065));
AN2X1 gate11837(.O (g23957), .I1 (g4138), .I2 (g19589));
AN2X1 gate11838(.O (g29516), .I1 (g28895), .I2 (g22369));
AN4X1 gate11839(.O (g14496), .I1 (g12411), .I2 (g12244), .I3 (g12197), .I4 (I16618));
AN2X1 gate11840(.O (g22670), .I1 (g20114), .I2 (g9104));
AN2X1 gate11841(.O (g21739), .I1 (g3080), .I2 (g20330));
AN4X1 gate11842(.O (I31356), .I1 (g31327), .I2 (g31859), .I3 (g32968), .I4 (g32969));
AN2X1 gate11843(.O (g25163), .I1 (g20217), .I2 (g23566));
AN2X1 gate11844(.O (g18561), .I1 (g2841), .I2 (g15277));
AN2X1 gate11845(.O (g18656), .I1 (g15120), .I2 (g17128));
AN2X1 gate11846(.O (g30121), .I1 (g28577), .I2 (g21052));
AN2X1 gate11847(.O (g25012), .I1 (g20644), .I2 (g23419));
AN2X1 gate11848(.O (g18353), .I1 (g1772), .I2 (g17955));
AN2X1 gate11849(.O (g18295), .I1 (g1489), .I2 (g16449));
AN2X1 gate11850(.O (g21738), .I1 (g3072), .I2 (g20330));
AN3X1 gate11851(.O (g10590), .I1 (g7246), .I2 (g7392), .I3 (I13937));
AN2X1 gate11852(.O (g17156), .I1 (g305), .I2 (g13385));
AN2X1 gate11853(.O (g17655), .I1 (g7897), .I2 (g13342));
AN2X1 gate11854(.O (g18680), .I1 (g15128), .I2 (g15885));
AN2X1 gate11855(.O (g18144), .I1 (g590), .I2 (g17533));
AN2X1 gate11856(.O (g18823), .I1 (g6727), .I2 (g15680));
AN2X1 gate11857(.O (g34344), .I1 (g34107), .I2 (g20038));
AN2X1 gate11858(.O (g21699), .I1 (g142), .I2 (g20283));
AN2X1 gate11859(.O (g28706), .I1 (g27584), .I2 (g20681));
AN2X1 gate11860(.O (g28597), .I1 (g27515), .I2 (g20508));
AN4X1 gate11861(.O (I31182), .I1 (g32719), .I2 (g32720), .I3 (g32721), .I4 (g32722));
AN2X1 gate11862(.O (g18336), .I1 (g1700), .I2 (g17873));
AN2X1 gate11863(.O (g24545), .I1 (g3333), .I2 (g23285));
AN3X1 gate11864(.O (g33474), .I1 (g32556), .I2 (I31066), .I3 (I31067));
AN2X1 gate11865(.O (g28256), .I1 (g11398), .I2 (g27984));
AN2X1 gate11866(.O (g15820), .I1 (g3578), .I2 (g13955));
AN2X1 gate11867(.O (g28689), .I1 (g27575), .I2 (g20651));
AN2X1 gate11868(.O (g32149), .I1 (g31658), .I2 (g29983));
AN2X1 gate11869(.O (g27042), .I1 (g25774), .I2 (g19343));
AN3X1 gate11870(.O (g33711), .I1 (g33176), .I2 (g10727), .I3 (g22332));
AN2X1 gate11871(.O (g30173), .I1 (g28118), .I2 (g13082));
AN2X1 gate11872(.O (g34291), .I1 (g34055), .I2 (g19366));
AN2X1 gate11873(.O (g31327), .I1 (g19200), .I2 (g29814));
AN2X1 gate11874(.O (g27255), .I1 (g25936), .I2 (g19689));
AN2X1 gate11875(.O (g28280), .I1 (g23761), .I2 (g27724));
AN2X1 gate11876(.O (g22131), .I1 (g6641), .I2 (g19277));
AN2X1 gate11877(.O (g29834), .I1 (g28368), .I2 (g23278));
AN2X1 gate11878(.O (g33327), .I1 (g32208), .I2 (g20561));
AN2X1 gate11879(.O (g34173), .I1 (g33679), .I2 (g24368));
AN3X1 gate11880(.O (I24064), .I1 (g3385), .I2 (g3391), .I3 (g8492));
AN3X1 gate11881(.O (g29208), .I1 (g24138), .I2 (I27538), .I3 (I27539));
AN2X1 gate11882(.O (g25788), .I1 (g8010), .I2 (g24579));
AN2X1 gate11883(.O (g32148), .I1 (g31631), .I2 (g29981));
AN2X1 gate11884(.O (g28624), .I1 (g22357), .I2 (g27009));
AN2X1 gate11885(.O (g28300), .I1 (g27771), .I2 (g26605));
AN2X1 gate11886(.O (g27270), .I1 (g26805), .I2 (g26793));
AN2X1 gate11887(.O (g32097), .I1 (g25960), .I2 (g31021));
AN4X1 gate11888(.O (I31331), .I1 (g30825), .I2 (g31854), .I3 (g32933), .I4 (g32934));
AN2X1 gate11889(.O (g27678), .I1 (g947), .I2 (g25830));
AN2X1 gate11890(.O (g18631), .I1 (g3694), .I2 (g17226));
AN2X1 gate11891(.O (g32104), .I1 (g31616), .I2 (g29906));
AN3X1 gate11892(.O (g7520), .I1 (g2704), .I2 (g2697), .I3 (g2689));
AN2X1 gate11893(.O (g18364), .I1 (g1844), .I2 (g17955));
AN2X1 gate11894(.O (g32343), .I1 (g31473), .I2 (g20710));
AN2X1 gate11895(.O (g31283), .I1 (g30156), .I2 (g27837));
AN2X1 gate11896(.O (g27460), .I1 (g26549), .I2 (g17610));
AN2X1 gate11897(.O (g27686), .I1 (g1291), .I2 (g25849));
AN2X1 gate11898(.O (g25946), .I1 (g24496), .I2 (g19537));
AN2X1 gate11899(.O (g31492), .I1 (g29790), .I2 (g23431));
AN2X1 gate11900(.O (g24817), .I1 (g22929), .I2 (g7235));
AN2X1 gate11901(.O (g30029), .I1 (g29164), .I2 (g12936));
AN3X1 gate11902(.O (g33492), .I1 (g32686), .I2 (I31156), .I3 (I31157));
AN2X1 gate11903(.O (g19674), .I1 (g2819), .I2 (g15867));
AN2X1 gate11904(.O (g24322), .I1 (g4423), .I2 (g22228));
AN2X1 gate11905(.O (g12939), .I1 (g405), .I2 (g11048));
AN2X1 gate11906(.O (g27030), .I1 (g26343), .I2 (g7947));
AN2X1 gate11907(.O (g20977), .I1 (g10123), .I2 (g17301));
AN2X1 gate11908(.O (g13299), .I1 (g437), .I2 (g11048));
AN2X1 gate11909(.O (g24532), .I1 (g22331), .I2 (g19478));
AN2X1 gate11910(.O (g32369), .I1 (g2130), .I2 (g31672));
AN2X1 gate11911(.O (g27267), .I1 (g26026), .I2 (g17124));
AN2X1 gate11912(.O (g27294), .I1 (g9975), .I2 (g26656));
AN2X1 gate11913(.O (g29614), .I1 (g28860), .I2 (g22369));
AN2X1 gate11914(.O (g30028), .I1 (g29069), .I2 (g9311));
AN3X1 gate11915(.O (g28231), .I1 (g27187), .I2 (g22763), .I3 (g27074));
AN2X1 gate11916(.O (g24977), .I1 (g23209), .I2 (g20232));
AN2X1 gate11917(.O (g34506), .I1 (g8833), .I2 (g34354));
AN2X1 gate11918(.O (g16803), .I1 (g5933), .I2 (g14810));
AN2X1 gate11919(.O (g31750), .I1 (g30103), .I2 (g23925));
AN2X1 gate11920(.O (g29607), .I1 (g28509), .I2 (g14208));
AN2X1 gate11921(.O (g18289), .I1 (g1448), .I2 (g16449));
AN4X1 gate11922(.O (I31026), .I1 (g31194), .I2 (g31800), .I3 (g32492), .I4 (g32493));
AN2X1 gate11923(.O (g29320), .I1 (g29068), .I2 (g22147));
AN2X1 gate11924(.O (g33381), .I1 (g11842), .I2 (g32318));
AN4X1 gate11925(.O (I31212), .I1 (g32761), .I2 (g32762), .I3 (g32763), .I4 (g32764));
AN4X1 gate11926(.O (g29073), .I1 (g27163), .I2 (g10290), .I3 (g21012), .I4 (I27409));
AN2X1 gate11927(.O (g12065), .I1 (g9557), .I2 (g9805));
AN2X1 gate11928(.O (g18309), .I1 (g1339), .I2 (g16931));
AN2X1 gate11929(.O (g29530), .I1 (g1612), .I2 (g28820));
AN2X1 gate11930(.O (g24656), .I1 (g11736), .I2 (g22926));
AN2X1 gate11931(.O (g29593), .I1 (g28470), .I2 (g7985));
AN2X1 gate11932(.O (g33091), .I1 (g32392), .I2 (g18897));
AN2X1 gate11933(.O (g18288), .I1 (g1454), .I2 (g16449));
AN2X1 gate11934(.O (g18224), .I1 (g1036), .I2 (g16100));
AN2X1 gate11935(.O (g21715), .I1 (g160), .I2 (g20283));
AN2X1 gate11936(.O (g22039), .I1 (g5949), .I2 (g19147));
AN2X1 gate11937(.O (g29346), .I1 (g4894), .I2 (g28381));
AN2X1 gate11938(.O (g25173), .I1 (g12234), .I2 (g23589));
AN2X1 gate11939(.O (g24295), .I1 (g4434), .I2 (g22550));
AN2X1 gate11940(.O (g18571), .I1 (g2856), .I2 (g16349));
AN2X1 gate11941(.O (g18308), .I1 (g6832), .I2 (g16931));
AN2X1 gate11942(.O (g24680), .I1 (g16422), .I2 (g22986));
AN2X1 gate11943(.O (g27219), .I1 (g26026), .I2 (g16742));
AN2X1 gate11944(.O (g32412), .I1 (g4765), .I2 (g30998));
AN2X1 gate11945(.O (g24144), .I1 (g17727), .I2 (g21660));
AN2X1 gate11946(.O (g33796), .I1 (g33117), .I2 (g25267));
AN2X1 gate11947(.O (g19692), .I1 (g12066), .I2 (g17086));
AN3X1 gate11948(.O (I24555), .I1 (g9559), .I2 (g9809), .I3 (g6093));
AN2X1 gate11949(.O (g29565), .I1 (g1932), .I2 (g28590));
AN2X1 gate11950(.O (g26604), .I1 (g13248), .I2 (g25051));
AN2X1 gate11951(.O (g17469), .I1 (g4076), .I2 (g13217));
AN2X1 gate11952(.O (g13737), .I1 (g4501), .I2 (g10571));
AN2X1 gate11953(.O (g22038), .I1 (g5945), .I2 (g19147));
AN2X1 gate11954(.O (g23551), .I1 (g10793), .I2 (g18948));
AN2X1 gate11955(.O (g23572), .I1 (g20230), .I2 (g20656));
AN2X1 gate11956(.O (g10917), .I1 (g9174), .I2 (g1087));
AN2X1 gate11957(.O (g12219), .I1 (g1189), .I2 (g7532));
AN2X1 gate11958(.O (g27218), .I1 (g25997), .I2 (g16740));
AN2X1 gate11959(.O (g30927), .I1 (g29910), .I2 (g24795));
AN2X1 gate11960(.O (g18495), .I1 (g2533), .I2 (g15426));
AN2X1 gate11961(.O (g33840), .I1 (g33253), .I2 (g20267));
AN2X1 gate11962(.O (g29641), .I1 (g28520), .I2 (g14237));
AN2X1 gate11963(.O (g29797), .I1 (g28347), .I2 (g23259));
AN2X1 gate11964(.O (g16662), .I1 (g4552), .I2 (g14753));
AN2X1 gate11965(.O (g13697), .I1 (g11166), .I2 (g8608));
AN2X1 gate11966(.O (g28660), .I1 (g27824), .I2 (g20623));
AN2X1 gate11967(.O (g18816), .I1 (g6527), .I2 (g15483));
AN2X1 gate11968(.O (g32011), .I1 (g8287), .I2 (g31134));
AN2X1 gate11969(.O (g27160), .I1 (g14163), .I2 (g26340));
AN2X1 gate11970(.O (g10706), .I1 (g3338), .I2 (g8691));
AN2X1 gate11971(.O (g15113), .I1 (g4291), .I2 (g14454));
AN2X1 gate11972(.O (g19207), .I1 (g7803), .I2 (g15992));
AN2X1 gate11973(.O (g18687), .I1 (g4664), .I2 (g15885));
AN2X1 gate11974(.O (g28456), .I1 (g27290), .I2 (g20104));
AN4X1 gate11975(.O (I31097), .I1 (g32596), .I2 (g32597), .I3 (g32598), .I4 (g32599));
AN2X1 gate11976(.O (g17601), .I1 (g9616), .I2 (g14572));
AN2X1 gate11977(.O (g22143), .I1 (g19568), .I2 (g10971));
AN2X1 gate11978(.O (g21784), .I1 (g3423), .I2 (g20391));
AN2X1 gate11979(.O (g22937), .I1 (g753), .I2 (g20540));
AN2X1 gate11980(.O (g26845), .I1 (g24391), .I2 (g21426));
AN2X1 gate11981(.O (g14256), .I1 (g2079), .I2 (g11872));
AN2X1 gate11982(.O (g21956), .I1 (g5360), .I2 (g21514));
AN2X1 gate11983(.O (g18752), .I1 (g15146), .I2 (g17926));
AN2X1 gate11984(.O (g27455), .I1 (g26488), .I2 (g17603));
AN2X1 gate11985(.O (g26395), .I1 (g22547), .I2 (g25561));
AN2X1 gate11986(.O (g30604), .I1 (g18911), .I2 (g29878));
AN3X1 gate11987(.O (g33522), .I1 (g32902), .I2 (I31306), .I3 (I31307));
AN2X1 gate11988(.O (g18374), .I1 (g1878), .I2 (g15171));
AN2X1 gate11989(.O (g29635), .I1 (g28910), .I2 (g22432));
AN2X1 gate11990(.O (g21889), .I1 (g4169), .I2 (g19801));
AN2X1 gate11991(.O (g23103), .I1 (g10143), .I2 (g20765));
AN4X1 gate11992(.O (g27617), .I1 (g23032), .I2 (g26264), .I3 (g26424), .I4 (g24982));
AN2X1 gate11993(.O (g15105), .I1 (g4235), .I2 (g14454));
AN2X1 gate11994(.O (g21980), .I1 (g5567), .I2 (g19074));
AN2X1 gate11995(.O (g10624), .I1 (g8387), .I2 (g3072));
AN2X1 gate11996(.O (g28550), .I1 (g12009), .I2 (g27092));
AN2X1 gate11997(.O (g18643), .I1 (g3849), .I2 (g17096));
AN2X1 gate11998(.O (g7469), .I1 (g4382), .I2 (g4438));
AN2X1 gate11999(.O (g32310), .I1 (g27577), .I2 (g31376));
AN2X1 gate12000(.O (g16204), .I1 (g6537), .I2 (g14348));
AN2X1 gate12001(.O (g28314), .I1 (g27552), .I2 (g14205));
AN2X1 gate12002(.O (g21888), .I1 (g4165), .I2 (g19801));
AN2X1 gate12003(.O (g21824), .I1 (g3706), .I2 (g20453));
AN2X1 gate12004(.O (g26633), .I1 (g24964), .I2 (g20616));
AN2X1 gate12005(.O (g34563), .I1 (g34372), .I2 (g17465));
AN3X1 gate12006(.O (I17542), .I1 (g13156), .I2 (g6767), .I3 (g6756));
AN2X1 gate12007(.O (g27201), .I1 (g25997), .I2 (g16685));
AN2X1 gate12008(.O (g27277), .I1 (g26359), .I2 (g14191));
AN4X1 gate12009(.O (I24675), .I1 (g24022), .I2 (g24023), .I3 (g24024), .I4 (g24025));
AN3X1 gate12010(.O (g33483), .I1 (g32621), .I2 (I31111), .I3 (I31112));
AN2X1 gate12011(.O (g26719), .I1 (g10709), .I2 (g24438));
AN2X1 gate12012(.O (g24289), .I1 (g4427), .I2 (g22550));
AN2X1 gate12013(.O (g18669), .I1 (g4608), .I2 (g17367));
AN2X1 gate12014(.O (g32112), .I1 (g31646), .I2 (g29923));
AN2X1 gate12015(.O (g25927), .I1 (g25004), .I2 (g20375));
AN2X1 gate12016(.O (g32050), .I1 (g11003), .I2 (g30825));
AN2X1 gate12017(.O (g24309), .I1 (g4480), .I2 (g22228));
AN2X1 gate12018(.O (g33862), .I1 (g33272), .I2 (g20504));
AN2X1 gate12019(.O (g18260), .I1 (g1252), .I2 (g16000));
AN2X1 gate12020(.O (g28243), .I1 (g27879), .I2 (g23423));
AN2X1 gate12021(.O (g24288), .I1 (g4417), .I2 (g22550));
AN2X1 gate12022(.O (g27595), .I1 (g26733), .I2 (g26703));
AN2X1 gate12023(.O (g24224), .I1 (g269), .I2 (g22594));
AN2X1 gate12024(.O (g18668), .I1 (g4322), .I2 (g17367));
AN2X1 gate12025(.O (g27467), .I1 (g269), .I2 (g26832));
AN4X1 gate12026(.O (g27494), .I1 (g8038), .I2 (g26314), .I3 (g518), .I4 (g9077));
AN2X1 gate12027(.O (g31949), .I1 (g1287), .I2 (g30825));
AN2X1 gate12028(.O (g18392), .I1 (g1988), .I2 (g15171));
AN2X1 gate12029(.O (g29891), .I1 (g28420), .I2 (g23356));
AN2X1 gate12030(.O (g24308), .I1 (g4489), .I2 (g22228));
AN2X1 gate12031(.O (g21931), .I1 (g5188), .I2 (g18997));
AN2X1 gate12032(.O (g18195), .I1 (g847), .I2 (g17821));
AN2X1 gate12033(.O (g22015), .I1 (g5719), .I2 (g21562));
AN2X1 gate12034(.O (g18489), .I1 (g2509), .I2 (g15426));
AN2X1 gate12035(.O (g34395), .I1 (g34193), .I2 (g21336));
AN2X1 gate12036(.O (g31948), .I1 (g30670), .I2 (g18884));
AN2X1 gate12037(.O (g32096), .I1 (g31601), .I2 (g29893));
AN2X1 gate12038(.O (g28269), .I1 (g27205), .I2 (g19712));
AN2X1 gate12039(.O (g29575), .I1 (g2066), .I2 (g28604));
AN2X1 gate12040(.O (g15881), .I1 (g3582), .I2 (g13983));
AN2X1 gate12041(.O (g18559), .I1 (g12856), .I2 (g15277));
AN2X1 gate12042(.O (g25491), .I1 (g23615), .I2 (g21355));
AN2X1 gate12043(.O (g18525), .I1 (g2610), .I2 (g15509));
AN2X1 gate12044(.O (g18488), .I1 (g2495), .I2 (g15426));
AN2X1 gate12045(.O (g18424), .I1 (g2165), .I2 (g18008));
AN2X1 gate12046(.O (g28341), .I1 (g27240), .I2 (g19790));
AN2X1 gate12047(.O (g29711), .I1 (g2541), .I2 (g29134));
AN2X1 gate12048(.O (g33904), .I1 (g33321), .I2 (g21059));
AN2X1 gate12049(.O (g24495), .I1 (g6928), .I2 (g23127));
AN2X1 gate12050(.O (g28268), .I1 (g8572), .I2 (g27990));
AN2X1 gate12051(.O (g31252), .I1 (g29643), .I2 (g20101));
AN2X1 gate12052(.O (g29327), .I1 (g29070), .I2 (g22156));
AN2X1 gate12053(.O (g26861), .I1 (g25021), .I2 (g25003));
AN2X1 gate12054(.O (g33252), .I1 (g32155), .I2 (g20064));
AN2X1 gate12055(.O (g13080), .I1 (g6923), .I2 (g11357));
AN2X1 gate12056(.O (g18558), .I1 (g2803), .I2 (g15277));
AN2X1 gate12057(.O (g28655), .I1 (g27561), .I2 (g20603));
AN2X1 gate12058(.O (g30191), .I1 (g28647), .I2 (g23843));
AN2X1 gate12059(.O (g16233), .I1 (g6137), .I2 (g14251));
AN2X1 gate12060(.O (g29537), .I1 (g28976), .I2 (g22472));
AN2X1 gate12061(.O (g34191), .I1 (g33713), .I2 (g24404));
AN2X1 gate12062(.O (g16672), .I1 (g6295), .I2 (g15008));
AN2X1 gate12063(.O (g27822), .I1 (g4157), .I2 (g25893));
AN4X1 gate12064(.O (I27539), .I1 (g28040), .I2 (g24135), .I3 (g24136), .I4 (g24137));
AN2X1 gate12065(.O (g26389), .I1 (g19949), .I2 (g25553));
AN2X1 gate12066(.O (g18893), .I1 (g16215), .I2 (g16030));
AN2X1 gate12067(.O (g25981), .I1 (g2051), .I2 (g25007));
AN2X1 gate12068(.O (g24687), .I1 (g5827), .I2 (g23666));
AN4X1 gate12069(.O (I31011), .I1 (g30735), .I2 (g31797), .I3 (g32471), .I4 (g32472));
AN2X1 gate12070(.O (g27266), .I1 (g26789), .I2 (g26770));
AN2X1 gate12071(.O (g26612), .I1 (g901), .I2 (g24407));
AN4X1 gate12072(.O (I27538), .I1 (g21209), .I2 (g24132), .I3 (g24133), .I4 (g24134));
AN2X1 gate12073(.O (g26388), .I1 (g19595), .I2 (g25552));
AN2X1 gate12074(.O (g18544), .I1 (g2791), .I2 (g15277));
AN2X1 gate12075(.O (g26324), .I1 (g2661), .I2 (g25439));
AN2X1 gate12076(.O (g32428), .I1 (g31133), .I2 (g16261));
AN2X1 gate12077(.O (g29606), .I1 (g28480), .I2 (g8011));
AN2X1 gate12078(.O (g21024), .I1 (g16306), .I2 (g4871));
AN2X1 gate12079(.O (g18713), .I1 (g4836), .I2 (g15915));
AN2X1 gate12080(.O (g13461), .I1 (g2719), .I2 (g11819));
AN2X1 gate12081(.O (g22084), .I1 (g6291), .I2 (g19210));
AN2X1 gate12082(.O (g31183), .I1 (g30249), .I2 (g25174));
AN2X1 gate12083(.O (g26251), .I1 (g1988), .I2 (g25341));
AN2X1 gate12084(.O (g22110), .I1 (g15167), .I2 (g19277));
AN2X1 gate12085(.O (g24643), .I1 (g22636), .I2 (g19696));
AN2X1 gate12086(.O (g26272), .I1 (g2036), .I2 (g25470));
AN2X1 gate12087(.O (g33847), .I1 (g33260), .I2 (g20383));
AN2X1 gate12088(.O (g21860), .I1 (g3945), .I2 (g21070));
AN2X1 gate12089(.O (g16513), .I1 (g8345), .I2 (g13708));
AN2X1 gate12090(.O (g28694), .I1 (g27579), .I2 (g20664));
AN2X1 gate12091(.O (g29750), .I1 (g28296), .I2 (g23215));
AN2X1 gate12092(.O (g29982), .I1 (g23656), .I2 (g28998));
AN2X1 gate12093(.O (g29381), .I1 (g28135), .I2 (g19399));
AN2X1 gate12094(.O (g18610), .I1 (g15088), .I2 (g17059));
AN2X1 gate12095(.O (g34861), .I1 (g16540), .I2 (g34827));
AN2X1 gate12096(.O (g30247), .I1 (g28735), .I2 (g23937));
AN2X1 gate12097(.O (g18705), .I1 (g4801), .I2 (g16782));
AN2X1 gate12098(.O (g13887), .I1 (g5204), .I2 (g12402));
AN2X1 gate12099(.O (g25990), .I1 (g9461), .I2 (g25017));
AN2X1 gate12100(.O (g23497), .I1 (g20169), .I2 (g20569));
AN3X1 gate12101(.O (g33509), .I1 (g32809), .I2 (I31241), .I3 (I31242));
AN2X1 gate12102(.O (g24669), .I1 (g22653), .I2 (g19742));
AN2X1 gate12103(.O (g31933), .I1 (g939), .I2 (g30735));
AN2X1 gate12104(.O (g30926), .I1 (g29903), .I2 (g21163));
AN2X1 gate12105(.O (g30045), .I1 (g29200), .I2 (g12419));
AN2X1 gate12106(.O (g18255), .I1 (g1087), .I2 (g16897));
AN2X1 gate12107(.O (g18189), .I1 (g812), .I2 (g17821));
AN2X1 gate12108(.O (g27588), .I1 (g26690), .I2 (g26673));
AN2X1 gate12109(.O (g15779), .I1 (g13909), .I2 (g11214));
AN2X1 gate12110(.O (g18679), .I1 (g4633), .I2 (g15758));
AN2X1 gate12111(.O (g31508), .I1 (g29813), .I2 (g23459));
AN2X1 gate12112(.O (g34389), .I1 (g34170), .I2 (g20715));
AN2X1 gate12113(.O (g17321), .I1 (g1418), .I2 (g13105));
AN4X1 gate12114(.O (I31112), .I1 (g32617), .I2 (g32618), .I3 (g32619), .I4 (g32620));
AN2X1 gate12115(.O (g34045), .I1 (g33766), .I2 (g22942));
AN2X1 gate12116(.O (g30612), .I1 (g26338), .I2 (g29597));
AN3X1 gate12117(.O (g33508), .I1 (g32802), .I2 (I31236), .I3 (I31237));
AN2X1 gate12118(.O (g24668), .I1 (g11754), .I2 (g22979));
AN2X1 gate12119(.O (g21700), .I1 (g150), .I2 (g20283));
AN2X1 gate12120(.O (g30099), .I1 (g28549), .I2 (g20776));
AN2X1 gate12121(.O (g33872), .I1 (g33282), .I2 (g20548));
AN2X1 gate12122(.O (g18270), .I1 (g1291), .I2 (g16031));
AN2X1 gate12123(.O (g29796), .I1 (g28345), .I2 (g23258));
AN2X1 gate12124(.O (g17179), .I1 (g1041), .I2 (g13211));
AN2X1 gate12125(.O (g24392), .I1 (g3115), .I2 (g23067));
AN2X1 gate12126(.O (g22685), .I1 (g11891), .I2 (g20192));
AN2X1 gate12127(.O (g18188), .I1 (g807), .I2 (g17328));
AN2X1 gate12128(.O (g18124), .I1 (g102), .I2 (g16886));
AN2X1 gate12129(.O (g21987), .I1 (g5579), .I2 (g19074));
AN2X1 gate12130(.O (g18678), .I1 (g66), .I2 (g15758));
AN2X1 gate12131(.O (g34388), .I1 (g10802), .I2 (g34062));
AN2X1 gate12132(.O (g16026), .I1 (g854), .I2 (g14065));
AN2X1 gate12133(.O (g28557), .I1 (g27772), .I2 (g15647));
AN2X1 gate12134(.O (g34324), .I1 (g14064), .I2 (g34161));
AN2X1 gate12135(.O (g15081), .I1 (g2689), .I2 (g12983));
AN2X1 gate12136(.O (g13393), .I1 (g703), .I2 (g11048));
AN2X1 gate12137(.O (g16212), .I1 (g6167), .I2 (g14321));
AN2X1 gate12138(.O (g24195), .I1 (g74), .I2 (g22722));
AN2X1 gate12139(.O (g28210), .I1 (g9229), .I2 (g27554));
AN2X1 gate12140(.O (g32317), .I1 (g5507), .I2 (g31542));
AN2X1 gate12141(.O (g27119), .I1 (g25877), .I2 (g22542));
AN2X1 gate12142(.O (g30098), .I1 (g28548), .I2 (g20774));
AN2X1 gate12143(.O (g34701), .I1 (g34536), .I2 (g20179));
AN4X1 gate12144(.O (g10721), .I1 (g3288), .I2 (g6875), .I3 (g3274), .I4 (g8481));
AN2X1 gate12145(.O (g20559), .I1 (g336), .I2 (g15831));
AN2X1 gate12146(.O (g30251), .I1 (g28745), .I2 (g23940));
AN2X1 gate12147(.O (g34534), .I1 (g34321), .I2 (g19743));
AN2X1 gate12148(.O (g23658), .I1 (g14687), .I2 (g20852));
AN2X1 gate12149(.O (g30272), .I1 (g28814), .I2 (g23982));
AN3X1 gate12150(.O (g34098), .I1 (g33744), .I2 (g9104), .I3 (g18957));
AN2X1 gate12151(.O (g19206), .I1 (g460), .I2 (g16206));
AN2X1 gate12152(.O (g15786), .I1 (g13940), .I2 (g11233));
AN2X1 gate12153(.O (g18460), .I1 (g2351), .I2 (g15224));
AN2X1 gate12154(.O (g18686), .I1 (g4659), .I2 (g15885));
AN2X1 gate12155(.O (g24559), .I1 (g22993), .I2 (g19567));
AN2X1 gate12156(.O (g18383), .I1 (g1950), .I2 (g15171));
AN2X1 gate12157(.O (g29840), .I1 (g2153), .I2 (g29056));
AN2X1 gate12158(.O (g24488), .I1 (g6905), .I2 (g23082));
AN4X1 gate12159(.O (I31096), .I1 (g31376), .I2 (g31812), .I3 (g32594), .I4 (g32595));
AN2X1 gate12160(.O (g24016), .I1 (g14528), .I2 (g21610));
AN2X1 gate12161(.O (g27118), .I1 (g26055), .I2 (g16529));
AN3X1 gate12162(.O (g22417), .I1 (g7753), .I2 (g9285), .I3 (g21186));
AN2X1 gate12163(.O (g11960), .I1 (g2495), .I2 (g7424));
AN2X1 gate12164(.O (g32129), .I1 (g31658), .I2 (g29955));
AN2X1 gate12165(.O (g21943), .I1 (g5240), .I2 (g18997));
AN2X1 gate12166(.O (g25832), .I1 (g8219), .I2 (g24625));
AN2X1 gate12167(.O (g21296), .I1 (g7879), .I2 (g16072));
AN2X1 gate12168(.O (g24558), .I1 (g22516), .I2 (g19566));
AN2X1 gate12169(.O (g18267), .I1 (g1266), .I2 (g16000));
AN2X1 gate12170(.O (g18294), .I1 (g15072), .I2 (g16449));
AN2X1 gate12171(.O (g27616), .I1 (g26349), .I2 (g20449));
AN2X1 gate12172(.O (g26871), .I1 (g25038), .I2 (g25020));
AN2X1 gate12173(.O (g17654), .I1 (g962), .I2 (g13284));
AN2X1 gate12174(.O (g32128), .I1 (g31631), .I2 (g29953));
AN3X1 gate12175(.O (I17575), .I1 (g13156), .I2 (g11450), .I3 (g6756));
AN2X1 gate12176(.O (g27313), .I1 (g1982), .I2 (g26701));
AN2X1 gate12177(.O (g29192), .I1 (g27163), .I2 (g10290));
AN2X1 gate12178(.O (g30032), .I1 (g29072), .I2 (g9326));
AN2X1 gate12179(.O (g21969), .I1 (g5373), .I2 (g21514));
AN2X1 gate12180(.O (g26360), .I1 (g10589), .I2 (g25533));
AN2X1 gate12181(.O (g25573), .I1 (I24704), .I2 (I24705));
AN2X1 gate12182(.O (g30140), .I1 (g28600), .I2 (g23749));
AN2X1 gate12183(.O (g27276), .I1 (g9750), .I2 (g26607));
AN2X1 gate12184(.O (g27285), .I1 (g9912), .I2 (g26632));
AN2X1 gate12185(.O (g29522), .I1 (g28923), .I2 (g22369));
AN2X1 gate12186(.O (g32323), .I1 (g31311), .I2 (g20610));
AN2X1 gate12187(.O (g24865), .I1 (g11323), .I2 (g23253));
AN2X1 gate12188(.O (g29663), .I1 (g1950), .I2 (g28693));
AN2X1 gate12189(.O (g34140), .I1 (g33931), .I2 (g23802));
AN2X1 gate12190(.O (g22762), .I1 (g9305), .I2 (g20645));
AN2X1 gate12191(.O (g15651), .I1 (g429), .I2 (g13414));
AN2X1 gate12192(.O (g21968), .I1 (g5459), .I2 (g21514));
AN2X1 gate12193(.O (g10655), .I1 (g8440), .I2 (g3423));
AN2X1 gate12194(.O (g15672), .I1 (g433), .I2 (g13458));
AN2X1 gate12195(.O (g27305), .I1 (g10041), .I2 (g26683));
AN2X1 gate12196(.O (g25926), .I1 (g25005), .I2 (g24839));
AN2X1 gate12197(.O (g24713), .I1 (g5831), .I2 (g23666));
AN2X1 gate12198(.O (g25045), .I1 (g17525), .I2 (g23448));
AN2X1 gate12199(.O (g18219), .I1 (g969), .I2 (g16100));
AN2X1 gate12200(.O (g27254), .I1 (g25935), .I2 (g19688));
AN2X1 gate12201(.O (g30061), .I1 (g1036), .I2 (g28188));
AN2X1 gate12202(.O (g33311), .I1 (g31942), .I2 (g12925));
AN2X1 gate12203(.O (g21855), .I1 (g3925), .I2 (g21070));
AN2X1 gate12204(.O (g34061), .I1 (g33800), .I2 (g23076));
AN2X1 gate12205(.O (g14180), .I1 (g872), .I2 (g10632));
AN2X1 gate12206(.O (g23855), .I1 (g4112), .I2 (g19455));
AN2X1 gate12207(.O (g22216), .I1 (g13660), .I2 (g20000));
AN2X1 gate12208(.O (g18218), .I1 (g1008), .I2 (g16100));
AN2X1 gate12209(.O (g21870), .I1 (g4093), .I2 (g19801));
AN3X1 gate12210(.O (I17606), .I1 (g14988), .I2 (g11450), .I3 (g6756));
AN2X1 gate12211(.O (g28601), .I1 (g27506), .I2 (g20514));
AN2X1 gate12212(.O (g28677), .I1 (g27571), .I2 (g20635));
AN2X1 gate12213(.O (g27036), .I1 (g26329), .I2 (g11038));
AN2X1 gate12214(.O (g29553), .I1 (g2437), .I2 (g28911));
AN2X1 gate12215(.O (g26629), .I1 (g14173), .I2 (g24418));
AN2X1 gate12216(.O (g27177), .I1 (g25997), .I2 (g16651));
AN2X1 gate12217(.O (g27560), .I1 (g26299), .I2 (g20191));
AN2X1 gate12218(.O (g34871), .I1 (g34823), .I2 (g19908));
AN2X1 gate12219(.O (g24189), .I1 (g324), .I2 (g22722));
AN2X1 gate12220(.O (g31756), .I1 (g30114), .I2 (g23942));
AN2X1 gate12221(.O (g24679), .I1 (g13289), .I2 (g22985));
AN2X1 gate12222(.O (g11244), .I1 (g8346), .I2 (g8566));
AN2X1 gate12223(.O (g29949), .I1 (g23575), .I2 (g28924));
AN2X1 gate12224(.O (g32232), .I1 (g31241), .I2 (g20266));
AN2X1 gate12225(.O (g20188), .I1 (g5849), .I2 (g17772));
AN2X1 gate12226(.O (g18160), .I1 (g645), .I2 (g17433));
AN2X1 gate12227(.O (g29326), .I1 (g29105), .I2 (g22155));
AN3X1 gate12228(.O (g10838), .I1 (g7738), .I2 (g5527), .I3 (g5535));
AN2X1 gate12229(.O (g28143), .I1 (g27344), .I2 (g26083));
AN2X1 gate12230(.O (g31780), .I1 (g30163), .I2 (g23999));
AN3X1 gate12231(.O (g25462), .I1 (g6404), .I2 (g22300), .I3 (I24585));
AN2X1 gate12232(.O (g24188), .I1 (g316), .I2 (g22722));
AN2X1 gate12233(.O (g22117), .I1 (g6597), .I2 (g19277));
AN2X1 gate12234(.O (g29536), .I1 (g28969), .I2 (g22432));
AN2X1 gate12235(.O (g22000), .I1 (g5727), .I2 (g21562));
AN2X1 gate12236(.O (g21867), .I1 (g4082), .I2 (g19801));
AN2X1 gate12237(.O (g18455), .I1 (g2327), .I2 (g15224));
AN2X1 gate12238(.O (g24686), .I1 (g5485), .I2 (g23630));
AN2X1 gate12239(.O (g24939), .I1 (g23771), .I2 (g21012));
AN2X1 gate12240(.O (g29757), .I1 (g28305), .I2 (g23221));
AN4X1 gate12241(.O (I31317), .I1 (g32914), .I2 (g32915), .I3 (g32916), .I4 (g32917));
AN2X1 gate12242(.O (g33350), .I1 (g32235), .I2 (g20702));
AN2X1 gate12243(.O (g32261), .I1 (g31251), .I2 (g20386));
AN2X1 gate12244(.O (g18617), .I1 (g3462), .I2 (g17062));
AN2X1 gate12245(.O (g18470), .I1 (g2403), .I2 (g15224));
AN2X1 gate12246(.O (g20093), .I1 (g15372), .I2 (g14584));
AN2X1 gate12247(.O (g33820), .I1 (g33075), .I2 (g26830));
AN2X1 gate12248(.O (g29621), .I1 (g2449), .I2 (g28994));
AN3X1 gate12249(.O (I24576), .I1 (g5390), .I2 (g5396), .I3 (g9792));
AN3X1 gate12250(.O (I24585), .I1 (g9621), .I2 (g9892), .I3 (g6439));
AN2X1 gate12251(.O (g10619), .I1 (g3080), .I2 (g7907));
AN2X1 gate12252(.O (g21714), .I1 (g278), .I2 (g20283));
AN2X1 gate12253(.O (g23581), .I1 (g20183), .I2 (g11900));
AN2X1 gate12254(.O (g24294), .I1 (g4452), .I2 (g22550));
AN2X1 gate12255(.O (g31152), .I1 (g10039), .I2 (g30067));
AN2X1 gate12256(.O (g25061), .I1 (g17586), .I2 (g23461));
AN4X1 gate12257(.O (I31002), .I1 (g32459), .I2 (g32460), .I3 (g32461), .I4 (g32462));
AN2X1 gate12258(.O (g18201), .I1 (g15061), .I2 (g15938));
AN2X1 gate12259(.O (g33846), .I1 (g33259), .I2 (g20380));
AN4X1 gate12260(.O (I31057), .I1 (g32538), .I2 (g32539), .I3 (g32540), .I4 (g32541));
AN2X1 gate12261(.O (g21707), .I1 (g191), .I2 (g20283));
AN2X1 gate12262(.O (g21819), .I1 (g3614), .I2 (g20924));
AN2X1 gate12263(.O (g29564), .I1 (g1882), .I2 (g28896));
AN2X1 gate12264(.O (g18277), .I1 (g1312), .I2 (g16136));
AN2X1 gate12265(.O (g14210), .I1 (g4392), .I2 (g10590));
AN2X1 gate12266(.O (g21910), .I1 (g5016), .I2 (g21468));
AN2X1 gate12267(.O (g26147), .I1 (g6513), .I2 (g25133));
AN2X1 gate12268(.O (g30220), .I1 (g28699), .I2 (g23888));
AN2X1 gate12269(.O (g28666), .I1 (g27567), .I2 (g20625));
AN2X1 gate12270(.O (g33731), .I1 (g33116), .I2 (g19520));
AN2X1 gate12271(.O (g28217), .I1 (g27733), .I2 (g23391));
AN2X1 gate12272(.O (g22123), .I1 (g6609), .I2 (g19277));
AN2X1 gate12273(.O (g21818), .I1 (g3610), .I2 (g20924));
AN4X1 gate12274(.O (g17747), .I1 (g6772), .I2 (g11592), .I3 (g11640), .I4 (I18740));
AN2X1 gate12275(.O (g21979), .I1 (g5559), .I2 (g19074));
AN2X1 gate12276(.O (g16896), .I1 (g262), .I2 (g13120));
AN2X1 gate12277(.O (g27665), .I1 (g26872), .I2 (g23519));
AN2X1 gate12278(.O (g30246), .I1 (g28734), .I2 (g23936));
AN2X1 gate12279(.O (g25871), .I1 (g8334), .I2 (g24804));
AN2X1 gate12280(.O (g20875), .I1 (g16281), .I2 (g4681));
AN2X1 gate12281(.O (g18595), .I1 (g2927), .I2 (g16349));
AN2X1 gate12282(.O (g28478), .I1 (g27007), .I2 (g12345));
AN2X1 gate12283(.O (g18467), .I1 (g2380), .I2 (g15224));
AN2X1 gate12284(.O (g18494), .I1 (g2527), .I2 (g15426));
AN2X1 gate12285(.O (g19500), .I1 (g504), .I2 (g16712));
AN2X1 gate12286(.O (g24219), .I1 (g225), .I2 (g22594));
AN2X1 gate12287(.O (g26858), .I1 (g2970), .I2 (g24540));
AN2X1 gate12288(.O (g21978), .I1 (g5551), .I2 (g19074));
AN2X1 gate12289(.O (g11967), .I1 (g311), .I2 (g7802));
AN2X1 gate12290(.O (g18623), .I1 (g3484), .I2 (g17062));
AN2X1 gate12291(.O (g20218), .I1 (g6541), .I2 (g17815));
AN2X1 gate12292(.O (g30071), .I1 (g29184), .I2 (g12975));
AN2X1 gate12293(.O (g17123), .I1 (g225), .I2 (g13209));
AN2X1 gate12294(.O (g24218), .I1 (g872), .I2 (g22594));
AN2X1 gate12295(.O (g21986), .I1 (g5575), .I2 (g19074));
AN2X1 gate12296(.O (g34071), .I1 (g8854), .I2 (g33799));
AN2X1 gate12297(.O (g18782), .I1 (g5835), .I2 (g18065));
AN2X1 gate12298(.O (g27485), .I1 (g26519), .I2 (g17644));
AN2X1 gate12299(.O (g28556), .I1 (g27431), .I2 (g20374));
AN2X1 gate12300(.O (g29509), .I1 (g1600), .I2 (g28755));
AN2X1 gate12301(.O (g32316), .I1 (g31307), .I2 (g23522));
AN2X1 gate12302(.O (g33405), .I1 (g32354), .I2 (g21398));
AN2X1 gate12303(.O (g21741), .I1 (g15086), .I2 (g20330));
AN2X1 gate12304(.O (g26844), .I1 (g25261), .I2 (g21418));
AN2X1 gate12305(.O (g18419), .I1 (g2051), .I2 (g15373));
AN2X1 gate12306(.O (g27454), .I1 (g26488), .I2 (g17602));
AN2X1 gate12307(.O (g26394), .I1 (g22530), .I2 (g25560));
AN2X1 gate12308(.O (g18352), .I1 (g1798), .I2 (g17955));
AN2X1 gate12309(.O (g29634), .I1 (g2108), .I2 (g29121));
AN2X1 gate12310(.O (g29851), .I1 (g1668), .I2 (g29079));
AN2X1 gate12311(.O (g29872), .I1 (g28401), .I2 (g23333));
AN2X1 gate12312(.O (g28223), .I1 (g27338), .I2 (g17194));
AN2X1 gate12313(.O (g15104), .I1 (g6955), .I2 (g14454));
AN2X1 gate12314(.O (g34754), .I1 (g34677), .I2 (g19602));
AN2X1 gate12315(.O (g18155), .I1 (g15056), .I2 (g17533));
AN2X1 gate12316(.O (g21067), .I1 (g10085), .I2 (g17625));
AN2X1 gate12317(.O (g18418), .I1 (g2122), .I2 (g15373));
AN2X1 gate12318(.O (g18822), .I1 (g6723), .I2 (g15680));
AN2X1 gate12319(.O (g30825), .I1 (g29814), .I2 (g22332));
AN2X1 gate12320(.O (g19613), .I1 (g1437), .I2 (g16713));
AN2X1 gate12321(.O (g32056), .I1 (g27271), .I2 (g31021));
AN2X1 gate12322(.O (g18266), .I1 (g1274), .I2 (g16000));
AN2X1 gate12323(.O (g11010), .I1 (g4698), .I2 (g8933));
AN2X1 gate12324(.O (g34859), .I1 (g16540), .I2 (g34820));
AN2X1 gate12325(.O (g18170), .I1 (g661), .I2 (g17433));
AN4X1 gate12326(.O (I31232), .I1 (g32791), .I2 (g32792), .I3 (g32793), .I4 (g32794));
AN2X1 gate12327(.O (g10677), .I1 (g4141), .I2 (g7611));
AN2X1 gate12328(.O (g22992), .I1 (g1227), .I2 (g19765));
AN2X1 gate12329(.O (g34370), .I1 (g34067), .I2 (g10554));
AN4X1 gate12330(.O (I24674), .I1 (g19919), .I2 (g24019), .I3 (g24020), .I4 (g24021));
AN2X1 gate12331(.O (g21801), .I1 (g3554), .I2 (g20924));
AN2X1 gate12332(.O (g28110), .I1 (g27974), .I2 (g18886));
AN2X1 gate12333(.O (g21735), .I1 (g3057), .I2 (g20330));
AN2X1 gate12334(.O (g21877), .I1 (g6888), .I2 (g19801));
AN2X1 gate12335(.O (g23801), .I1 (g1448), .I2 (g19362));
AN2X1 gate12336(.O (g34858), .I1 (g16540), .I2 (g34816));
AN2X1 gate12337(.O (g30151), .I1 (g28607), .I2 (g21249));
AN2X1 gate12338(.O (g30172), .I1 (g28625), .I2 (g21286));
AN2X1 gate12339(.O (g24915), .I1 (g23087), .I2 (g20158));
AN4X1 gate12340(.O (I31261), .I1 (g30937), .I2 (g31842), .I3 (g32831), .I4 (g32832));
AN2X1 gate12341(.O (g27594), .I1 (g26721), .I2 (g26694));
AN2X1 gate12342(.O (g28531), .I1 (g27722), .I2 (g15608));
AN2X1 gate12343(.O (g17391), .I1 (g9556), .I2 (g14378));
AN2X1 gate12344(.O (g22835), .I1 (g15803), .I2 (g19633));
AN2X1 gate12345(.O (g28178), .I1 (g27019), .I2 (g19397));
AN2X1 gate12346(.O (g18167), .I1 (g718), .I2 (g17433));
AN2X1 gate12347(.O (g18194), .I1 (g843), .I2 (g17821));
AN2X1 gate12348(.O (g18589), .I1 (g2902), .I2 (g16349));
AN2X1 gate12349(.O (g22014), .I1 (g5805), .I2 (g21562));
AN2X1 gate12350(.O (g34367), .I1 (g7404), .I2 (g34042));
AN2X1 gate12351(.O (g31787), .I1 (g21281), .I2 (g29385));
AN2X1 gate12352(.O (g34394), .I1 (g34190), .I2 (g21305));
AN2X1 gate12353(.O (g25071), .I1 (g12804), .I2 (g23478));
AN2X1 gate12354(.O (g33113), .I1 (g31964), .I2 (g22339));
AN2X1 gate12355(.O (g33787), .I1 (g33103), .I2 (g20595));
AN2X1 gate12356(.O (g32342), .I1 (g6545), .I2 (g31579));
AN2X1 gate12357(.O (g29574), .I1 (g2016), .I2 (g28931));
AN2X1 gate12358(.O (g31282), .I1 (g30130), .I2 (g27779));
AN2X1 gate12359(.O (g22007), .I1 (g5770), .I2 (g21562));
AN2X1 gate12360(.O (g15850), .I1 (g3606), .I2 (g14151));
AN3X1 gate12361(.O (g29205), .I1 (g24117), .I2 (I27523), .I3 (I27524));
AN2X1 gate12362(.O (g18588), .I1 (g2970), .I2 (g16349));
AN2X1 gate12363(.O (g18524), .I1 (g2681), .I2 (g15509));
AN2X1 gate12364(.O (g28676), .I1 (g27570), .I2 (g20632));
AN2X1 gate12365(.O (g32145), .I1 (g31609), .I2 (g29977));
AN2X1 gate12366(.O (g14791), .I1 (g1146), .I2 (g10909));
AN2X1 gate12367(.O (g32031), .I1 (g31372), .I2 (g13464));
AN2X1 gate12368(.O (g24467), .I1 (g13761), .I2 (g23047));
AN2X1 gate12369(.O (g27519), .I1 (g26488), .I2 (g17710));
AN2X1 gate12370(.O (g33357), .I1 (g32247), .I2 (g20775));
AN3X1 gate12371(.O (g27185), .I1 (g26190), .I2 (g8302), .I3 (g1917));
AN2X1 gate12372(.O (g25147), .I1 (g20202), .I2 (g23542));
AN2X1 gate12373(.O (g32199), .I1 (g30916), .I2 (g25506));
AN2X1 gate12374(.O (g18401), .I1 (g2036), .I2 (g15373));
AN2X1 gate12375(.O (g28654), .I1 (g1030), .I2 (g27108));
AN2X1 gate12376(.O (g33105), .I1 (g26298), .I2 (g32138));
AN2X1 gate12377(.O (g14168), .I1 (g887), .I2 (g10632));
AN2X1 gate12378(.O (g18477), .I1 (g2429), .I2 (g15426));
AN2X1 gate12379(.O (g26203), .I1 (g1632), .I2 (g25337));
AN2X1 gate12380(.O (g33743), .I1 (g33119), .I2 (g19574));
AN2X1 gate12381(.O (g16802), .I1 (g5567), .I2 (g14807));
AN2X1 gate12382(.O (g18119), .I1 (g475), .I2 (g17015));
AN2X1 gate12383(.O (g27518), .I1 (g26488), .I2 (g17709));
AN2X1 gate12384(.O (g27154), .I1 (g26055), .I2 (g16630));
AN2X1 gate12385(.O (g34319), .I1 (g9535), .I2 (g34156));
AN2X1 gate12386(.O (g32198), .I1 (g4253), .I2 (g31327));
AN2X1 gate12387(.O (g22116), .I1 (g6589), .I2 (g19277));
AN2X1 gate12388(.O (g16730), .I1 (g5212), .I2 (g14723));
AN2X1 gate12389(.O (g24984), .I1 (g22929), .I2 (g12818));
AN2X1 gate12390(.O (g18118), .I1 (g471), .I2 (g17015));
AN2X1 gate12391(.O (g21866), .I1 (g4072), .I2 (g19801));
AN2X1 gate12392(.O (g21917), .I1 (g5092), .I2 (g21468));
AN2X1 gate12393(.O (g30227), .I1 (g28708), .I2 (g23899));
AN2X1 gate12394(.O (g31769), .I1 (g30141), .I2 (g23986));
AN2X1 gate12395(.O (g23917), .I1 (g1472), .I2 (g19428));
AN2X1 gate12396(.O (g33640), .I1 (g33387), .I2 (g18831));
AN4X1 gate12397(.O (g26281), .I1 (g24688), .I2 (g8812), .I3 (g8778), .I4 (g8757));
AN2X1 gate12398(.O (g32330), .I1 (g31320), .I2 (g20631));
AN2X1 gate12399(.O (g29592), .I1 (g28469), .I2 (g11832));
AN2X1 gate12400(.O (g30059), .I1 (g28106), .I2 (g12467));
AN2X1 gate12401(.O (g22720), .I1 (g9253), .I2 (g20619));
AN4X1 gate12402(.O (I31316), .I1 (g29385), .I2 (g32911), .I3 (g32912), .I4 (g32913));
AN2X1 gate12403(.O (g30025), .I1 (g28492), .I2 (g23502));
AN2X1 gate12404(.O (g25151), .I1 (g17719), .I2 (g23549));
AN2X1 gate12405(.O (g16765), .I1 (g6581), .I2 (g15045));
AN2X1 gate12406(.O (g15716), .I1 (g468), .I2 (g13437));
AN2X1 gate12407(.O (g18749), .I1 (g5148), .I2 (g17847));
AN2X1 gate12408(.O (g22041), .I1 (g5957), .I2 (g19147));
AN2X1 gate12409(.O (g26301), .I1 (g2145), .I2 (g25244));
AN2X1 gate12410(.O (g13656), .I1 (g278), .I2 (g11144));
AN2X1 gate12411(.O (g18616), .I1 (g6875), .I2 (g17200));
AN2X1 gate12412(.O (g18313), .I1 (g1430), .I2 (g16931));
AN2X1 gate12413(.O (g33803), .I1 (g33231), .I2 (g20071));
AN3X1 gate12414(.O (g24822), .I1 (g3010), .I2 (g23534), .I3 (I24003));
AN2X1 gate12415(.O (g26120), .I1 (g9809), .I2 (g25293));
AN2X1 gate12416(.O (g30058), .I1 (g29180), .I2 (g12950));
AN2X1 gate12417(.O (g16690), .I1 (g8399), .I2 (g13867));
AN4X1 gate12418(.O (g11144), .I1 (g239), .I2 (g8136), .I3 (g246), .I4 (I14198));
AN2X1 gate12419(.O (g18748), .I1 (g5142), .I2 (g17847));
AN2X1 gate12420(.O (g8643), .I1 (g2927), .I2 (g2922));
AN2X1 gate12421(.O (g25367), .I1 (g6946), .I2 (g22407));
AN4X1 gate12422(.O (I31056), .I1 (g30735), .I2 (g31805), .I3 (g32536), .I4 (g32537));
AN2X1 gate12423(.O (g21706), .I1 (g222), .I2 (g20283));
AN2X1 gate12424(.O (g18276), .I1 (g1351), .I2 (g16136));
AN2X1 gate12425(.O (g18285), .I1 (g1395), .I2 (g16164));
AN2X1 gate12426(.O (g29350), .I1 (g4939), .I2 (g28395));
AN2X1 gate12427(.O (g26146), .I1 (g9892), .I2 (g25334));
AN2X1 gate12428(.O (g30203), .I1 (g28668), .I2 (g23864));
AN2X1 gate12429(.O (g18704), .I1 (g4793), .I2 (g16782));
AN2X1 gate12430(.O (g34203), .I1 (g33726), .I2 (g24537));
AN2X1 gate12431(.O (g18305), .I1 (g1521), .I2 (g16489));
AN2X1 gate12432(.O (g33881), .I1 (g33292), .I2 (g20586));
AN2X1 gate12433(.O (g30044), .I1 (g29174), .I2 (g12944));
AN2X1 gate12434(.O (g18254), .I1 (g1236), .I2 (g16897));
AN2X1 gate12435(.O (g18809), .I1 (g7074), .I2 (g15656));
AN2X1 gate12436(.O (g21923), .I1 (g5029), .I2 (g21468));
AN2X1 gate12437(.O (g22340), .I1 (g19605), .I2 (g13522));
AN2X1 gate12438(.O (g32161), .I1 (g3151), .I2 (g31154));
AN2X1 gate12439(.O (g22035), .I1 (g5933), .I2 (g19147));
AN2X1 gate12440(.O (g28587), .I1 (g27487), .I2 (g20498));
AN2X1 gate12441(.O (g26290), .I1 (g2595), .I2 (g25498));
AN2X1 gate12442(.O (g18466), .I1 (g2389), .I2 (g15224));
AN2X1 gate12443(.O (g23280), .I1 (g19417), .I2 (g20146));
AN2X1 gate12444(.O (g27215), .I1 (g26055), .I2 (g16724));
AN2X1 gate12445(.O (g27501), .I1 (g26400), .I2 (g17673));
AN2X1 gate12446(.O (g15112), .I1 (g4284), .I2 (g14454));
AN4X1 gate12447(.O (I31271), .I1 (g29385), .I2 (g32846), .I3 (g32847), .I4 (g32848));
AN2X1 gate12448(.O (g30281), .I1 (g28850), .I2 (g23992));
AN2X1 gate12449(.O (g18808), .I1 (g6390), .I2 (g15656));
AN3X1 gate12450(.O (g25420), .I1 (g6058), .I2 (g22220), .I3 (I24555));
AN2X1 gate12451(.O (g24194), .I1 (g106), .I2 (g22722));
AN2X1 gate12452(.O (g24589), .I1 (g5471), .I2 (g23630));
AN2X1 gate12453(.O (g34281), .I1 (g34043), .I2 (g19276));
AN2X1 gate12454(.O (g29731), .I1 (g2089), .I2 (g29118));
AN2X1 gate12455(.O (g22142), .I1 (g7957), .I2 (g19140));
AN2X1 gate12456(.O (g27439), .I1 (g232), .I2 (g26831));
AN2X1 gate12457(.O (g34301), .I1 (g34064), .I2 (g19415));
AN2X1 gate12458(.O (g18177), .I1 (g749), .I2 (g17328));
AN2X1 gate12459(.O (g18560), .I1 (g2837), .I2 (g15277));
AN2X1 gate12460(.O (g30120), .I1 (g28576), .I2 (g21051));
AN2X1 gate12461(.O (g28543), .I1 (g27735), .I2 (g15628));
AN2X1 gate12462(.O (g24588), .I1 (g5142), .I2 (g23590));
AN2X1 gate12463(.O (g32087), .I1 (g1291), .I2 (g30825));
AN2X1 gate12464(.O (g34120), .I1 (g33930), .I2 (g25158));
AN4X1 gate12465(.O (I31342), .I1 (g32949), .I2 (g32950), .I3 (g32951), .I4 (g32952));
AN2X1 gate12466(.O (g32258), .I1 (g31624), .I2 (g30303));
AN2X1 gate12467(.O (g28117), .I1 (g8075), .I2 (g27245));
AN2X1 gate12468(.O (g18642), .I1 (g15097), .I2 (g17096));
AN2X1 gate12469(.O (g25059), .I1 (g20870), .I2 (g23460));
AN2X1 gate12470(.O (g33890), .I1 (g33310), .I2 (g20659));
AN2X1 gate12471(.O (g19788), .I1 (g9983), .I2 (g17216));
AN4X1 gate12472(.O (I31031), .I1 (g30614), .I2 (g31801), .I3 (g32499), .I4 (g32500));
AN2X1 gate12473(.O (g16128), .I1 (g14333), .I2 (g14166));
AN2X1 gate12474(.O (g34146), .I1 (g33788), .I2 (g20091));
AN2X1 gate12475(.O (g34738), .I1 (g34660), .I2 (g33442));
AN2X1 gate12476(.O (g33249), .I1 (g32144), .I2 (g20026));
AN2X1 gate12477(.O (g34562), .I1 (g34369), .I2 (g17411));
AN2X1 gate12478(.O (g28569), .I1 (g27453), .I2 (g20433));
AN2X1 gate12479(.O (g21066), .I1 (g10043), .I2 (g17625));
AN2X1 gate12480(.O (g25058), .I1 (g23276), .I2 (g20513));
AN2X1 gate12481(.O (g16245), .I1 (g14278), .I2 (g14708));
AN2X1 gate12482(.O (g32043), .I1 (g31482), .I2 (g16173));
AN3X1 gate12483(.O (g33482), .I1 (g32614), .I2 (I31106), .I3 (I31107));
AN2X1 gate12484(.O (g32244), .I1 (g31609), .I2 (g30297));
AN2X1 gate12485(.O (g31710), .I1 (g29814), .I2 (g19128));
AN2X1 gate12486(.O (g33248), .I1 (g32131), .I2 (g19996));
AN2X1 gate12487(.O (g10676), .I1 (g8506), .I2 (g3774));
AN4X1 gate12488(.O (I27514), .I1 (g24091), .I2 (g24092), .I3 (g24093), .I4 (g24094));
AN2X1 gate12489(.O (g18733), .I1 (g15141), .I2 (g16877));
AN2X1 gate12490(.O (g27083), .I1 (g25819), .I2 (g22456));
AN2X1 gate12491(.O (g27348), .I1 (g26488), .I2 (g17392));
AN2X1 gate12492(.O (g33710), .I1 (g14037), .I2 (g33246));
AN2X1 gate12493(.O (g22130), .I1 (g6637), .I2 (g19277));
AN2X1 gate12494(.O (g27284), .I1 (g9908), .I2 (g26631));
AN2X1 gate12495(.O (g24864), .I1 (g11201), .I2 (g22305));
AN2X1 gate12496(.O (g22193), .I1 (g19880), .I2 (g20682));
AN2X1 gate12497(.O (g28242), .I1 (g27769), .I2 (g23626));
AN2X1 gate12498(.O (g21876), .I1 (g4119), .I2 (g19801));
AN2X1 gate12499(.O (g21885), .I1 (g4122), .I2 (g19801));
AN2X1 gate12500(.O (g26547), .I1 (g13283), .I2 (g25027));
AN2X1 gate12501(.O (g10654), .I1 (g3085), .I2 (g8434));
AN2X1 gate12502(.O (g11023), .I1 (g9669), .I2 (g5084));
AN2X1 gate12503(.O (g15857), .I1 (g3199), .I2 (g14038));
AN2X1 gate12504(.O (g23885), .I1 (g4132), .I2 (g19513));
AN2X1 gate12505(.O (g27304), .I1 (g2273), .I2 (g26682));
AN2X1 gate12506(.O (g24749), .I1 (g17511), .I2 (g22432));
AN2X1 gate12507(.O (g32069), .I1 (g10878), .I2 (g30735));
AN2X1 gate12508(.O (g12284), .I1 (g1532), .I2 (g7557));
AN2X1 gate12509(.O (g14654), .I1 (g7178), .I2 (g10476));
AN2X1 gate12510(.O (g24313), .I1 (g4504), .I2 (g22228));
AN2X1 gate12511(.O (g22165), .I1 (g15594), .I2 (g18903));
AN2X1 gate12512(.O (g18630), .I1 (g3689), .I2 (g17226));
AN2X1 gate12513(.O (g21854), .I1 (g3921), .I2 (g21070));
AN2X1 gate12514(.O (g15793), .I1 (g3219), .I2 (g13873));
AN2X1 gate12515(.O (g18693), .I1 (g4717), .I2 (g16053));
AN2X1 gate12516(.O (g23854), .I1 (g4093), .I2 (g19506));
AN2X1 gate12517(.O (g31778), .I1 (g21369), .I2 (g29385));
AN2X1 gate12518(.O (g24748), .I1 (g17656), .I2 (g22457));
AN4X1 gate12519(.O (g26226), .I1 (g24688), .I2 (g8812), .I3 (g10658), .I4 (g10627));
AN2X1 gate12520(.O (g32068), .I1 (g31515), .I2 (g10862));
AN2X1 gate12521(.O (g33081), .I1 (g32388), .I2 (g18875));
AN2X1 gate12522(.O (g17193), .I1 (g2504), .I2 (g13023));
AN2X1 gate12523(.O (g21763), .I1 (g3223), .I2 (g20785));
AN2X1 gate12524(.O (g18166), .I1 (g655), .I2 (g17433));
AN2X1 gate12525(.O (g24285), .I1 (g4388), .I2 (g22550));
AN2X1 gate12526(.O (g25902), .I1 (g24398), .I2 (g19373));
AN2X1 gate12527(.O (g18665), .I1 (g4584), .I2 (g17367));
AN4X1 gate12528(.O (I31132), .I1 (g32645), .I2 (g32646), .I3 (g32647), .I4 (g32648));
AN2X1 gate12529(.O (g31786), .I1 (g30189), .I2 (g24010));
AN2X1 gate12530(.O (g25957), .I1 (g17190), .I2 (g24960));
AN2X1 gate12531(.O (g24704), .I1 (g17593), .I2 (g22384));
AN3X1 gate12532(.O (g25377), .I1 (g5712), .I2 (g22210), .I3 (I24530));
AN2X1 gate12533(.O (g33786), .I1 (g33130), .I2 (g20572));
AN2X1 gate12534(.O (g24305), .I1 (g4477), .I2 (g22228));
AN2X1 gate12535(.O (g16737), .I1 (g6645), .I2 (g15042));
AN2X1 gate12536(.O (g26572), .I1 (g7443), .I2 (g24439));
AN2X1 gate12537(.O (g22006), .I1 (g5767), .I2 (g21562));
AN2X1 gate12538(.O (g28639), .I1 (g27767), .I2 (g20597));
AN3X1 gate12539(.O (g24900), .I1 (g3752), .I2 (g23582), .I3 (I24067));
AN2X1 gate12540(.O (g33647), .I1 (g33390), .I2 (g18878));
AN2X1 gate12541(.O (g32337), .I1 (g31465), .I2 (g20663));
AN2X1 gate12542(.O (g27139), .I1 (g26055), .I2 (g16608));
AN3X1 gate12543(.O (g28293), .I1 (g7424), .I2 (g2495), .I3 (g27474));
AN2X1 gate12544(.O (g33356), .I1 (g32245), .I2 (g20772));
AN2X1 gate12545(.O (g22863), .I1 (g9547), .I2 (g20388));
AN2X1 gate12546(.O (g27653), .I1 (g26549), .I2 (g15562));
AN2X1 gate12547(.O (g28638), .I1 (g27551), .I2 (g20583));
AN2X1 gate12548(.O (g32171), .I1 (g31706), .I2 (g27800));
AN4X1 gate12549(.O (I31161), .I1 (g30614), .I2 (g31824), .I3 (g32687), .I4 (g32688));
AN2X1 gate12550(.O (g18476), .I1 (g2433), .I2 (g15426));
AN2X1 gate12551(.O (g18485), .I1 (g2465), .I2 (g15426));
AN2X1 gate12552(.O (g29787), .I1 (g28334), .I2 (g23249));
AN2X1 gate12553(.O (g26127), .I1 (g2236), .I2 (g25119));
AN2X1 gate12554(.O (g27138), .I1 (g26055), .I2 (g16607));
AN2X1 gate12555(.O (g28265), .I1 (g11367), .I2 (g27989));
AN2X1 gate12556(.O (g34661), .I1 (g34575), .I2 (g18907));
AN2X1 gate12557(.O (g18555), .I1 (g2834), .I2 (g15277));
AN2X1 gate12558(.O (g18454), .I1 (g2303), .I2 (g15224));
AN3X1 gate12559(.O (g25290), .I1 (g5022), .I2 (g22173), .I3 (I24482));
AN2X1 gate12560(.O (g14216), .I1 (g7631), .I2 (g10608));
AN2X1 gate12561(.O (g21916), .I1 (g5084), .I2 (g21468));
AN2X1 gate12562(.O (g30226), .I1 (g28707), .I2 (g23898));
AN2X1 gate12563(.O (g18570), .I1 (g2848), .I2 (g16349));
AN2X1 gate12564(.O (g18712), .I1 (g4843), .I2 (g15915));
AN2X1 gate12565(.O (g33233), .I1 (g32094), .I2 (g23005));
AN2X1 gate12566(.O (g31182), .I1 (g30240), .I2 (g20682));
AN2X1 gate12567(.O (g31672), .I1 (g29814), .I2 (g19050));
AN2X1 gate12568(.O (g27333), .I1 (g10180), .I2 (g26765));
AN2X1 gate12569(.O (g24642), .I1 (g8290), .I2 (g22898));
AN2X1 gate12570(.O (g34226), .I1 (g33914), .I2 (g21467));
AN2X1 gate12571(.O (g14587), .I1 (g10584), .I2 (g10567));
AN2X1 gate12572(.O (g29743), .I1 (g28206), .I2 (g10233));
AN4X1 gate12573(.O (I31087), .I1 (g32580), .I2 (g32581), .I3 (g32582), .I4 (g32583));
AN2X1 gate12574(.O (g34715), .I1 (g34570), .I2 (g33375));
AN2X1 gate12575(.O (g34481), .I1 (g34404), .I2 (g18916));
AN2X1 gate12576(.O (g23314), .I1 (g9104), .I2 (g19200));
AN2X1 gate12577(.O (g32425), .I1 (g31668), .I2 (g21604));
AN2X1 gate12578(.O (g26103), .I1 (g2185), .I2 (g25100));
AN2X1 gate12579(.O (g34572), .I1 (g34387), .I2 (g33326));
AN2X1 gate12580(.O (g10543), .I1 (g8238), .I2 (g437));
AN2X1 gate12581(.O (g26095), .I1 (g11923), .I2 (g25090));
AN2X1 gate12582(.O (g27963), .I1 (g25952), .I2 (g16047));
AN2X1 gate12583(.O (g23076), .I1 (g19128), .I2 (g9104));
AN2X1 gate12584(.O (g29640), .I1 (g28498), .I2 (g8125));
AN2X1 gate12585(.O (g25366), .I1 (g7733), .I2 (g22406));
AN2X1 gate12586(.O (g29769), .I1 (g28319), .I2 (g23237));
AN2X1 gate12587(.O (g18239), .I1 (g1135), .I2 (g16326));
AN2X1 gate12588(.O (g21721), .I1 (g385), .I2 (g21037));
AN2X1 gate12589(.O (g33331), .I1 (g32216), .I2 (g20607));
AN2X1 gate12590(.O (g27664), .I1 (g1024), .I2 (g25911));
AN2X1 gate12591(.O (g18567), .I1 (g2894), .I2 (g16349));
AN2X1 gate12592(.O (g18594), .I1 (g12858), .I2 (g16349));
AN2X1 gate12593(.O (g31513), .I1 (g2606), .I2 (g29318));
AN2X1 gate12594(.O (g32010), .I1 (g31785), .I2 (g22303));
AN3X1 gate12595(.O (g33513), .I1 (g32837), .I2 (I31261), .I3 (I31262));
AN2X1 gate12596(.O (g29803), .I1 (g28414), .I2 (g26836));
AN2X1 gate12597(.O (g18238), .I1 (g1152), .I2 (g16326));
AN2X1 gate12598(.O (g26181), .I1 (g2652), .I2 (g25157));
AN2X1 gate12599(.O (g26671), .I1 (g316), .I2 (g24429));
AN2X1 gate12600(.O (g28586), .I1 (g27484), .I2 (g20497));
AN2X1 gate12601(.O (g24630), .I1 (g23255), .I2 (g14149));
AN2X1 gate12602(.O (g31961), .I1 (g31751), .I2 (g22154));
AN2X1 gate12603(.O (g33897), .I1 (g33315), .I2 (g20777));
AN4X1 gate12604(.O (g17781), .I1 (g6772), .I2 (g11592), .I3 (g6789), .I4 (I18785));
AN2X1 gate12605(.O (g31505), .I1 (g30195), .I2 (g24379));
AN2X1 gate12606(.O (g28442), .I1 (g27278), .I2 (g20072));
AN3X1 gate12607(.O (g33505), .I1 (g32779), .I2 (I31221), .I3 (I31222));
AN2X1 gate12608(.O (g18382), .I1 (g1936), .I2 (g15171));
AN2X1 gate12609(.O (g24009), .I1 (g19671), .I2 (g10971));
AN2X1 gate12610(.O (g33404), .I1 (g32353), .I2 (g21397));
AN2X1 gate12611(.O (g29881), .I1 (g2040), .I2 (g29150));
AN2X1 gate12612(.O (g21773), .I1 (g3263), .I2 (g20785));
AN2X1 gate12613(.O (g18519), .I1 (g2648), .I2 (g15509));
AN2X1 gate12614(.O (g11016), .I1 (g4888), .I2 (g8984));
AN2X1 gate12615(.O (g21942), .I1 (g5236), .I2 (g18997));
AN2X1 gate12616(.O (g13525), .I1 (g10019), .I2 (g11911));
AN2X1 gate12617(.O (g18176), .I1 (g732), .I2 (g17328));
AN2X1 gate12618(.O (g18185), .I1 (g790), .I2 (g17328));
AN2X1 gate12619(.O (g22063), .I1 (g6109), .I2 (g21611));
AN2X1 gate12620(.O (g18675), .I1 (g4349), .I2 (g15758));
AN2X1 gate12621(.O (g34385), .I1 (g34168), .I2 (g20642));
AN2X1 gate12622(.O (g33717), .I1 (g14092), .I2 (g33306));
AN2X1 gate12623(.O (g24008), .I1 (g7909), .I2 (g19502));
AN2X1 gate12624(.O (g32086), .I1 (g7597), .I2 (g30735));
AN2X1 gate12625(.O (g30095), .I1 (g28545), .I2 (g20768));
AN2X1 gate12626(.O (g31212), .I1 (g20028), .I2 (g29669));
AN2X1 gate12627(.O (g28116), .I1 (g27366), .I2 (g26183));
AN2X1 gate12628(.O (g18518), .I1 (g2657), .I2 (g15509));
AN2X1 gate12629(.O (g18154), .I1 (g622), .I2 (g17533));
AN2X1 gate12630(.O (g27312), .I1 (g12019), .I2 (g26700));
AN2X1 gate12631(.O (g24892), .I1 (g11559), .I2 (g23264));
AN4X1 gate12632(.O (g26190), .I1 (g25357), .I2 (g11724), .I3 (g7586), .I4 (g11686));
AN2X1 gate12633(.O (g24485), .I1 (g10710), .I2 (g22319));
AN2X1 gate12634(.O (g24476), .I1 (g18879), .I2 (g22330));
AN4X1 gate12635(.O (I31337), .I1 (g32942), .I2 (g32943), .I3 (g32944), .I4 (g32945));
AN2X1 gate12636(.O (g16611), .I1 (g5583), .I2 (g14727));
AN2X1 gate12637(.O (g27115), .I1 (g26026), .I2 (g16526));
AN2X1 gate12638(.O (g11893), .I1 (g1668), .I2 (g7268));
AN4X1 gate12639(.O (g13830), .I1 (g11543), .I2 (g11424), .I3 (g11395), .I4 (I16143));
AN2X1 gate12640(.O (g22873), .I1 (g19854), .I2 (g19683));
AN2X1 gate12641(.O (g25551), .I1 (g23822), .I2 (g21511));
AN2X1 gate12642(.O (g18637), .I1 (g3821), .I2 (g17096));
AN2X1 gate12643(.O (g25572), .I1 (I24699), .I2 (I24700));
AN4X1 gate12644(.O (I31171), .I1 (g31528), .I2 (g31826), .I3 (g32701), .I4 (g32702));
AN2X1 gate12645(.O (g30181), .I1 (g28636), .I2 (g23821));
AN2X1 gate12646(.O (g30671), .I1 (g29319), .I2 (g22317));
AN2X1 gate12647(.O (g18935), .I1 (g4322), .I2 (g15574));
AN2X1 gate12648(.O (g32322), .I1 (g31308), .I2 (g20605));
AN2X1 gate12649(.O (g24555), .I1 (g23184), .I2 (g21024));
AN2X1 gate12650(.O (g29662), .I1 (g1848), .I2 (g29049));
AN2X1 gate12651(.O (g9217), .I1 (g632), .I2 (g626));
AN2X1 gate12652(.O (g21734), .I1 (g3040), .I2 (g20330));
AN2X1 gate12653(.O (g32159), .I1 (g31658), .I2 (g30040));
AN2X1 gate12654(.O (g24712), .I1 (g19592), .I2 (g23001));
AN2X1 gate12655(.O (g29890), .I1 (g28419), .I2 (g23355));
AN2X1 gate12656(.O (g24914), .I1 (g8721), .I2 (g23301));
AN2X1 gate12657(.O (g21839), .I1 (g3763), .I2 (g20453));
AN2X1 gate12658(.O (g21930), .I1 (g5180), .I2 (g18997));
AN2X1 gate12659(.O (g25127), .I1 (g13997), .I2 (g23524));
AN2X1 gate12660(.O (g21993), .I1 (g5603), .I2 (g19074));
AN2X1 gate12661(.O (g32158), .I1 (g31658), .I2 (g30022));
AN2X1 gate12662(.O (g22209), .I1 (g19907), .I2 (g20751));
AN2X1 gate12663(.O (g15856), .I1 (g9056), .I2 (g14223));
AN3X1 gate12664(.O (g15995), .I1 (g13314), .I2 (g1157), .I3 (g10666));
AN2X1 gate12665(.O (g33723), .I1 (g14091), .I2 (g33299));
AN2X1 gate12666(.O (g28237), .I1 (g9492), .I2 (g27597));
AN2X1 gate12667(.O (g21838), .I1 (g3747), .I2 (g20453));
AN2X1 gate12668(.O (g22834), .I1 (g102), .I2 (g19630));
AN2X1 gate12669(.O (g15880), .I1 (g3211), .I2 (g13980));
AN2X1 gate12670(.O (g31149), .I1 (g29508), .I2 (g23021));
AN2X1 gate12671(.O (g21965), .I1 (g15149), .I2 (g21514));
AN2X1 gate12672(.O (g26088), .I1 (g6545), .I2 (g25080));
AN2X1 gate12673(.O (g26024), .I1 (g2619), .I2 (g25039));
AN2X1 gate12674(.O (g22208), .I1 (g19906), .I2 (g20739));
AN2X1 gate12675(.O (g29710), .I1 (g2380), .I2 (g29094));
AN3X1 gate12676(.O (g28035), .I1 (g24103), .I2 (I26530), .I3 (I26531));
AN2X1 gate12677(.O (g29552), .I1 (g2223), .I2 (g28579));
AN2X1 gate12678(.O (g33433), .I1 (g32238), .I2 (g29694));
AN2X1 gate12679(.O (g23131), .I1 (g13919), .I2 (g19930));
AN2X1 gate12680(.O (g32295), .I1 (g27931), .I2 (g31376));
AN2X1 gate12681(.O (g10841), .I1 (g8509), .I2 (g8567));
AN3X1 gate12682(.O (g29204), .I1 (g24110), .I2 (I27518), .I3 (I27519));
AN2X1 gate12683(.O (g31148), .I1 (g2661), .I2 (g30055));
AN2X1 gate12684(.O (g30190), .I1 (g28646), .I2 (g23842));
AN2X1 gate12685(.O (g13042), .I1 (g433), .I2 (g11048));
AN2X1 gate12686(.O (g16199), .I1 (g3614), .I2 (g14051));
AN2X1 gate12687(.O (g18215), .I1 (g943), .I2 (g15979));
AN2X1 gate12688(.O (g25103), .I1 (g4927), .I2 (g22908));
AN2X1 gate12689(.O (g27184), .I1 (g26628), .I2 (g13756));
AN2X1 gate12690(.O (g16736), .I1 (g6303), .I2 (g15036));
AN2X1 gate12691(.O (g18501), .I1 (g12854), .I2 (g15509));
AN2X1 gate12692(.O (g18729), .I1 (g15139), .I2 (g16821));
AN2X1 gate12693(.O (g22021), .I1 (g5869), .I2 (g19147));
AN2X1 gate12694(.O (g27674), .I1 (g26873), .I2 (g23543));
AN2X1 gate12695(.O (g25980), .I1 (g1926), .I2 (g25006));
AN2X1 gate12696(.O (g18577), .I1 (g2988), .I2 (g16349));
AN2X1 gate12697(.O (g33104), .I1 (g26296), .I2 (g32137));
AN2X1 gate12698(.O (g25095), .I1 (g23319), .I2 (g20556));
AN2X1 gate12699(.O (g33811), .I1 (g33439), .I2 (g17573));
AN2X1 gate12700(.O (g33646), .I1 (g33389), .I2 (g18876));
AN2X1 gate12701(.O (g19767), .I1 (g16810), .I2 (g14203));
AN2X1 gate12702(.O (g32336), .I1 (g31596), .I2 (g11842));
AN2X1 gate12703(.O (g34520), .I1 (g34294), .I2 (g19505));
AN2X1 gate12704(.O (g23619), .I1 (g19453), .I2 (g13045));
AN2X1 gate12705(.O (g33343), .I1 (g32227), .I2 (g20665));
AN2X1 gate12706(.O (g21557), .I1 (g12980), .I2 (g15674));
AN2X1 gate12707(.O (g18728), .I1 (g4939), .I2 (g16821));
AN2X1 gate12708(.O (g18439), .I1 (g2250), .I2 (g18008));
AN2X1 gate12709(.O (g30089), .I1 (g28538), .I2 (g20709));
AN2X1 gate12710(.O (g24941), .I1 (g23171), .I2 (g20190));
AN2X1 gate12711(.O (g26126), .I1 (g1959), .I2 (g25118));
AN2X1 gate12712(.O (g30211), .I1 (g28685), .I2 (g23878));
AN2X1 gate12713(.O (g11939), .I1 (g2361), .I2 (g7380));
AN2X1 gate12714(.O (g23618), .I1 (g19388), .I2 (g11917));
AN2X1 gate12715(.O (g25181), .I1 (g23405), .I2 (g20696));
AN3X1 gate12716(.O (g34089), .I1 (g22957), .I2 (g9104), .I3 (g33744));
AN2X1 gate12717(.O (g16843), .I1 (g6251), .I2 (g14864));
AN2X1 gate12718(.O (g18438), .I1 (g2236), .I2 (g18008));
AN2X1 gate12719(.O (g34211), .I1 (g33891), .I2 (g21349));
AN2X1 gate12720(.O (g26250), .I1 (g1902), .I2 (g25429));
AN2X1 gate12721(.O (g13383), .I1 (g4765), .I2 (g11797));
AN2X1 gate12722(.O (g24675), .I1 (g17568), .I2 (g22342));
AN2X1 gate12723(.O (g29647), .I1 (g28934), .I2 (g22457));
AN2X1 gate12724(.O (g30024), .I1 (g28497), .I2 (g23501));
AN2X1 gate12725(.O (g33369), .I1 (g32277), .I2 (g21060));
AN3X1 gate12726(.O (I24048), .I1 (g3034), .I2 (g3040), .I3 (g8426));
AN2X1 gate12727(.O (g17726), .I1 (g1467), .I2 (g13315));
AN2X1 gate12728(.O (g16764), .I1 (g6307), .I2 (g14776));
AN3X1 gate12729(.O (g34088), .I1 (g33736), .I2 (g9104), .I3 (g18957));
AN2X1 gate12730(.O (g13030), .I1 (g429), .I2 (g11048));
AN2X1 gate12731(.O (g22073), .I1 (g6235), .I2 (g19210));
AN2X1 gate12732(.O (g18349), .I1 (g1768), .I2 (g17955));
AN2X1 gate12733(.O (g14586), .I1 (g11953), .I2 (g11970));
AN2X1 gate12734(.O (g13294), .I1 (g1564), .I2 (g11513));
AN4X1 gate12735(.O (I31086), .I1 (g31554), .I2 (g31811), .I3 (g32578), .I4 (g32579));
AN2X1 gate12736(.O (g29380), .I1 (g28134), .I2 (g19396));
AN2X1 gate12737(.O (g33368), .I1 (g32275), .I2 (g21057));
AN2X1 gate12738(.O (g34860), .I1 (g16540), .I2 (g34823));
AN2X1 gate12739(.O (g16869), .I1 (g6259), .I2 (g14902));
AN2X1 gate12740(.O (g27692), .I1 (g26392), .I2 (g20697));
AN2X1 gate12741(.O (g28130), .I1 (g27353), .I2 (g23063));
AN2X1 gate12742(.O (g28193), .I1 (g8851), .I2 (g27629));
AN2X1 gate12743(.O (g26339), .I1 (g225), .I2 (g24836));
AN2X1 gate12744(.O (g25931), .I1 (g24574), .I2 (g19477));
AN2X1 gate12745(.O (g18906), .I1 (g13568), .I2 (g16264));
AN2X1 gate12746(.O (g18348), .I1 (g1744), .I2 (g17955));
AN2X1 gate12747(.O (g24637), .I1 (g16586), .I2 (g22884));
AN2X1 gate12748(.O (g19521), .I1 (g513), .I2 (g16739));
AN2X1 gate12749(.O (g22122), .I1 (g6601), .I2 (g19277));
AN3X1 gate12750(.O (g12692), .I1 (g10323), .I2 (g3522), .I3 (g3530));
AN2X1 gate12751(.O (g12761), .I1 (g969), .I2 (g7567));
AN2X1 gate12752(.O (g18284), .I1 (g15071), .I2 (g16164));
AN2X1 gate12753(.O (g16868), .I1 (g5813), .I2 (g14297));
AN2X1 gate12754(.O (g34497), .I1 (g34275), .I2 (g33072));
AN2X1 gate12755(.O (g28165), .I1 (g27018), .I2 (g22455));
AN2X1 gate12756(.O (g28523), .I1 (g27704), .I2 (g15585));
AN2X1 gate12757(.O (g18304), .I1 (g1542), .I2 (g16489));
AN2X1 gate12758(.O (g29182), .I1 (g27163), .I2 (g12730));
AN2X1 gate12759(.O (g29651), .I1 (g2537), .I2 (g29134));
AN2X1 gate12760(.O (g33412), .I1 (g32362), .I2 (g21411));
AN4X1 gate12761(.O (I31322), .I1 (g32921), .I2 (g32922), .I3 (g32923), .I4 (g32924));
AN2X1 gate12762(.O (g16161), .I1 (g5841), .I2 (g14297));
AN2X1 gate12763(.O (g15611), .I1 (g471), .I2 (g13437));
AN2X1 gate12764(.O (g15722), .I1 (g464), .I2 (g13437));
AN2X1 gate12765(.O (g18622), .I1 (g3480), .I2 (g17062));
AN2X1 gate12766(.O (g22034), .I1 (g5929), .I2 (g19147));
AN2X1 gate12767(.O (g15080), .I1 (g12855), .I2 (g12983));
AN2X1 gate12768(.O (g18566), .I1 (g2860), .I2 (g16349));
AN2X1 gate12769(.O (g30126), .I1 (g28582), .I2 (g21058));
AN2X1 gate12770(.O (g14615), .I1 (g10604), .I2 (g10587));
AN2X1 gate12771(.O (g27214), .I1 (g26026), .I2 (g13901));
AN2X1 gate12772(.O (g34700), .I1 (g34535), .I2 (g20129));
AN2X1 gate12773(.O (g31229), .I1 (g30288), .I2 (g23949));
AN3X1 gate12774(.O (g10720), .I1 (g2704), .I2 (g10219), .I3 (g2689));
AN2X1 gate12775(.O (g21815), .I1 (g3598), .I2 (g20924));
AN2X1 gate12776(.O (g30250), .I1 (g28744), .I2 (g23939));
AN2X1 gate12777(.O (g27329), .I1 (g12052), .I2 (g26743));
AN2X1 gate12778(.O (g32309), .I1 (g5160), .I2 (g31528));
AN2X1 gate12779(.O (g27207), .I1 (g26055), .I2 (g16692));
AN2X1 gate12780(.O (g33896), .I1 (g33314), .I2 (g20771));
AN2X1 gate12781(.O (g31228), .I1 (g20028), .I2 (g29713));
AN2X1 gate12782(.O (g27539), .I1 (g26576), .I2 (g17745));
AN2X1 gate12783(.O (g29331), .I1 (g29143), .I2 (g22169));
AN2X1 gate12784(.O (g32224), .I1 (g4300), .I2 (g31327));
AN2X1 gate12785(.O (g34658), .I1 (g34574), .I2 (g18896));
AN2X1 gate12786(.O (g23187), .I1 (g13989), .I2 (g20010));
AN2X1 gate12787(.O (g26855), .I1 (g2960), .I2 (g24535));
AN2X1 gate12788(.O (g21975), .I1 (g5523), .I2 (g19074));
AN2X1 gate12789(.O (g27328), .I1 (g12482), .I2 (g26736));
AN2X1 gate12790(.O (g25089), .I1 (g23317), .I2 (g20553));
AN2X1 gate12791(.O (g32308), .I1 (g31293), .I2 (g23503));
AN2X1 gate12792(.O (g20215), .I1 (g16479), .I2 (g10476));
AN2X1 gate12793(.O (g29513), .I1 (g28448), .I2 (g14095));
AN2X1 gate12794(.O (g18139), .I1 (g542), .I2 (g17249));
AN2X1 gate12795(.O (g27538), .I1 (g26549), .I2 (g14744));
AN2X1 gate12796(.O (g18653), .I1 (g4176), .I2 (g16249));
AN2X1 gate12797(.O (g24501), .I1 (g14000), .I2 (g23182));
AN2X1 gate12798(.O (g24729), .I1 (g22719), .I2 (g23018));
AN2X1 gate12799(.O (g25088), .I1 (g17601), .I2 (g23491));
AN2X1 gate12800(.O (g17292), .I1 (g1075), .I2 (g13093));
AN4X1 gate12801(.O (g11160), .I1 (g6336), .I2 (g7074), .I3 (g6322), .I4 (g10003));
AN2X1 gate12802(.O (g17153), .I1 (g6311), .I2 (g14943));
AN3X1 gate12803(.O (I24033), .I1 (g8219), .I2 (g8443), .I3 (g3747));
AN2X1 gate12804(.O (g18138), .I1 (g546), .I2 (g17249));
AN4X1 gate12805(.O (I26531), .I1 (g24099), .I2 (g24100), .I3 (g24101), .I4 (g24102));
AN2X1 gate12806(.O (g21937), .I1 (g5208), .I2 (g18997));
AN3X1 gate12807(.O (I17552), .I1 (g13156), .I2 (g11450), .I3 (g11498));
AN2X1 gate12808(.O (g34338), .I1 (g34099), .I2 (g19905));
AN2X1 gate12809(.O (g24728), .I1 (g16513), .I2 (g23017));
AN4X1 gate12810(.O (g16244), .I1 (g11547), .I2 (g11592), .I3 (g6789), .I4 (I17585));
AN4X1 gate12811(.O (I31336), .I1 (g31672), .I2 (g31855), .I3 (g32940), .I4 (g32941));
AN2X1 gate12812(.O (g14035), .I1 (g699), .I2 (g11048));
AN2X1 gate12813(.O (g15650), .I1 (g8362), .I2 (g13413));
AN2X1 gate12814(.O (g34969), .I1 (g34960), .I2 (g19570));
AN2X1 gate12815(.O (g10684), .I1 (g7998), .I2 (g411));
AN2X1 gate12816(.O (g28703), .I1 (g27925), .I2 (g20680));
AN2X1 gate12817(.O (g18636), .I1 (g3817), .I2 (g17096));
AN2X1 gate12818(.O (g18415), .I1 (g2108), .I2 (g15373));
AN2X1 gate12819(.O (g31310), .I1 (g30157), .I2 (g27886));
AN2X1 gate12820(.O (g18333), .I1 (g1691), .I2 (g17873));
AN2X1 gate12821(.O (g30060), .I1 (g29146), .I2 (g10581));
AN2X1 gate12822(.O (g21791), .I1 (g3368), .I2 (g20391));
AN2X1 gate12823(.O (g28253), .I1 (g23719), .I2 (g27700));
AN2X1 gate12824(.O (g21884), .I1 (g4104), .I2 (g19801));
AN2X1 gate12825(.O (g11915), .I1 (g1802), .I2 (g7315));
AN2X1 gate12826(.O (g34968), .I1 (g34952), .I2 (g23203));
AN2X1 gate12827(.O (g23884), .I1 (g4119), .I2 (g19510));
AN2X1 gate12828(.O (g30197), .I1 (g28661), .I2 (g23859));
AN2X1 gate12829(.O (g31959), .I1 (g4907), .I2 (g30673));
AN2X1 gate12830(.O (g33379), .I1 (g30984), .I2 (g32364));
AN4X1 gate12831(.O (g19462), .I1 (g7850), .I2 (g14182), .I3 (g14177), .I4 (g16646));
AN2X1 gate12832(.O (g25126), .I1 (g16839), .I2 (g23523));
AN2X1 gate12833(.O (g25987), .I1 (g9501), .I2 (g25015));
AN4X1 gate12834(.O (I31017), .I1 (g32480), .I2 (g32481), .I3 (g32482), .I4 (g32483));
AN2X1 gate12835(.O (g13277), .I1 (g3195), .I2 (g11432));
AN2X1 gate12836(.O (g28236), .I1 (g8515), .I2 (g27971));
AN2X1 gate12837(.O (g34870), .I1 (g34820), .I2 (g19882));
AN2X1 gate12838(.O (g34527), .I1 (g34303), .I2 (g19603));
AN2X1 gate12839(.O (g24284), .I1 (g4375), .I2 (g22550));
AN2X1 gate12840(.O (g18664), .I1 (g4332), .I2 (g17367));
AN2X1 gate12841(.O (g27235), .I1 (g25910), .I2 (g19579));
AN2X1 gate12842(.O (g24304), .I1 (g12875), .I2 (g22228));
AN2X1 gate12843(.O (g26819), .I1 (g106), .I2 (g24490));
AN2X1 gate12844(.O (g27683), .I1 (g25770), .I2 (g23567));
AN2X1 gate12845(.O (g24622), .I1 (g19856), .I2 (g22866));
AN3X1 gate12846(.O (g33742), .I1 (g7828), .I2 (g33142), .I3 (I31600));
AN2X1 gate12847(.O (g26257), .I1 (g4253), .I2 (g25197));
AN2X1 gate12848(.O (g31944), .I1 (g31745), .I2 (g22146));
AN2X1 gate12849(.O (g11037), .I1 (g6128), .I2 (g9184));
AN2X1 gate12850(.O (g18576), .I1 (g2868), .I2 (g16349));
AN2X1 gate12851(.O (g18585), .I1 (g2960), .I2 (g16349));
AN2X1 gate12852(.O (g14193), .I1 (g7178), .I2 (g10590));
AN2X1 gate12853(.O (g18484), .I1 (g2491), .I2 (g15426));
AN2X1 gate12854(.O (g22109), .I1 (g6455), .I2 (g18833));
AN2X1 gate12855(.O (g32260), .I1 (g31250), .I2 (g20385));
AN3X1 gate12856(.O (g28264), .I1 (g7315), .I2 (g1802), .I3 (g27416));
AN2X1 gate12857(.O (g34503), .I1 (g34278), .I2 (g19437));
AN2X1 gate12858(.O (g34867), .I1 (g34826), .I2 (g20145));
AN2X1 gate12859(.O (g25969), .I1 (g9310), .I2 (g24987));
AN2X1 gate12860(.O (g18554), .I1 (g2831), .I2 (g15277));
AN2X1 gate12861(.O (g29620), .I1 (g2399), .I2 (g29097));
AN2X1 gate12862(.O (g33681), .I1 (g33129), .I2 (g7991));
AN2X1 gate12863(.O (g22108), .I1 (g6439), .I2 (g18833));
AN2X1 gate12864(.O (g18609), .I1 (g3147), .I2 (g16987));
AN2X1 gate12865(.O (g27414), .I1 (g255), .I2 (g26827));
AN2X1 gate12866(.O (g32195), .I1 (g30734), .I2 (g25451));
AN2X1 gate12867(.O (g24139), .I1 (g17619), .I2 (g21653));
AN2X1 gate12868(.O (g25968), .I1 (g25215), .I2 (g20739));
AN2X1 gate12869(.O (g18312), .I1 (g1579), .I2 (g16931));
AN2X1 gate12870(.O (g33802), .I1 (g33097), .I2 (g14545));
AN2X1 gate12871(.O (g33429), .I1 (g32231), .I2 (g29676));
AN2X1 gate12872(.O (g33857), .I1 (g33267), .I2 (g20445));
AN2X1 gate12873(.O (g29646), .I1 (g1816), .I2 (g28675));
AN3X1 gate12874(.O (g30315), .I1 (g29182), .I2 (g7028), .I3 (g5644));
AN2X1 gate12875(.O (g34581), .I1 (g22864), .I2 (g34312));
AN2X1 gate12876(.O (g18608), .I1 (g15087), .I2 (g16987));
AN2X1 gate12877(.O (g27407), .I1 (g26488), .I2 (g17522));
AN2X1 gate12878(.O (g18115), .I1 (g460), .I2 (g17015));
AN4X1 gate12879(.O (I27534), .I1 (g28039), .I2 (g24128), .I3 (g24129), .I4 (g24130));
AN4X1 gate12880(.O (g33730), .I1 (g7202), .I2 (g4621), .I3 (g33127), .I4 (g4633));
AN2X1 gate12881(.O (g32016), .I1 (g8522), .I2 (g31138));
AN2X1 gate12882(.O (g33428), .I1 (g32230), .I2 (g29672));
AN2X1 gate12883(.O (g34707), .I1 (g34544), .I2 (g20579));
AN2X1 gate12884(.O (g30202), .I1 (g28667), .I2 (g23863));
AN2X1 gate12885(.O (g25870), .I1 (g24840), .I2 (g16182));
AN2X1 gate12886(.O (g30257), .I1 (g28750), .I2 (g23952));
AN3X1 gate12887(.O (g25411), .I1 (g5062), .I2 (g23764), .I3 (I24546));
AN2X1 gate12888(.O (g26094), .I1 (g24936), .I2 (g9664));
AN2X1 gate12889(.O (g31765), .I1 (g30128), .I2 (g23968));
AN2X1 gate12890(.O (g24415), .I1 (g4760), .I2 (g22869));
AN2X1 gate12891(.O (g7763), .I1 (g2965), .I2 (g2960));
AN2X1 gate12892(.O (g24333), .I1 (g4512), .I2 (g22228));
AN2X1 gate12893(.O (g29369), .I1 (g28209), .I2 (g22341));
AN2X1 gate12894(.O (g14222), .I1 (g8655), .I2 (g11826));
AN2X1 gate12895(.O (g21922), .I1 (g5112), .I2 (g21468));
AN2X1 gate12896(.O (g22982), .I1 (g19535), .I2 (g19747));
AN2X1 gate12897(.O (g30111), .I1 (g28565), .I2 (g20917));
AN2X1 gate12898(.O (g18745), .I1 (g5128), .I2 (g17847));
AN2X1 gate12899(.O (g33690), .I1 (g33146), .I2 (g16280));
AN2X1 gate12900(.O (g30070), .I1 (g29167), .I2 (g9529));
AN2X1 gate12901(.O (g34111), .I1 (g33733), .I2 (g22936));
AN2X1 gate12902(.O (g18799), .I1 (g6181), .I2 (g15348));
AN2X1 gate12903(.O (g22091), .I1 (g6415), .I2 (g18833));
AN2X1 gate12904(.O (g23531), .I1 (g10760), .I2 (g18930));
AN2X1 gate12905(.O (g13853), .I1 (g4549), .I2 (g10620));
AN2X1 gate12906(.O (g18813), .I1 (g6513), .I2 (g15483));
AN2X1 gate12907(.O (g30590), .I1 (g18911), .I2 (g29812));
AN2X1 gate12908(.O (g21740), .I1 (g3085), .I2 (g20330));
AN2X1 gate12909(.O (g16599), .I1 (g6601), .I2 (g15030));
AN2X1 gate12910(.O (g26019), .I1 (g5507), .I2 (g25032));
AN2X1 gate12911(.O (g25503), .I1 (g6888), .I2 (g22529));
AN2X1 gate12912(.O (g18798), .I1 (g6177), .I2 (g15348));
AN2X1 gate12913(.O (g28542), .I1 (g27405), .I2 (g20275));
AN2X1 gate12914(.O (g31504), .I1 (g29370), .I2 (g10553));
AN2X1 gate12915(.O (g28453), .I1 (g27582), .I2 (g10233));
AN2X1 gate12916(.O (g27206), .I1 (g26055), .I2 (g16691));
AN3X1 gate12917(.O (g33504), .I1 (g32772), .I2 (I31216), .I3 (I31217));
AN2X1 gate12918(.O (g24664), .I1 (g22652), .I2 (g19741));
AN2X1 gate12919(.O (g29850), .I1 (g28340), .I2 (g24893));
AN2X1 gate12920(.O (g19911), .I1 (g14707), .I2 (g17748));
AN2X1 gate12921(.O (g34741), .I1 (g8899), .I2 (g34697));
AN2X1 gate12922(.O (g16598), .I1 (g6283), .I2 (g14899));
AN2X1 gate12923(.O (g15810), .I1 (g3937), .I2 (g14055));
AN2X1 gate12924(.O (g13524), .I1 (g9995), .I2 (g11910));
AN2X1 gate12925(.O (g17091), .I1 (g8659), .I2 (g12940));
AN2X1 gate12926(.O (g18184), .I1 (g785), .I2 (g17328));
AN2X1 gate12927(.O (g21953), .I1 (g5377), .I2 (g21514));
AN2X1 gate12928(.O (g18805), .I1 (g6377), .I2 (g15656));
AN2X1 gate12929(.O (g18674), .I1 (g4340), .I2 (g15758));
AN2X1 gate12930(.O (g23373), .I1 (g13699), .I2 (g20195));
AN2X1 gate12931(.O (g30094), .I1 (g28544), .I2 (g20767));
AN4X1 gate12932(.O (g27759), .I1 (g22457), .I2 (g25224), .I3 (g26424), .I4 (g26213));
AN2X1 gate12933(.O (g25581), .I1 (g19338), .I2 (g24150));
AN2X1 gate12934(.O (g25450), .I1 (g6888), .I2 (g22497));
AN2X1 gate12935(.O (g32042), .I1 (g27244), .I2 (g31070));
AN2X1 gate12936(.O (g21800), .I1 (g3546), .I2 (g20924));
AN2X1 gate12937(.O (g24484), .I1 (g16288), .I2 (g23208));
AN2X1 gate12938(.O (g29896), .I1 (g2599), .I2 (g29171));
AN2X1 gate12939(.O (g27114), .I1 (g25997), .I2 (g16523));
AN2X1 gate12940(.O (g32255), .I1 (g31248), .I2 (g20381));
AN2X1 gate12941(.O (g31129), .I1 (g1968), .I2 (g30017));
AN2X1 gate12942(.O (g32189), .I1 (g30824), .I2 (g25369));
AN2X1 gate12943(.O (g21936), .I1 (g5200), .I2 (g18997));
AN2X1 gate12944(.O (g18732), .I1 (g4961), .I2 (g16877));
AN2X1 gate12945(.O (g27435), .I1 (g26549), .I2 (g17585));
AN2X1 gate12946(.O (g18934), .I1 (g3133), .I2 (g16096));
AN2X1 gate12947(.O (g30735), .I1 (g29814), .I2 (g22319));
AN2X1 gate12948(.O (g24554), .I1 (g22490), .I2 (g19541));
AN2X1 gate12949(.O (g27107), .I1 (g26055), .I2 (g16514));
AN2X1 gate12950(.O (g32270), .I1 (g31254), .I2 (g20444));
AN2X1 gate12951(.O (g16125), .I1 (g5152), .I2 (g14238));
AN2X1 gate12952(.O (g16532), .I1 (g5252), .I2 (g14841));
AN2X1 gate12953(.O (g25818), .I1 (g8124), .I2 (g24605));
AN2X1 gate12954(.O (g28530), .I1 (g27383), .I2 (g20240));
AN2X1 gate12955(.O (g31128), .I1 (g12187), .I2 (g30016));
AN2X1 gate12956(.O (g32188), .I1 (g27586), .I2 (g31376));
AN2X1 gate12957(.O (g25979), .I1 (g24517), .I2 (g19650));
AN2X1 gate12958(.O (g28346), .I1 (g27243), .I2 (g19800));
AN2X1 gate12959(.O (g7251), .I1 (g452), .I2 (g392));
AN2X1 gate12960(.O (g24312), .I1 (g4501), .I2 (g22228));
AN2X1 gate12961(.O (g18692), .I1 (g4732), .I2 (g16053));
AN2X1 gate12962(.O (g18761), .I1 (g5471), .I2 (g17929));
AN2X1 gate12963(.O (g33245), .I1 (g32125), .I2 (g19961));
AN2X1 gate12964(.O (g24608), .I1 (g6500), .I2 (g23425));
AN2X1 gate12965(.O (g25978), .I1 (g9391), .I2 (g25001));
AN2X1 gate12966(.O (g13313), .I1 (g475), .I2 (g11048));
AN2X1 gate12967(.O (g15967), .I1 (g3913), .I2 (g14058));
AN2X1 gate12968(.O (g30196), .I1 (g28659), .I2 (g23858));
AN2X1 gate12969(.O (g31323), .I1 (g30150), .I2 (g27907));
AN2X1 gate12970(.O (g29582), .I1 (g27766), .I2 (g28608));
AN2X1 gate12971(.O (g31299), .I1 (g30123), .I2 (g27800));
AN2X1 gate12972(.O (g17192), .I1 (g1677), .I2 (g13022));
AN2X1 gate12973(.O (g34196), .I1 (g33682), .I2 (g24485));
AN2X1 gate12974(.O (g21762), .I1 (g3219), .I2 (g20785));
AN2X1 gate12975(.O (g21964), .I1 (g5441), .I2 (g21514));
AN2X1 gate12976(.O (g25986), .I1 (g5160), .I2 (g25013));
AN2X1 gate12977(.O (g32030), .I1 (g4172), .I2 (g30937));
AN2X1 gate12978(.O (g24921), .I1 (g23721), .I2 (g20739));
AN4X1 gate12979(.O (I31016), .I1 (g30825), .I2 (g31798), .I3 (g32478), .I4 (g32479));
AN2X1 gate12980(.O (g31298), .I1 (g30169), .I2 (g27886));
AN2X1 gate12981(.O (g34526), .I1 (g34300), .I2 (g19569));
AN2X1 gate12982(.O (g18400), .I1 (g2012), .I2 (g15373));
AN2X1 gate12983(.O (g10873), .I1 (g3004), .I2 (g9015));
AN2X1 gate12984(.O (g26077), .I1 (g9607), .I2 (g25233));
AN2X1 gate12985(.O (g24745), .I1 (g650), .I2 (g23550));
AN2X1 gate12986(.O (g29627), .I1 (g28493), .I2 (g11884));
AN2X1 gate12987(.O (g18214), .I1 (g939), .I2 (g15979));
AN2X1 gate12988(.O (g28292), .I1 (g23781), .I2 (g27762));
AN2X1 gate12989(.O (g29959), .I1 (g28953), .I2 (g12823));
AN2X1 gate12990(.O (g22862), .I1 (g1570), .I2 (g19673));
AN3X1 gate12991(.O (g28153), .I1 (g26424), .I2 (g22763), .I3 (g27031));
AN2X1 gate12992(.O (g18329), .I1 (g1612), .I2 (g17873));
AN2X1 gate12993(.O (g25067), .I1 (g4722), .I2 (g22885));
AN2X1 gate12994(.O (g25094), .I1 (g23318), .I2 (g20554));
AN2X1 gate12995(.O (g18207), .I1 (g925), .I2 (g15938));
AN2X1 gate12996(.O (g26689), .I1 (g15754), .I2 (g24431));
AN2X1 gate12997(.O (g29378), .I1 (g28137), .I2 (g22493));
AN2X1 gate12998(.O (g13808), .I1 (g4543), .I2 (g10607));
AN2X1 gate12999(.O (g18539), .I1 (g2763), .I2 (g15277));
AN2X1 gate13000(.O (g11036), .I1 (g9806), .I2 (g5774));
AN2X1 gate13001(.O (g26280), .I1 (g13051), .I2 (g25248));
AN2X1 gate13002(.O (g18328), .I1 (g1657), .I2 (g17873));
AN2X1 gate13003(.O (g27263), .I1 (g25940), .I2 (g19713));
AN2X1 gate13004(.O (g21909), .I1 (g5041), .I2 (g21468));
AN2X1 gate13005(.O (g31232), .I1 (g30294), .I2 (g23972));
AN2X1 gate13006(.O (g25150), .I1 (g17480), .I2 (g23547));
AN2X1 gate13007(.O (g22040), .I1 (g5953), .I2 (g19147));
AN2X1 gate13008(.O (g25801), .I1 (g8097), .I2 (g24585));
AN2X1 gate13009(.O (g26300), .I1 (g1968), .I2 (g25341));
AN2X1 gate13010(.O (g34866), .I1 (g34819), .I2 (g20106));
AN2X1 gate13011(.O (g28136), .I1 (g27382), .I2 (g23135));
AN2X1 gate13012(.O (g18538), .I1 (g2759), .I2 (g15277));
AN2X1 gate13013(.O (g15079), .I1 (g2151), .I2 (g12955));
AN2X1 gate13014(.O (g27332), .I1 (g12538), .I2 (g26758));
AN2X1 gate13015(.O (g29603), .I1 (g2265), .I2 (g29060));
AN2X1 gate13016(.O (g24674), .I1 (g446), .I2 (g23496));
AN2X1 gate13017(.O (g29742), .I1 (g28288), .I2 (g10233));
AN2X1 gate13018(.O (g21908), .I1 (g5037), .I2 (g21468));
AN2X1 gate13019(.O (g15078), .I1 (g10361), .I2 (g12955));
AN2X1 gate13020(.O (g33697), .I1 (g33160), .I2 (g13330));
AN2X1 gate13021(.O (g30001), .I1 (g28490), .I2 (g23486));
AN2X1 gate13022(.O (g31995), .I1 (g28274), .I2 (g30569));
AN2X1 gate13023(.O (g33856), .I1 (g33266), .I2 (g20442));
AN2X1 gate13024(.O (g26102), .I1 (g1825), .I2 (g25099));
AN2X1 gate13025(.O (g12135), .I1 (g9684), .I2 (g9959));
AN2X1 gate13026(.O (g31261), .I1 (g14754), .I2 (g30259));
AN2X1 gate13027(.O (g26157), .I1 (g2093), .I2 (g25136));
AN2X1 gate13028(.O (g27406), .I1 (g26488), .I2 (g17521));
AN3X1 gate13029(.O (g34077), .I1 (g22957), .I2 (g9104), .I3 (g33736));
AN2X1 gate13030(.O (g27962), .I1 (g25954), .I2 (g19597));
AN2X1 gate13031(.O (g27361), .I1 (g26519), .I2 (g17419));
AN2X1 gate13032(.O (g33880), .I1 (g33290), .I2 (g20568));
AN4X1 gate13033(.O (I31042), .I1 (g32515), .I2 (g32516), .I3 (g32517), .I4 (g32518));
AN2X1 gate13034(.O (g18241), .I1 (g1183), .I2 (g16431));
AN2X1 gate13035(.O (g34706), .I1 (g34496), .I2 (g10570));
AN2X1 gate13036(.O (g21747), .I1 (g3061), .I2 (g20330));
AN2X1 gate13037(.O (g32160), .I1 (g31001), .I2 (g22995));
AN2X1 gate13038(.O (g30256), .I1 (g28749), .I2 (g23947));
AN2X1 gate13039(.O (g25526), .I1 (g23720), .I2 (g21400));
AN2X1 gate13040(.O (g28164), .I1 (g8651), .I2 (g27528));
AN2X1 gate13041(.O (g26231), .I1 (g1854), .I2 (g25300));
AN3X1 gate13042(.O (g33512), .I1 (g32830), .I2 (I31256), .I3 (I31257));
AN2X1 gate13043(.O (g14913), .I1 (g1442), .I2 (g10939));
AN2X1 gate13044(.O (g27500), .I1 (g26400), .I2 (g17672));
AN2X1 gate13045(.O (g29857), .I1 (g28386), .I2 (g23304));
AN2X1 gate13046(.O (g15817), .I1 (g3921), .I2 (g13929));
AN2X1 gate13047(.O (g14614), .I1 (g11975), .I2 (g11997));
AN2X1 gate13048(.O (g24761), .I1 (g22751), .I2 (g19852));
AN2X1 gate13049(.O (g19540), .I1 (g1124), .I2 (g15904));
AN2X1 gate13050(.O (g21814), .I1 (g3594), .I2 (g20924));
AN2X1 gate13051(.O (g18771), .I1 (g5685), .I2 (g15615));
AN2X1 gate13052(.O (g16023), .I1 (g3813), .I2 (g13584));
AN2X1 gate13053(.O (g16224), .I1 (g14583), .I2 (g14232));
AN4X1 gate13054(.O (g11166), .I1 (g8363), .I2 (g269), .I3 (g8296), .I4 (I14225));
AN2X1 gate13055(.O (g18235), .I1 (g1141), .I2 (g16326));
AN2X1 gate13056(.O (g21751), .I1 (g3167), .I2 (g20785));
AN2X1 gate13057(.O (g21807), .I1 (g3566), .I2 (g20924));
AN2X1 gate13058(.O (g21772), .I1 (g3259), .I2 (g20785));
AN2X1 gate13059(.O (g26854), .I1 (g2868), .I2 (g24534));
AN2X1 gate13060(.O (g15783), .I1 (g3215), .I2 (g14098));
AN2X1 gate13061(.O (g21974), .I1 (g5517), .I2 (g19074));
AN2X1 gate13062(.O (g22062), .I1 (g6093), .I2 (g21611));
AN2X1 gate13063(.O (g18683), .I1 (g4674), .I2 (g15885));
AN2X1 gate13064(.O (g25866), .I1 (g3853), .I2 (g24648));
AN2X1 gate13065(.O (g24400), .I1 (g3466), .I2 (g23112));
AN2X1 gate13066(.O (g27221), .I1 (g26055), .I2 (g16747));
AN3X1 gate13067(.O (g33831), .I1 (g23088), .I2 (g33149), .I3 (g9104));
AN2X1 gate13068(.O (g28327), .I1 (g27365), .I2 (g19785));
AN2X1 gate13069(.O (g29549), .I1 (g2012), .I2 (g28900));
AN2X1 gate13070(.O (g34102), .I1 (g33912), .I2 (g23599));
AN2X1 gate13071(.O (g26511), .I1 (g19265), .I2 (g24364));
AN2X1 gate13072(.O (g34157), .I1 (g33794), .I2 (g20159));
AN2X1 gate13073(.O (g23639), .I1 (g19050), .I2 (g9104));
AN4X1 gate13074(.O (I31267), .I1 (g32840), .I2 (g32841), .I3 (g32842), .I4 (g32843));
AN2X1 gate13075(.O (g10565), .I1 (g8182), .I2 (g424));
AN2X1 gate13076(.O (g28537), .I1 (g6832), .I2 (g27089));
AN2X1 gate13077(.O (g31499), .I1 (g29801), .I2 (g23446));
AN3X1 gate13078(.O (g33499), .I1 (g32737), .I2 (I31191), .I3 (I31192));
AN2X1 gate13079(.O (g14565), .I1 (g11934), .I2 (g11952));
AN2X1 gate13080(.O (g29548), .I1 (g1798), .I2 (g28575));
AN2X1 gate13081(.O (g23293), .I1 (g9104), .I2 (g19200));
AN2X1 gate13082(.O (g24329), .I1 (g4462), .I2 (g22228));
AN2X1 gate13083(.O (g30066), .I1 (g28518), .I2 (g20636));
AN2X1 gate13084(.O (g22851), .I1 (g496), .I2 (g19654));
AN2X1 gate13085(.O (g28108), .I1 (g7975), .I2 (g27237));
AN2X1 gate13086(.O (g30231), .I1 (g28718), .I2 (g23907));
AN2X1 gate13087(.O (g15823), .I1 (g3945), .I2 (g14116));
AN2X1 gate13088(.O (g34066), .I1 (g33730), .I2 (g19352));
AN2X1 gate13089(.O (g10034), .I1 (g1521), .I2 (g1500));
AN2X1 gate13090(.O (g25077), .I1 (g23297), .I2 (g20536));
AN3X1 gate13091(.O (g33498), .I1 (g32730), .I2 (I31186), .I3 (I31187));
AN2X1 gate13092(.O (g23265), .I1 (g20069), .I2 (g20132));
AN2X1 gate13093(.O (g24328), .I1 (g4567), .I2 (g22228));
AN3X1 gate13094(.O (g28283), .I1 (g7380), .I2 (g2361), .I3 (g27445));
AN2X1 gate13095(.O (g18515), .I1 (g2643), .I2 (g15509));
AN2X1 gate13096(.O (g23416), .I1 (g20082), .I2 (g20321));
AN2X1 gate13097(.O (g18414), .I1 (g2102), .I2 (g15373));
AN2X1 gate13098(.O (g31989), .I1 (g31770), .I2 (g22200));
AN2X1 gate13099(.O (g14641), .I1 (g11994), .I2 (g12020));
AN3X1 gate13100(.O (g28303), .I1 (g7462), .I2 (g2629), .I3 (g27494));
AN2X1 gate13101(.O (g27106), .I1 (g26026), .I2 (g16512));
AN2X1 gate13102(.O (g21841), .I1 (g3857), .I2 (g21070));
AN2X1 gate13103(.O (g21992), .I1 (g5599), .I2 (g19074));
AN2X1 gate13104(.O (g34876), .I1 (g34844), .I2 (g20534));
AN2X1 gate13105(.O (g18407), .I1 (g2016), .I2 (g15373));
AN2X1 gate13106(.O (g25923), .I1 (g24443), .I2 (g19443));
AN2X1 gate13107(.O (g31988), .I1 (g31768), .I2 (g22199));
AN2X1 gate13108(.O (g33722), .I1 (g33175), .I2 (g19445));
AN2X1 gate13109(.O (g33924), .I1 (g33335), .I2 (g33346));
AN2X1 gate13110(.O (g32419), .I1 (g4955), .I2 (g31000));
AN2X1 gate13111(.O (g15966), .I1 (g3462), .I2 (g13555));
AN4X1 gate13112(.O (g28982), .I1 (g27163), .I2 (g12687), .I3 (g20682), .I4 (I27349));
AN2X1 gate13113(.O (g31271), .I1 (g29706), .I2 (g23300));
AN2X1 gate13114(.O (g12812), .I1 (g518), .I2 (g9158));
AN2X1 gate13115(.O (g34763), .I1 (g34689), .I2 (g19915));
AN2X1 gate13116(.O (g15631), .I1 (g168), .I2 (g13437));
AN2X1 gate13117(.O (g27033), .I1 (g25767), .I2 (g19273));
AN2X1 gate13118(.O (g27371), .I1 (g26400), .I2 (g17473));
AN2X1 gate13119(.O (g32418), .I1 (g31126), .I2 (g16239));
AN2X1 gate13120(.O (g26287), .I1 (g2138), .I2 (g25225));
AN2X1 gate13121(.O (g27234), .I1 (g26055), .I2 (g16814));
AN2X1 gate13122(.O (g25102), .I1 (g4727), .I2 (g22885));
AN2X1 gate13123(.O (g21835), .I1 (g3802), .I2 (g20453));
AN2X1 gate13124(.O (g32170), .I1 (g31671), .I2 (g27779));
AN2X1 gate13125(.O (g13567), .I1 (g10102), .I2 (g11948));
AN2X1 gate13126(.O (g22047), .I1 (g6077), .I2 (g21611));
AN2X1 gate13127(.O (g26307), .I1 (g13070), .I2 (g25288));
AN2X1 gate13128(.O (g26085), .I1 (g11906), .I2 (g25070));
AN2X1 gate13129(.O (g29626), .I1 (g28584), .I2 (g11415));
AN3X1 gate13130(.O (g33461), .I1 (g32463), .I2 (I31001), .I3 (I31002));
AN2X1 gate13131(.O (g16669), .I1 (g5611), .I2 (g14993));
AN2X1 gate13132(.O (g33342), .I1 (g32226), .I2 (g20660));
AN3X1 gate13133(.O (g29323), .I1 (g28539), .I2 (g6905), .I3 (g3639));
AN2X1 gate13134(.O (g23007), .I1 (g681), .I2 (g20248));
AN2X1 gate13135(.O (g31145), .I1 (g9970), .I2 (g30052));
AN2X1 gate13136(.O (g18441), .I1 (g2246), .I2 (g18008));
AN2X1 gate13137(.O (g18584), .I1 (g2950), .I2 (g16349));
AN2X1 gate13138(.O (g24771), .I1 (g7028), .I2 (g23605));
AN2X1 gate13139(.O (g18206), .I1 (g918), .I2 (g15938));
AN2X1 gate13140(.O (g29533), .I1 (g28958), .I2 (g22417));
AN2X1 gate13141(.O (g12795), .I1 (g1312), .I2 (g7601));
AN2X1 gate13142(.O (g16668), .I1 (g5543), .I2 (g14962));
AN2X1 gate13143(.O (g16842), .I1 (g6279), .I2 (g14861));
AN2X1 gate13144(.O (g17574), .I1 (g9554), .I2 (g14546));
AN2X1 gate13145(.O (g33887), .I1 (g33298), .I2 (g20615));
AN2X1 gate13146(.O (g18759), .I1 (g5467), .I2 (g17929));
AN2X1 gate13147(.O (g22051), .I1 (g6105), .I2 (g21611));
AN2X1 gate13148(.O (g22072), .I1 (g6259), .I2 (g19210));
AN2X1 gate13149(.O (g18725), .I1 (g4912), .I2 (g16077));
AN2X1 gate13150(.O (g32167), .I1 (g3853), .I2 (g31194));
AN2X1 gate13151(.O (g32194), .I1 (g30601), .I2 (g28436));
AN2X1 gate13152(.O (g25876), .I1 (g3470), .I2 (g24667));
AN3X1 gate13153(.O (g33529), .I1 (g32953), .I2 (I31341), .I3 (I31342));
AN4X1 gate13154(.O (I31201), .I1 (g31672), .I2 (g31831), .I3 (g32745), .I4 (g32746));
AN2X1 gate13155(.O (g27507), .I1 (g26549), .I2 (g17683));
AN4X1 gate13156(.O (I31277), .I1 (g32856), .I2 (g32857), .I3 (g32858), .I4 (g32859));
AN2X1 gate13157(.O (g18114), .I1 (g452), .I2 (g17015));
AN2X1 gate13158(.O (g28192), .I1 (g8891), .I2 (g27415));
AN2X1 gate13159(.O (g18758), .I1 (g7004), .I2 (g15595));
AN2X1 gate13160(.O (g31528), .I1 (g19050), .I2 (g29814));
AN2X1 gate13161(.O (g26341), .I1 (g24746), .I2 (g20105));
AN2X1 gate13162(.O (g18435), .I1 (g2173), .I2 (g18008));
AN3X1 gate13163(.O (g33528), .I1 (g32946), .I2 (I31336), .I3 (I31337));
AN2X1 gate13164(.O (g34287), .I1 (g11370), .I2 (g34124));
AN2X1 gate13165(.O (g19661), .I1 (g5489), .I2 (g16969));
AN2X1 gate13166(.O (g33843), .I1 (g33256), .I2 (g20325));
AN2X1 gate13167(.O (g21720), .I1 (g376), .I2 (g21037));
AN2X1 gate13168(.O (g33330), .I1 (g32211), .I2 (g20588));
AN2X1 gate13169(.O (g26156), .I1 (g2028), .I2 (g25135));
AN2X1 gate13170(.O (g18107), .I1 (g429), .I2 (g17015));
AN4X1 gate13171(.O (g27421), .I1 (g8038), .I2 (g26314), .I3 (g9187), .I4 (g9077));
AN3X1 gate13172(.O (g34085), .I1 (g33761), .I2 (g9104), .I3 (g18957));
AN2X1 gate13173(.O (g28663), .I1 (g27566), .I2 (g20624));
AN2X1 gate13174(.O (g32401), .I1 (g31116), .I2 (g13432));
AN2X1 gate13175(.O (g34076), .I1 (g33694), .I2 (g19519));
AN2X1 gate13176(.O (g30596), .I1 (g30279), .I2 (g18947));
AN2X1 gate13177(.O (g26180), .I1 (g2587), .I2 (g25156));
AN2X1 gate13178(.O (g26670), .I1 (g13385), .I2 (g24428));
AN2X1 gate13179(.O (g21746), .I1 (g3045), .I2 (g20330));
AN2X1 gate13180(.O (g33365), .I1 (g32267), .I2 (g20994));
AN2X1 gate13181(.O (g32119), .I1 (g31609), .I2 (g29939));
AN2X1 gate13182(.O (g30243), .I1 (g28731), .I2 (g23929));
AN2X1 gate13183(.O (g31132), .I1 (g29504), .I2 (g22987));
AN2X1 gate13184(.O (g18744), .I1 (g5124), .I2 (g17847));
AN2X1 gate13185(.O (g34054), .I1 (g33778), .I2 (g22942));
AN2X1 gate13186(.O (g31960), .I1 (g31749), .I2 (g22153));
AN2X1 gate13187(.O (g33869), .I1 (g33279), .I2 (g20543));
AN2X1 gate13188(.O (g14537), .I1 (g10550), .I2 (g10529));
AN2X1 gate13189(.O (g18345), .I1 (g1736), .I2 (g17955));
AN2X1 gate13190(.O (g19715), .I1 (g9679), .I2 (g17120));
AN4X1 gate13191(.O (I31037), .I1 (g32508), .I2 (g32509), .I3 (g32510), .I4 (g32511));
AN2X1 gate13192(.O (g29856), .I1 (g28385), .I2 (g23303));
AN4X1 gate13193(.O (g17780), .I1 (g6772), .I2 (g11592), .I3 (g11640), .I4 (I18782));
AN2X1 gate13194(.O (g21465), .I1 (g16155), .I2 (g13663));
AN2X1 gate13195(.O (g18399), .I1 (g2024), .I2 (g15373));
AN2X1 gate13196(.O (g29880), .I1 (g1936), .I2 (g29149));
AN2X1 gate13197(.O (g33868), .I1 (g33278), .I2 (g20542));
AN2X1 gate13198(.O (g26839), .I1 (g2988), .I2 (g24516));
AN2X1 gate13199(.O (g27541), .I1 (g26278), .I2 (g23334));
AN2X1 gate13200(.O (g30269), .I1 (g28778), .I2 (g23970));
AN2X1 gate13201(.O (g22846), .I1 (g9386), .I2 (g20676));
AN2X1 gate13202(.O (g21983), .I1 (g5555), .I2 (g19074));
AN2X1 gate13203(.O (g28553), .I1 (g27187), .I2 (g10290));
AN3X1 gate13204(.O (g25456), .I1 (g5752), .I2 (g22210), .I3 (I24579));
AN2X1 gate13205(.O (g18398), .I1 (g2020), .I2 (g15373));
AN2X1 gate13206(.O (g29512), .I1 (g2161), .I2 (g28793));
AN2X1 gate13207(.O (g32313), .I1 (g31303), .I2 (g23515));
AN4X1 gate13208(.O (I31352), .I1 (g32963), .I2 (g32964), .I3 (g32965), .I4 (g32966));
AN2X1 gate13209(.O (g21806), .I1 (g3558), .I2 (g20924));
AN2X1 gate13210(.O (g26838), .I1 (g2860), .I2 (g24515));
AN2X1 gate13211(.O (g18141), .I1 (g568), .I2 (g17533));
AN2X1 gate13212(.O (g30268), .I1 (g28777), .I2 (g23969));
AN2X1 gate13213(.O (g18652), .I1 (g4172), .I2 (g16249));
AN2X1 gate13214(.O (g18804), .I1 (g15163), .I2 (g15656));
AN2X1 gate13215(.O (g34341), .I1 (g34101), .I2 (g19952));
AN2X1 gate13216(.O (g25916), .I1 (g24432), .I2 (g19434));
AN2X1 gate13217(.O (g16610), .I1 (g5260), .I2 (g14918));
AN2X1 gate13218(.O (g16705), .I1 (g6299), .I2 (g15024));
AN2X1 gate13219(.O (g17152), .I1 (g8635), .I2 (g12997));
AN2X1 gate13220(.O (g31225), .I1 (g30276), .I2 (g21012));
AN2X1 gate13221(.O (g32276), .I1 (g31646), .I2 (g30313));
AN4X1 gate13222(.O (g27724), .I1 (g22417), .I2 (g25208), .I3 (g26424), .I4 (g26190));
AN2X1 gate13223(.O (g34655), .I1 (g34573), .I2 (g18885));
AN4X1 gate13224(.O (I31266), .I1 (g31327), .I2 (g31843), .I3 (g32838), .I4 (g32839));
AN2X1 gate13225(.O (g27359), .I1 (g26488), .I2 (g17416));
AN2X1 gate13226(.O (g30180), .I1 (g28635), .I2 (g23820));
AN2X1 gate13227(.O (g27325), .I1 (g12478), .I2 (g26724));
AN2X1 gate13228(.O (g30670), .I1 (g11330), .I2 (g29359));
AN2X1 gate13229(.O (g31471), .I1 (g29754), .I2 (g23399));
AN2X1 gate13230(.O (g32305), .I1 (g31287), .I2 (g20567));
AN2X1 gate13231(.O (g32053), .I1 (g14176), .I2 (g31509));
AN3X1 gate13232(.O (g33471), .I1 (g32535), .I2 (I31051), .I3 (I31052));
AN2X1 gate13233(.O (g34180), .I1 (g33716), .I2 (g24373));
AN2X1 gate13234(.O (g33087), .I1 (g32391), .I2 (g18888));
AN2X1 gate13235(.O (g18263), .I1 (g1249), .I2 (g16000));
AN2X1 gate13236(.O (g32254), .I1 (g31247), .I2 (g20379));
AN2X1 gate13237(.O (g27535), .I1 (g26519), .I2 (g17737));
AN2X1 gate13238(.O (g26487), .I1 (g15702), .I2 (g24359));
AN2X1 gate13239(.O (g27434), .I1 (g26549), .I2 (g17584));
AN2X1 gate13240(.O (g27358), .I1 (g26400), .I2 (g17415));
AN2X1 gate13241(.O (g25076), .I1 (g12805), .I2 (g23479));
AN2X1 gate13242(.O (g25085), .I1 (g4912), .I2 (g22908));
AN2X1 gate13243(.O (g18332), .I1 (g1677), .I2 (g17873));
AN2X1 gate13244(.O (g19784), .I1 (g2775), .I2 (g15877));
AN2X1 gate13245(.O (g28252), .I1 (g27159), .I2 (g19682));
AN2X1 gate13246(.O (g12920), .I1 (g1227), .I2 (g10960));
AN2X1 gate13247(.O (g18135), .I1 (g136), .I2 (g17249));
AN2X1 gate13248(.O (g34335), .I1 (g8461), .I2 (g34197));
AN2X1 gate13249(.O (g25054), .I1 (g12778), .I2 (g23452));
AN2X1 gate13250(.O (g24725), .I1 (g19587), .I2 (g23012));
AN2X1 gate13251(.O (g30930), .I1 (g29915), .I2 (g23342));
AN2X1 gate13252(.O (g32036), .I1 (g31469), .I2 (g13486));
AN2X1 gate13253(.O (g27121), .I1 (g136), .I2 (g26326));
AN3X1 gate13254(.O (g29316), .I1 (g28528), .I2 (g6875), .I3 (g3288));
AN2X1 gate13255(.O (g19354), .I1 (g471), .I2 (g16235));
AN2X1 gate13256(.O (g33244), .I1 (g32190), .I2 (g23152));
AN2X1 gate13257(.O (g32177), .I1 (g30608), .I2 (g25214));
AN2X1 gate13258(.O (g18406), .I1 (g2060), .I2 (g15373));
AN2X1 gate13259(.O (g13349), .I1 (g4933), .I2 (g11780));
AN4X1 gate13260(.O (I31167), .I1 (g32696), .I2 (g32697), .I3 (g32698), .I4 (g32699));
AN3X1 gate13261(.O (I18785), .I1 (g13156), .I2 (g6767), .I3 (g11498));
AN2X1 gate13262(.O (g26279), .I1 (g4249), .I2 (g25213));
AN2X1 gate13263(.O (g18361), .I1 (g1821), .I2 (g17955));
AN2X1 gate13264(.O (g24758), .I1 (g6523), .I2 (g23733));
AN2X1 gate13265(.O (g23130), .I1 (g728), .I2 (g20248));
AN2X1 gate13266(.O (g34667), .I1 (g34471), .I2 (g33424));
AN2X1 gate13267(.O (g34694), .I1 (g34530), .I2 (g19885));
AN2X1 gate13268(.O (g17405), .I1 (g1422), .I2 (g13137));
AN2X1 gate13269(.O (g11083), .I1 (g8836), .I2 (g802));
AN2X1 gate13270(.O (g34965), .I1 (g34949), .I2 (g23084));
AN2X1 gate13271(.O (g30131), .I1 (g28589), .I2 (g21178));
AN2X1 gate13272(.O (g31069), .I1 (g29793), .I2 (g14150));
AN2X1 gate13273(.O (g19671), .I1 (g1454), .I2 (g16155));
AN2X1 gate13274(.O (g29989), .I1 (g29006), .I2 (g10489));
AN2X1 gate13275(.O (g18500), .I1 (g2421), .I2 (g15426));
AN2X1 gate13276(.O (g22020), .I1 (g5863), .I2 (g19147));
AN2X1 gate13277(.O (g27682), .I1 (g25777), .I2 (g23565));
AN2X1 gate13278(.O (g23165), .I1 (g13954), .I2 (g19964));
AN2X1 gate13279(.O (g28183), .I1 (g27024), .I2 (g19421));
AN2X1 gate13280(.O (g28673), .I1 (g1373), .I2 (g27122));
AN2X1 gate13281(.O (g33810), .I1 (g33427), .I2 (g12768));
AN2X1 gate13282(.O (g27291), .I1 (g11969), .I2 (g26653));
AN2X1 gate13283(.O (g29611), .I1 (g28540), .I2 (g14209));
AN2X1 gate13284(.O (g33657), .I1 (g30991), .I2 (g33443));
AN2X1 gate13285(.O (g26286), .I1 (g2126), .I2 (g25389));
AN2X1 gate13286(.O (g29988), .I1 (g29187), .I2 (g12235));
AN2X1 gate13287(.O (g29924), .I1 (g13031), .I2 (g29190));
AN2X1 gate13288(.O (g34487), .I1 (g34416), .I2 (g18983));
AN2X1 gate13289(.O (g13566), .I1 (g7092), .I2 (g12358));
AN2X1 gate13290(.O (g22046), .I1 (g6073), .I2 (g21611));
AN2X1 gate13291(.O (g26306), .I1 (g13087), .I2 (g25286));
AN2X1 gate13292(.O (g24849), .I1 (g4165), .I2 (g22227));
AN2X1 gate13293(.O (g33879), .I1 (g33289), .I2 (g20566));
AN2X1 gate13294(.O (g24940), .I1 (g5011), .I2 (g23971));
AN2X1 gate13295(.O (g24399), .I1 (g3133), .I2 (g23067));
AN2X1 gate13296(.O (g34502), .I1 (g26363), .I2 (g34343));
AN2X1 gate13297(.O (g30210), .I1 (g28684), .I2 (g23877));
AN2X1 gate13298(.O (g34557), .I1 (g34352), .I2 (g20555));
AN2X1 gate13299(.O (g23006), .I1 (g19575), .I2 (g19776));
AN2X1 gate13300(.O (g23475), .I1 (g19070), .I2 (g8971));
AN2X1 gate13301(.O (g33878), .I1 (g33288), .I2 (g20565));
AN4X1 gate13302(.O (I31022), .I1 (g32487), .I2 (g32488), .I3 (g32489), .I4 (g32490));
AN2X1 gate13303(.O (g18221), .I1 (g1018), .I2 (g16100));
AN2X1 gate13304(.O (g22113), .I1 (g6561), .I2 (g19277));
AN2X1 gate13305(.O (g21863), .I1 (g3957), .I2 (g21070));
AN2X1 gate13306(.O (g26815), .I1 (g4108), .I2 (g24528));
AN2X1 gate13307(.O (g24141), .I1 (g17657), .I2 (g21656));
AN2X1 gate13308(.O (g34279), .I1 (g34231), .I2 (g19208));
AN4X1 gate13309(.O (g11139), .I1 (g5990), .I2 (g7051), .I3 (g5976), .I4 (g9935));
AN2X1 gate13310(.O (g33886), .I1 (g33297), .I2 (g20614));
AN2X1 gate13311(.O (g27134), .I1 (g25997), .I2 (g16602));
AN2X1 gate13312(.O (g30278), .I1 (g28818), .I2 (g23988));
AN2X1 gate13313(.O (g27029), .I1 (g26327), .I2 (g11031));
AN2X1 gate13314(.O (g18613), .I1 (g3338), .I2 (g17200));
AN2X1 gate13315(.O (g31792), .I1 (g30214), .I2 (g24017));
AN2X1 gate13316(.O (g32166), .I1 (g31007), .I2 (g23029));
AN2X1 gate13317(.O (g32009), .I1 (g31782), .I2 (g22224));
AN2X1 gate13318(.O (g25993), .I1 (g2610), .I2 (g25025));
AN2X1 gate13319(.O (g31967), .I1 (g31755), .I2 (g22167));
AN2X1 gate13320(.O (g31994), .I1 (g31775), .I2 (g22215));
AN2X1 gate13321(.O (g22105), .I1 (g6494), .I2 (g18833));
AN4X1 gate13322(.O (I31276), .I1 (g31376), .I2 (g31844), .I3 (g32854), .I4 (g32855));
AN2X1 gate13323(.O (g27028), .I1 (g26342), .I2 (g1157));
AN2X1 gate13324(.O (g29199), .I1 (g27187), .I2 (g12687));
AN2X1 gate13325(.O (g32008), .I1 (g31781), .I2 (g22223));
AN2X1 gate13326(.O (g25965), .I1 (g2208), .I2 (g24980));
AN2X1 gate13327(.O (g29650), .I1 (g28949), .I2 (g22472));
AN2X1 gate13328(.O (g29736), .I1 (g28522), .I2 (g10233));
AN2X1 gate13329(.O (g16160), .I1 (g5499), .I2 (g14262));
AN2X1 gate13330(.O (g29887), .I1 (g28417), .I2 (g23351));
AN2X1 gate13331(.O (g21703), .I1 (g146), .I2 (g20283));
AN2X1 gate13332(.O (g18273), .I1 (g1287), .I2 (g16031));
AN2X1 gate13333(.O (g24332), .I1 (g4459), .I2 (g22228));
AN2X1 gate13334(.O (g18106), .I1 (g411), .I2 (g17015));
AN2X1 gate13335(.O (g20135), .I1 (g16258), .I2 (g16695));
AN2X1 gate13336(.O (g18605), .I1 (g3129), .I2 (g16987));
AN2X1 gate13337(.O (g13415), .I1 (g837), .I2 (g11048));
AN2X1 gate13338(.O (g21347), .I1 (g1339), .I2 (g15750));
AN2X1 gate13339(.O (g13333), .I1 (g4743), .I2 (g11755));
AN2X1 gate13340(.O (g33425), .I1 (g32380), .I2 (g21466));
AN2X1 gate13341(.O (g28213), .I1 (g27720), .I2 (g23380));
AN2X1 gate13342(.O (g15679), .I1 (g3470), .I2 (g13555));
AN2X1 gate13343(.O (g18812), .I1 (g6509), .I2 (g15483));
AN2X1 gate13344(.O (g10948), .I1 (g7880), .I2 (g1478));
AN2X1 gate13345(.O (g18463), .I1 (g2375), .I2 (g15224));
AN2X1 gate13346(.O (g33919), .I1 (g33438), .I2 (g10795));
AN2X1 gate13347(.O (g24406), .I1 (g13623), .I2 (g22860));
AN2X1 gate13348(.O (g29528), .I1 (g2429), .I2 (g28874));
AN4X1 gate13349(.O (I31036), .I1 (g30673), .I2 (g31802), .I3 (g32506), .I4 (g32507));
AN2X1 gate13350(.O (g24962), .I1 (g23194), .I2 (g20210));
AN2X1 gate13351(.O (g29843), .I1 (g28373), .I2 (g23289));
AN2X1 gate13352(.O (g21781), .I1 (g3408), .I2 (g20391));
AN2X1 gate13353(.O (g29330), .I1 (g29114), .I2 (g18894));
AN2X1 gate13354(.O (g16617), .I1 (g6287), .I2 (g14940));
AN2X1 gate13355(.O (g25502), .I1 (g6946), .I2 (g22527));
AN2X1 gate13356(.O (g15678), .I1 (g1094), .I2 (g13846));
AN4X1 gate13357(.O (I31101), .I1 (g30735), .I2 (g31813), .I3 (g32601), .I4 (g32602));
AN4X1 gate13358(.O (I31177), .I1 (g32710), .I2 (g32711), .I3 (g32712), .I4 (g32713));
AN2X1 gate13359(.O (g18951), .I1 (g3484), .I2 (g16124));
AN2X1 gate13360(.O (g30187), .I1 (g28643), .I2 (g23840));
AN2X1 gate13361(.O (g18371), .I1 (g1870), .I2 (g15171));
AN3X1 gate13362(.O (g8721), .I1 (g385), .I2 (g376), .I3 (g365));
AN2X1 gate13363(.O (g28205), .I1 (g27516), .I2 (g16746));
AN2X1 gate13364(.O (g18234), .I1 (g1129), .I2 (g16326));
AN2X1 gate13365(.O (g34187), .I1 (g33708), .I2 (g24397));
AN2X1 gate13366(.O (g17769), .I1 (g1146), .I2 (g13188));
AN2X1 gate13367(.O (g21952), .I1 (g5366), .I2 (g21514));
AN2X1 gate13368(.O (g28311), .I1 (g9792), .I2 (g27679));
AN2X1 gate13369(.O (g23372), .I1 (g16448), .I2 (g20194));
AN2X1 gate13370(.O (g29869), .I1 (g2331), .I2 (g29129));
AN2X1 gate13371(.O (g21821), .I1 (g3723), .I2 (g20453));
AN2X1 gate13372(.O (g17768), .I1 (g13325), .I2 (g10741));
AN4X1 gate13373(.O (I26530), .I1 (g26365), .I2 (g24096), .I3 (g24097), .I4 (g24098));
AN2X1 gate13374(.O (g18795), .I1 (g6163), .I2 (g15348));
AN2X1 gate13375(.O (g30937), .I1 (g22626), .I2 (g29814));
AN2X1 gate13376(.O (g29868), .I1 (g2227), .I2 (g29128));
AN2X1 gate13377(.O (g27649), .I1 (g10820), .I2 (g25820));
AN2X1 gate13378(.O (g34143), .I1 (g33934), .I2 (g23828));
AN2X1 gate13379(.O (g16595), .I1 (g5921), .I2 (g14697));
AN2X1 gate13380(.O (g21790), .I1 (g3454), .I2 (g20391));
AN2X1 gate13381(.O (g24004), .I1 (g37), .I2 (g21225));
AN2X1 gate13382(.O (g33086), .I1 (g32390), .I2 (g18887));
AN2X1 gate13383(.O (g27648), .I1 (g25882), .I2 (g8974));
AN2X1 gate13384(.O (g24221), .I1 (g232), .I2 (g22594));
AN2X1 gate13385(.O (g27491), .I1 (g26576), .I2 (g17652));
AN2X1 gate13386(.O (g26486), .I1 (g4423), .I2 (g24358));
AN2X1 gate13387(.O (g18514), .I1 (g2629), .I2 (g15509));
AN2X1 gate13388(.O (g29709), .I1 (g2116), .I2 (g29121));
AN2X1 gate13389(.O (g34169), .I1 (g33804), .I2 (g31227));
AN2X1 gate13390(.O (g21873), .I1 (g6946), .I2 (g19801));
AN2X1 gate13391(.O (g18507), .I1 (g2595), .I2 (g15509));
AN2X1 gate13392(.O (g22027), .I1 (g5889), .I2 (g19147));
AN2X1 gate13393(.O (g23873), .I1 (g21222), .I2 (g10815));
AN2X1 gate13394(.O (g15875), .I1 (g3961), .I2 (g13963));
AN2X1 gate13395(.O (g30168), .I1 (g28623), .I2 (g23794));
AN2X1 gate13396(.O (g29708), .I1 (g1955), .I2 (g29082));
AN2X1 gate13397(.O (g33817), .I1 (g33235), .I2 (g20102));
AN2X1 gate13398(.O (g11115), .I1 (g6133), .I2 (g9954));
AN2X1 gate13399(.O (g33322), .I1 (g32202), .I2 (g20450));
AN2X1 gate13400(.O (g34410), .I1 (g34204), .I2 (g21427));
AN2X1 gate13401(.O (g27981), .I1 (g26751), .I2 (g23924));
AN2X1 gate13402(.O (g25815), .I1 (g8155), .I2 (g24603));
AN2X1 gate13403(.O (g31125), .I1 (g29502), .I2 (g22973));
AN2X1 gate13404(.O (g32176), .I1 (g2779), .I2 (g31623));
AN4X1 gate13405(.O (I31166), .I1 (g30673), .I2 (g31825), .I3 (g32694), .I4 (g32695));
AN4X1 gate13406(.O (g26223), .I1 (g24688), .I2 (g10678), .I3 (g10658), .I4 (g8757));
AN2X1 gate13407(.O (g31977), .I1 (g31764), .I2 (g22179));
AN3X1 gate13408(.O (g33532), .I1 (g32974), .I2 (I31356), .I3 (I31357));
AN2X1 gate13409(.O (g33901), .I1 (g33317), .I2 (g20920));
AN2X1 gate13410(.O (g34479), .I1 (g34403), .I2 (g18905));
AN2X1 gate13411(.O (g34666), .I1 (g34587), .I2 (g19144));
AN2X1 gate13412(.O (g25187), .I1 (g12296), .I2 (g23629));
AN2X1 gate13413(.O (g18163), .I1 (g79), .I2 (g17433));
AN2X1 gate13414(.O (g15837), .I1 (g3255), .I2 (g14127));
AN2X1 gate13415(.O (g32154), .I1 (g31277), .I2 (g14184));
AN2X1 gate13416(.O (g34363), .I1 (g34148), .I2 (g20389));
AN2X1 gate13417(.O (g25975), .I1 (g9434), .I2 (g24999));
AN2X1 gate13418(.O (g34217), .I1 (g33736), .I2 (g22876));
AN2X1 gate13419(.O (g22710), .I1 (g19358), .I2 (g19600));
AN2X1 gate13420(.O (g30015), .I1 (g29040), .I2 (g10519));
AN2X1 gate13421(.O (g21834), .I1 (g3752), .I2 (g20453));
AN2X1 gate13422(.O (g22003), .I1 (g5736), .I2 (g21562));
AN2X1 gate13423(.O (g34478), .I1 (g34402), .I2 (g18904));
AN2X1 gate13424(.O (g28152), .I1 (g26297), .I2 (g27279));
AN2X1 gate13425(.O (g26084), .I1 (g24926), .I2 (g9602));
AN4X1 gate13426(.O (g28846), .I1 (g21434), .I2 (g26424), .I3 (g25399), .I4 (g27474));
AN2X1 gate13427(.O (g24812), .I1 (g19662), .I2 (g22192));
AN2X1 gate13428(.O (g19855), .I1 (g2787), .I2 (g15962));
AN2X1 gate13429(.O (g33353), .I1 (g32240), .I2 (g20732));
AN2X1 gate13430(.O (g25143), .I1 (g4922), .I2 (g22908));
AN2X1 gate13431(.O (g34486), .I1 (g34412), .I2 (g18953));
AN2X1 gate13432(.O (g18541), .I1 (g2767), .I2 (g15277));
AN4X1 gate13433(.O (g27395), .I1 (g8046), .I2 (g26314), .I3 (g9187), .I4 (g9077));
AN2X1 gate13434(.O (g33680), .I1 (g33128), .I2 (g4688));
AN2X1 gate13435(.O (g18473), .I1 (g2342), .I2 (g15224));
AN2X1 gate13436(.O (g27262), .I1 (g25997), .I2 (g17092));
AN2X1 gate13437(.O (g26179), .I1 (g2504), .I2 (g25155));
AN2X1 gate13438(.O (g12794), .I1 (g1008), .I2 (g7567));
AN3X1 gate13439(.O (I17529), .I1 (g13156), .I2 (g11450), .I3 (g6756));
AN2X1 gate13440(.O (g34556), .I1 (g34350), .I2 (g20537));
AN2X1 gate13441(.O (g18789), .I1 (g6035), .I2 (g15634));
AN2X1 gate13442(.O (g21453), .I1 (g16713), .I2 (g13625));
AN2X1 gate13443(.O (g22081), .I1 (g6279), .I2 (g19210));
AN2X1 gate13444(.O (g29602), .I1 (g2020), .I2 (g28962));
AN2X1 gate13445(.O (g29810), .I1 (g28259), .I2 (g11317));
AN2X1 gate13446(.O (g29774), .I1 (g28287), .I2 (g10233));
AN2X1 gate13447(.O (g34580), .I1 (g29539), .I2 (g34311));
AN2X1 gate13448(.O (g26178), .I1 (g2389), .I2 (g25473));
AN4X1 gate13449(.O (g16194), .I1 (g11547), .I2 (g6782), .I3 (g11640), .I4 (I17529));
AN2X1 gate13450(.O (g27633), .I1 (g13076), .I2 (g25766));
AN2X1 gate13451(.O (g21913), .I1 (g5069), .I2 (g21468));
AN2X1 gate13452(.O (g29375), .I1 (g13946), .I2 (g28370));
AN2X1 gate13453(.O (g30223), .I1 (g28702), .I2 (g23895));
AN4X1 gate13454(.O (g13805), .I1 (g11489), .I2 (g11394), .I3 (g11356), .I4 (I16129));
AN2X1 gate13455(.O (g18788), .I1 (g6031), .I2 (g15634));
AN2X1 gate13456(.O (g18724), .I1 (g4907), .I2 (g16077));
AN2X1 gate13457(.O (g25884), .I1 (g11153), .I2 (g24711));
AN2X1 gate13458(.O (g18359), .I1 (g1825), .I2 (g17955));
AN2X1 gate13459(.O (g34223), .I1 (g33744), .I2 (g22876));
AN2X1 gate13460(.O (g18325), .I1 (g1624), .I2 (g17873));
AN2X1 gate13461(.O (g26186), .I1 (g24580), .I2 (g23031));
AN2X1 gate13462(.O (g23436), .I1 (g676), .I2 (g20375));
AN2X1 gate13463(.O (g18535), .I1 (g2741), .I2 (g15277));
AN2X1 gate13464(.O (g18434), .I1 (g2217), .I2 (g18008));
AN2X1 gate13465(.O (g18358), .I1 (g1811), .I2 (g17955));
AN2X1 gate13466(.O (g31966), .I1 (g31754), .I2 (g22166));
AN2X1 gate13467(.O (g30084), .I1 (g28534), .I2 (g20700));
AN2X1 gate13468(.O (g27521), .I1 (g26519), .I2 (g14700));
AN2X1 gate13469(.O (g29337), .I1 (g29166), .I2 (g22180));
AN2X1 gate13470(.O (g17786), .I1 (g1489), .I2 (g13216));
AN2X1 gate13471(.O (g30110), .I1 (g28564), .I2 (g20916));
AN2X1 gate13472(.O (g25479), .I1 (g22646), .I2 (g9917));
AN2X1 gate13473(.O (g34084), .I1 (g9214), .I2 (g33851));
AN2X1 gate13474(.O (g15075), .I1 (g12850), .I2 (g12955));
AN2X1 gate13475(.O (g31017), .I1 (g29479), .I2 (g22841));
AN2X1 gate13476(.O (g34110), .I1 (g33732), .I2 (g22935));
AN2X1 gate13477(.O (g25217), .I1 (g12418), .I2 (g23698));
AN2X1 gate13478(.O (g33364), .I1 (g32264), .I2 (g20921));
AN2X1 gate13479(.O (g18121), .I1 (g424), .I2 (g17015));
AN2X1 gate13480(.O (g22090), .I1 (g6404), .I2 (g18833));
AN2X1 gate13481(.O (g30179), .I1 (g28634), .I2 (g23819));
AN2X1 gate13482(.O (g24507), .I1 (g22304), .I2 (g19429));
AN2X1 gate13483(.O (g18344), .I1 (g1740), .I2 (g17955));
AN3X1 gate13484(.O (g19581), .I1 (g15843), .I2 (g1500), .I3 (g10918));
AN2X1 gate13485(.O (g34179), .I1 (g33686), .I2 (g24372));
AN4X1 gate13486(.O (g27440), .I1 (g8046), .I2 (g26314), .I3 (g518), .I4 (g504));
AN2X1 gate13487(.O (g21464), .I1 (g16181), .I2 (g10872));
AN4X1 gate13488(.O (g28020), .I1 (g23032), .I2 (g26241), .I3 (g26424), .I4 (g25542));
AN2X1 gate13489(.O (g28583), .I1 (g12009), .I2 (g27112));
AN2X1 gate13490(.O (g30178), .I1 (g28632), .I2 (g23815));
AN2X1 gate13491(.O (g9479), .I1 (g305), .I2 (g324));
AN2X1 gate13492(.O (g24421), .I1 (g3835), .I2 (g23139));
AN2X1 gate13493(.O (g34178), .I1 (g33712), .I2 (g24361));
AN2X1 gate13494(.O (g34740), .I1 (g34664), .I2 (g19414));
AN2X1 gate13495(.O (g16616), .I1 (g6267), .I2 (g14741));
AN4X1 gate13496(.O (g10756), .I1 (g3990), .I2 (g6928), .I3 (g3976), .I4 (g8595));
AN2X1 gate13497(.O (g18682), .I1 (g4646), .I2 (g15885));
AN4X1 gate13498(.O (I31176), .I1 (g31579), .I2 (g31827), .I3 (g32708), .I4 (g32709));
AN2X1 gate13499(.O (g30186), .I1 (g28641), .I2 (g23839));
AN2X1 gate13500(.O (g27247), .I1 (g2759), .I2 (g26745));
AN4X1 gate13501(.O (I31092), .I1 (g32589), .I2 (g32590), .I3 (g32591), .I4 (g32592));
AN2X1 gate13502(.O (g18291), .I1 (g1437), .I2 (g16449));
AN2X1 gate13503(.O (g24012), .I1 (g14496), .I2 (g21561));
AN2X1 gate13504(.O (g17182), .I1 (g8579), .I2 (g13016));
AN2X1 gate13505(.O (g21797), .I1 (g3518), .I2 (g20924));
AN2X1 gate13506(.O (g34186), .I1 (g33705), .I2 (g24396));
AN2X1 gate13507(.O (g34685), .I1 (g14164), .I2 (g34550));
AN2X1 gate13508(.O (g25580), .I1 (g19268), .I2 (g24149));
AN2X1 gate13509(.O (g18173), .I1 (g736), .I2 (g17328));
AN2X1 gate13510(.O (g27389), .I1 (g26519), .I2 (g17503));
AN2X1 gate13511(.O (g34953), .I1 (g34935), .I2 (g19957));
AN4X1 gate13512(.O (g27045), .I1 (g10295), .I2 (g3171), .I3 (g3179), .I4 (g26244));
AN2X1 gate13513(.O (g31309), .I1 (g30132), .I2 (g27837));
AN4X1 gate13514(.O (I24699), .I1 (g21127), .I2 (g24054), .I3 (g24055), .I4 (g24056));
AN2X1 gate13515(.O (g32083), .I1 (g947), .I2 (g30735));
AN2X1 gate13516(.O (g32348), .I1 (g2145), .I2 (g31672));
AN2X1 gate13517(.O (g23292), .I1 (g19879), .I2 (g16726));
AN2X1 gate13518(.O (g25223), .I1 (g22523), .I2 (g10652));
AN2X1 gate13519(.O (g16704), .I1 (g5957), .I2 (g15018));
AN2X1 gate13520(.O (g27612), .I1 (g25887), .I2 (g8844));
AN2X1 gate13521(.O (g31224), .I1 (g30280), .I2 (g23932));
AN2X1 gate13522(.O (g32284), .I1 (g31260), .I2 (g20507));
AN2X1 gate13523(.O (g28113), .I1 (g8016), .I2 (g27242));
AN2X1 gate13524(.O (g26423), .I1 (g19488), .I2 (g24356));
AN2X1 gate13525(.O (g27099), .I1 (g14094), .I2 (g26352));
AN2X1 gate13526(.O (g15822), .I1 (g3925), .I2 (g13960));
AN2X1 gate13527(.O (g27388), .I1 (g26519), .I2 (g17502));
AN2X1 gate13528(.O (g27324), .I1 (g10150), .I2 (g26720));
AN2X1 gate13529(.O (g24541), .I1 (g22626), .I2 (g10851));
AN2X1 gate13530(.O (g32304), .I1 (g31284), .I2 (g20564));
AN2X1 gate13531(.O (g30936), .I1 (g8830), .I2 (g29916));
AN2X1 gate13532(.O (g28282), .I1 (g23762), .I2 (g27727));
AN2X1 gate13533(.O (g12099), .I1 (g9619), .I2 (g9888));
AN2X1 gate13534(.O (g27534), .I1 (g26488), .I2 (g17735));
AN2X1 gate13535(.O (g27098), .I1 (g25868), .I2 (g22528));
AN2X1 gate13536(.O (g28302), .I1 (g23809), .I2 (g27817));
AN2X1 gate13537(.O (g25084), .I1 (g4737), .I2 (g22885));
AN2X1 gate13538(.O (g27251), .I1 (g26721), .I2 (g26694));
AN2X1 gate13539(.O (g27272), .I1 (g26055), .I2 (g17144));
AN2X1 gate13540(.O (g25110), .I1 (g10427), .I2 (g23509));
AN2X1 gate13541(.O (g16808), .I1 (g6653), .I2 (g14825));
AN2X1 gate13542(.O (g19384), .I1 (g667), .I2 (g16310));
AN2X1 gate13543(.O (g18760), .I1 (g5462), .I2 (g17929));
AN2X1 gate13544(.O (g18134), .I1 (g534), .I2 (g17249));
AN2X1 gate13545(.O (g25922), .I1 (g24959), .I2 (g20065));
AN2X1 gate13546(.O (g34334), .I1 (g34090), .I2 (g19865));
AN2X1 gate13547(.O (g24788), .I1 (g11384), .I2 (g23111));
AN2X1 gate13548(.O (g31495), .I1 (g1913), .I2 (g30309));
AN2X1 gate13549(.O (g24724), .I1 (g17624), .I2 (g22432));
AN2X1 gate13550(.O (g29599), .I1 (g1710), .I2 (g29018));
AN3X1 gate13551(.O (g33495), .I1 (g32707), .I2 (I31171), .I3 (I31172));
AN2X1 gate13552(.O (g22717), .I1 (g9291), .I2 (g20212));
AN2X1 gate13553(.O (g16177), .I1 (g5128), .I2 (g14238));
AN2X1 gate13554(.O (g24325), .I1 (g4543), .I2 (g22228));
AN2X1 gate13555(.O (g25179), .I1 (g16928), .I2 (g23611));
AN2X1 gate13556(.O (g26543), .I1 (g12910), .I2 (g24377));
AN4X1 gate13557(.O (I27503), .I1 (g19890), .I2 (g24075), .I3 (g24076), .I4 (g28032));
AN2X1 gate13558(.O (g18506), .I1 (g2571), .I2 (g15509));
AN2X1 gate13559(.O (g22026), .I1 (g5913), .I2 (g19147));
AN2X1 gate13560(.O (g27462), .I1 (g26576), .I2 (g17612));
AN2X1 gate13561(.O (g33816), .I1 (g33234), .I2 (g20096));
AN2X1 gate13562(.O (g29598), .I1 (g28823), .I2 (g22342));
AN2X1 gate13563(.O (g16642), .I1 (g6633), .I2 (g14981));
AN2X1 gate13564(.O (g25178), .I1 (g20241), .I2 (g23608));
AN2X1 gate13565(.O (g15589), .I1 (g411), .I2 (g13334));
AN2X1 gate13566(.O (g32139), .I1 (g31601), .I2 (g29960));
AN4X1 gate13567(.O (g27032), .I1 (g7704), .I2 (g5180), .I3 (g5188), .I4 (g26200));
AN2X1 gate13568(.O (g34964), .I1 (g34947), .I2 (g23060));
AN2X1 gate13569(.O (g33687), .I1 (g33132), .I2 (g4878));
AN2X1 gate13570(.O (g31976), .I1 (g31762), .I2 (g22178));
AN2X1 gate13571(.O (g31985), .I1 (g4722), .I2 (g30614));
AN2X1 gate13572(.O (g19735), .I1 (g9740), .I2 (g17135));
AN2X1 gate13573(.O (g27140), .I1 (g25885), .I2 (g22593));
AN2X1 gate13574(.O (g30216), .I1 (g28691), .I2 (g23882));
AN2X1 gate13575(.O (g27997), .I1 (g26813), .I2 (g23995));
AN4X1 gate13576(.O (g28768), .I1 (g21434), .I2 (g26424), .I3 (g25308), .I4 (g27421));
AN2X1 gate13577(.O (g15836), .I1 (g3187), .I2 (g14104));
AN2X1 gate13578(.O (g31752), .I1 (g30104), .I2 (g23928));
AN2X1 gate13579(.O (g34216), .I1 (g33778), .I2 (g22689));
AN2X1 gate13580(.O (g31374), .I1 (g29748), .I2 (g23390));
AN3X1 gate13581(.O (g29322), .I1 (g29192), .I2 (g7074), .I3 (g6336));
AN2X1 gate13582(.O (g33374), .I1 (g32289), .I2 (g21221));
AN2X1 gate13583(.O (g16733), .I1 (g5893), .I2 (g14889));
AN3X1 gate13584(.O (I18671), .I1 (g13156), .I2 (g11450), .I3 (g6756));
AN2X1 gate13585(.O (g29532), .I1 (g1878), .I2 (g28861));
AN2X1 gate13586(.O (g29901), .I1 (g28429), .I2 (g23376));
AN2X1 gate13587(.O (g32333), .I1 (g31326), .I2 (g23559));
AN2X1 gate13588(.O (g15119), .I1 (g4249), .I2 (g14454));
AN2X1 gate13589(.O (g20682), .I1 (g16238), .I2 (g4646));
AN4X1 gate13590(.O (g13771), .I1 (g11441), .I2 (g11355), .I3 (g11302), .I4 (I16111));
AN3X1 gate13591(.O (g25417), .I1 (g5712), .I2 (g23816), .I3 (I24552));
AN2X1 gate13592(.O (g23474), .I1 (g13830), .I2 (g20533));
AN2X1 gate13593(.O (g24682), .I1 (g22662), .I2 (g19754));
AN2X1 gate13594(.O (g22149), .I1 (g14581), .I2 (g18880));
AN2X1 gate13595(.O (g29783), .I1 (g28329), .I2 (g23246));
AN2X1 gate13596(.O (g21711), .I1 (g291), .I2 (g20283));
AN2X1 gate13597(.O (g26123), .I1 (g1696), .I2 (g25382));
AN2X1 gate13598(.O (g15118), .I1 (g4253), .I2 (g14454));
AN2X1 gate13599(.O (g34909), .I1 (g34856), .I2 (g20130));
AN2X1 gate13600(.O (g24291), .I1 (g18660), .I2 (g22550));
AN2X1 gate13601(.O (g30000), .I1 (g23685), .I2 (g29029));
AN2X1 gate13602(.O (g29656), .I1 (g28515), .I2 (g11666));
AN2X1 gate13603(.O (g34117), .I1 (g33742), .I2 (g19755));
AN2X1 gate13604(.O (g15749), .I1 (g1454), .I2 (g13273));
AN2X1 gate13605(.O (g18649), .I1 (g4049), .I2 (g17271));
AN2X1 gate13606(.O (g22097), .I1 (g6451), .I2 (g18833));
AN2X1 gate13607(.O (g27360), .I1 (g26488), .I2 (g17417));
AN2X1 gate13608(.O (g33842), .I1 (g33255), .I2 (g20322));
AN2X1 gate13609(.O (g18240), .I1 (g15066), .I2 (g16431));
AN2X1 gate13610(.O (g22104), .I1 (g6444), .I2 (g18833));
AN2X1 gate13611(.O (g17149), .I1 (g232), .I2 (g13255));
AN2X1 gate13612(.O (g33392), .I1 (g32344), .I2 (g21362));
AN2X1 gate13613(.O (g18648), .I1 (g4045), .I2 (g17271));
AN2X1 gate13614(.O (g18491), .I1 (g2518), .I2 (g15426));
AN2X1 gate13615(.O (g31489), .I1 (g2204), .I2 (g30305));
AN2X1 gate13616(.O (g26230), .I1 (g1768), .I2 (g25385));
AN2X1 gate13617(.O (g25964), .I1 (g1783), .I2 (g24979));
AN3X1 gate13618(.O (g33489), .I1 (g32665), .I2 (I31141), .I3 (I31142));
AN2X1 gate13619(.O (g21606), .I1 (g15959), .I2 (g13763));
AN3X1 gate13620(.O (g27162), .I1 (g26171), .I2 (g8259), .I3 (g2208));
AN2X1 gate13621(.O (g34568), .I1 (g34379), .I2 (g17512));
AN2X1 gate13622(.O (g34747), .I1 (g34671), .I2 (g19527));
AN2X1 gate13623(.O (g23606), .I1 (g16927), .I2 (g20679));
AN2X1 gate13624(.O (g29336), .I1 (g4704), .I2 (g28363));
AN2X1 gate13625(.O (g15704), .I1 (g3440), .I2 (g13504));
AN2X1 gate13626(.O (g30242), .I1 (g28730), .I2 (g23927));
AN2X1 gate13627(.O (g18604), .I1 (g3125), .I2 (g16987));
AN2X1 gate13628(.O (g21303), .I1 (g10120), .I2 (g17625));
AN2X1 gate13629(.O (g16485), .I1 (g5563), .I2 (g14924));
AN2X1 gate13630(.O (g18755), .I1 (g5343), .I2 (g15595));
AN2X1 gate13631(.O (g31525), .I1 (g29892), .I2 (g23526));
AN2X1 gate13632(.O (g31488), .I1 (g1779), .I2 (g30302));
AN2X1 gate13633(.O (g31016), .I1 (g29478), .I2 (g22840));
AN3X1 gate13634(.O (g33525), .I1 (g32925), .I2 (I31321), .I3 (I31322));
AN3X1 gate13635(.O (g33488), .I1 (g32658), .I2 (I31136), .I3 (I31137));
AN2X1 gate13636(.O (g28249), .I1 (g27152), .I2 (g19677));
AN2X1 gate13637(.O (g15809), .I1 (g3917), .I2 (g14154));
AN2X1 gate13638(.O (g18770), .I1 (g15153), .I2 (g15615));
AN3X1 gate13639(.O (g22369), .I1 (g9354), .I2 (g7717), .I3 (g20783));
AN2X1 gate13640(.O (g18563), .I1 (g2890), .I2 (g16349));
AN2X1 gate13641(.O (g18981), .I1 (g11206), .I2 (g16158));
AN2X1 gate13642(.O (g21750), .I1 (g3161), .I2 (g20785));
AN2X1 gate13643(.O (g28248), .I1 (g27150), .I2 (g19676));
AN2X1 gate13644(.O (g29966), .I1 (g23617), .I2 (g28970));
AN2X1 gate13645(.O (g28710), .I1 (g27589), .I2 (g20703));
AN2X1 gate13646(.O (g15808), .I1 (g3590), .I2 (g14048));
AN2X1 gate13647(.O (g21982), .I1 (g5547), .I2 (g19074));
AN2X1 gate13648(.O (g27451), .I1 (g26400), .I2 (g17599));
AN2X1 gate13649(.O (g26391), .I1 (g19593), .I2 (g25555));
AN3X1 gate13650(.O (I26948), .I1 (g24981), .I2 (g26424), .I3 (g22698));
AN2X1 gate13651(.O (g23381), .I1 (g7239), .I2 (g21413));
AN2X1 gate13652(.O (g27220), .I1 (g26026), .I2 (g16743));
AN2X1 gate13653(.O (g33830), .I1 (g33382), .I2 (g20166));
AN2X1 gate13654(.O (g29631), .I1 (g1682), .I2 (g28656));
AN2X1 gate13655(.O (g32312), .I1 (g31302), .I2 (g20591));
AN2X1 gate13656(.O (g32200), .I1 (g27468), .I2 (g31376));
AN2X1 gate13657(.O (g33893), .I1 (g33313), .I2 (g20706));
AN2X1 gate13658(.O (g28204), .I1 (g26098), .I2 (g27654));
AN2X1 gate13659(.O (g27628), .I1 (g26400), .I2 (g18061));
AN2X1 gate13660(.O (g34751), .I1 (g34674), .I2 (g19543));
AN2X1 gate13661(.O (g29364), .I1 (g27400), .I2 (g28321));
AN2X1 gate13662(.O (g10827), .I1 (g8914), .I2 (g4258));
AN2X1 gate13663(.O (g25909), .I1 (g8745), .I2 (g24875));
AN2X1 gate13664(.O (g32115), .I1 (g31631), .I2 (g29928));
AN2X1 gate13665(.O (g25543), .I1 (g23795), .I2 (g21461));
AN2X1 gate13666(.O (g12220), .I1 (g1521), .I2 (g7535));
AN2X1 gate13667(.O (g27246), .I1 (g26690), .I2 (g26673));
AN2X1 gate13668(.O (g33865), .I1 (g33275), .I2 (g20526));
AN2X1 gate13669(.O (g21796), .I1 (g3512), .I2 (g20924));
AN2X1 gate13670(.O (g30230), .I1 (g28717), .I2 (g23906));
AN2X1 gate13671(.O (g25908), .I1 (g24782), .I2 (g22520));
AN2X1 gate13672(.O (g18767), .I1 (g15150), .I2 (g17929));
AN2X1 gate13673(.O (g18794), .I1 (g6154), .I2 (g15348));
AN2X1 gate13674(.O (g34230), .I1 (g33761), .I2 (g22942));
AN2X1 gate13675(.O (g18395), .I1 (g12849), .I2 (g15373));
AN2X1 gate13676(.O (g32052), .I1 (g31507), .I2 (g13885));
AN2X1 gate13677(.O (g18262), .I1 (g1259), .I2 (g16000));
AN2X1 gate13678(.O (g22133), .I1 (g6649), .I2 (g19277));
AN2X1 gate13679(.O (g25569), .I1 (I24684), .I2 (I24685));
AN2X1 gate13680(.O (g21840), .I1 (g15099), .I2 (g21070));
AN2X1 gate13681(.O (g25568), .I1 (I24679), .I2 (I24680));
AN2X1 gate13682(.O (g18633), .I1 (g6905), .I2 (g17226));
AN2X1 gate13683(.O (g17133), .I1 (g10683), .I2 (g13222));
AN2X1 gate13684(.O (g34841), .I1 (g34761), .I2 (g20080));
AN2X1 gate13685(.O (g18191), .I1 (g827), .I2 (g17821));
AN2X1 gate13686(.O (g18719), .I1 (g4894), .I2 (g16795));
AN2X1 gate13687(.O (g22011), .I1 (g15154), .I2 (g21562));
AN2X1 gate13688(.O (g15874), .I1 (g3893), .I2 (g14079));
AN2X1 gate13689(.O (g24649), .I1 (g6527), .I2 (g23733));
AN2X1 gate13690(.O (g29571), .I1 (g28452), .I2 (g11762));
AN2X1 gate13691(.O (g11114), .I1 (g5689), .I2 (g10160));
AN2X1 gate13692(.O (g31270), .I1 (g29692), .I2 (g23282));
AN2X1 gate13693(.O (g16519), .I1 (g5591), .I2 (g14804));
AN2X1 gate13694(.O (g16176), .I1 (g14596), .I2 (g11779));
AN2X1 gate13695(.O (g16185), .I1 (g3263), .I2 (g14011));
AN2X1 gate13696(.O (g25123), .I1 (g4732), .I2 (g22885));
AN2X1 gate13697(.O (g18718), .I1 (g4854), .I2 (g15915));
AN2X1 gate13698(.O (g15693), .I1 (g269), .I2 (g13474));
AN2X1 gate13699(.O (g18521), .I1 (g2667), .I2 (g15509));
AN2X1 gate13700(.O (g31188), .I1 (g20028), .I2 (g29653));
AN2X1 gate13701(.O (g25814), .I1 (g24760), .I2 (g13323));
AN2X1 gate13702(.O (g27370), .I1 (g26400), .I2 (g17472));
AN2X1 gate13703(.O (g31124), .I1 (g2259), .I2 (g29997));
AN2X1 gate13704(.O (g32184), .I1 (g30611), .I2 (g25249));
AN4X1 gate13705(.O (g28998), .I1 (g17424), .I2 (g25212), .I3 (g26424), .I4 (g27474));
AN2X1 gate13706(.O (g33124), .I1 (g8945), .I2 (g32296));
AN3X1 gate13707(.O (g33678), .I1 (g33149), .I2 (g10710), .I3 (g22319));
AN2X1 gate13708(.O (g24491), .I1 (g10727), .I2 (g22332));
AN2X1 gate13709(.O (g24903), .I1 (g128), .I2 (g23889));
AN2X1 gate13710(.O (g28233), .I1 (g27827), .I2 (g23411));
AN2X1 gate13711(.O (g16518), .I1 (g5571), .I2 (g14956));
AN2X1 gate13712(.O (g28182), .I1 (g8770), .I2 (g27349));
AN2X1 gate13713(.O (g25772), .I1 (g24944), .I2 (g24934));
AN2X1 gate13714(.O (g28672), .I1 (g7577), .I2 (g27017));
AN2X1 gate13715(.O (g24755), .I1 (g16022), .I2 (g23030));
AN2X1 gate13716(.O (g27151), .I1 (g26026), .I2 (g16626));
AN2X1 gate13717(.O (g34578), .I1 (g24578), .I2 (g34308));
AN2X1 gate13718(.O (g16637), .I1 (g5949), .I2 (g14968));
AN2X1 gate13719(.O (g22310), .I1 (g19662), .I2 (g20235));
AN2X1 gate13720(.O (g18440), .I1 (g2255), .I2 (g18008));
AN2X1 gate13721(.O (g13345), .I1 (g4754), .I2 (g11773));
AN2X1 gate13722(.O (g26275), .I1 (g2417), .I2 (g25349));
AN2X1 gate13723(.O (g30007), .I1 (g29141), .I2 (g12929));
AN3X1 gate13724(.O (I24546), .I1 (g5046), .I2 (g5052), .I3 (g9716));
AN2X1 gate13725(.O (g34586), .I1 (g11025), .I2 (g34317));
AN2X1 gate13726(.O (g18573), .I1 (g2898), .I2 (g16349));
AN2X1 gate13727(.O (g29687), .I1 (g2407), .I2 (g29097));
AN2X1 gate13728(.O (g22112), .I1 (g6555), .I2 (g19277));
AN2X1 gate13729(.O (g18247), .I1 (g1178), .I2 (g16431));
AN2X1 gate13730(.O (g29985), .I1 (g28127), .I2 (g20532));
AN2X1 gate13731(.O (g10890), .I1 (g7858), .I2 (g1105));
AN2X1 gate13732(.O (g21862), .I1 (g3953), .I2 (g21070));
AN2X1 gate13733(.O (g22050), .I1 (g6088), .I2 (g21611));
AN2X1 gate13734(.O (g23553), .I1 (g19413), .I2 (g11875));
AN2X1 gate13735(.O (g18389), .I1 (g1974), .I2 (g15171));
AN2X1 gate13736(.O (g29752), .I1 (g28516), .I2 (g10233));
AN4X1 gate13737(.O (I31312), .I1 (g32905), .I2 (g32906), .I3 (g32907), .I4 (g32908));
AN2X1 gate13738(.O (g29954), .I1 (g2299), .I2 (g28796));
AN2X1 gate13739(.O (g21949), .I1 (g5264), .I2 (g18997));
AN2X1 gate13740(.O (g15712), .I1 (g3791), .I2 (g13521));
AN2X1 gate13741(.O (g18612), .I1 (g3329), .I2 (g17200));
AN2X1 gate13742(.O (g15914), .I1 (g3905), .I2 (g14024));
AN2X1 gate13743(.O (g25992), .I1 (g2485), .I2 (g25024));
AN2X1 gate13744(.O (g18388), .I1 (g1968), .I2 (g15171));
AN2X1 gate13745(.O (g19660), .I1 (g12001), .I2 (g16968));
AN2X1 gate13746(.O (g18324), .I1 (g1644), .I2 (g17873));
AN2X1 gate13747(.O (g24794), .I1 (g11414), .I2 (g23138));
AN2X1 gate13748(.O (g31219), .I1 (g30265), .I2 (g20875));
AN2X1 gate13749(.O (g34116), .I1 (g33933), .I2 (g25140));
AN2X1 gate13750(.O (g24395), .I1 (g4704), .I2 (g22845));
AN3X1 gate13751(.O (g25510), .I1 (g6444), .I2 (g22300), .I3 (I24619));
AN2X1 gate13752(.O (g18701), .I1 (g4771), .I2 (g16856));
AN2X1 gate13753(.O (g26684), .I1 (g25407), .I2 (g20673));
AN2X1 gate13754(.O (g21948), .I1 (g5260), .I2 (g18997));
AN2X1 gate13755(.O (g22096), .I1 (g6434), .I2 (g18833));
AN2X1 gate13756(.O (g32400), .I1 (g4743), .I2 (g30989));
AN2X1 gate13757(.O (g18777), .I1 (g5808), .I2 (g18065));
AN2X1 gate13758(.O (g18534), .I1 (g2735), .I2 (g15277));
AN4X1 gate13759(.O (I14198), .I1 (g225), .I2 (g8237), .I3 (g232), .I4 (g8180));
AN2X1 gate13760(.O (g32013), .I1 (g8673), .I2 (g30614));
AN2X1 gate13761(.O (g30041), .I1 (g28511), .I2 (g23518));
AN4X1 gate13762(.O (I31052), .I1 (g32531), .I2 (g32532), .I3 (g32533), .I4 (g32534));
AN2X1 gate13763(.O (g18251), .I1 (g996), .I2 (g16897));
AN2X1 gate13764(.O (g21702), .I1 (g157), .I2 (g20283));
AN2X1 gate13765(.O (g31218), .I1 (g30271), .I2 (g23909));
AN2X1 gate13766(.O (g16729), .I1 (g5240), .I2 (g14720));
AN2X1 gate13767(.O (g18272), .I1 (g1283), .I2 (g16031));
AN2X1 gate13768(.O (g21757), .I1 (g3187), .I2 (g20785));
AN2X1 gate13769(.O (g25579), .I1 (g19422), .I2 (g24147));
AN2X1 gate13770(.O (g30275), .I1 (g28816), .I2 (g23984));
AN4X1 gate13771(.O (I24700), .I1 (g24057), .I2 (g24058), .I3 (g24059), .I4 (g24060));
AN2X1 gate13772(.O (g27227), .I1 (g26026), .I2 (g16771));
AN2X1 gate13773(.O (g33837), .I1 (g33251), .I2 (g20233));
AN3X1 gate13774(.O (I24625), .I1 (g6428), .I2 (g6434), .I3 (g10014));
AN2X1 gate13775(.O (g32207), .I1 (g31221), .I2 (g23323));
AN2X1 gate13776(.O (g26517), .I1 (g15708), .I2 (g24367));
AN2X1 gate13777(.O (g34746), .I1 (g34670), .I2 (g19526));
AN2X1 gate13778(.O (g34493), .I1 (g34273), .I2 (g19360));
AN2X1 gate13779(.O (g25578), .I1 (g19402), .I2 (g24146));
AN2X1 gate13780(.O (g15567), .I1 (g392), .I2 (g13312));
AN2X1 gate13781(.O (g27025), .I1 (g26334), .I2 (g7917));
AN2X1 gate13782(.O (g24191), .I1 (g319), .I2 (g22722));
AN2X1 gate13783(.O (g24719), .I1 (g681), .I2 (g23530));
AN2X1 gate13784(.O (g18462), .I1 (g2361), .I2 (g15224));
AN2X1 gate13785(.O (g25014), .I1 (g17474), .I2 (g23420));
AN2X1 gate13786(.O (g32328), .I1 (g5853), .I2 (g31554));
AN2X1 gate13787(.O (g29668), .I1 (g28527), .I2 (g14255));
AN2X1 gate13788(.O (g29842), .I1 (g28372), .I2 (g23284));
AN2X1 gate13789(.O (g27540), .I1 (g26576), .I2 (g17746));
AN2X1 gate13790(.O (g23564), .I1 (g16882), .I2 (g20648));
AN4X1 gate13791(.O (g27058), .I1 (g10323), .I2 (g3522), .I3 (g3530), .I4 (g26264));
AN2X1 gate13792(.O (g30035), .I1 (g22539), .I2 (g28120));
AN2X1 gate13793(.O (g18140), .I1 (g559), .I2 (g17533));
AN2X1 gate13794(.O (g34340), .I1 (g34100), .I2 (g19950));
AN2X1 gate13795(.O (g27203), .I1 (g26026), .I2 (g16688));
AN2X1 gate13796(.O (g19596), .I1 (g1094), .I2 (g16681));
AN2X1 gate13797(.O (g26130), .I1 (g24890), .I2 (g19772));
AN2X1 gate13798(.O (g29525), .I1 (g2169), .I2 (g28837));
AN2X1 gate13799(.O (g21847), .I1 (g3905), .I2 (g21070));
AN2X1 gate13800(.O (g34684), .I1 (g14178), .I2 (g34545));
AN2X1 gate13801(.O (g10999), .I1 (g7880), .I2 (g1472));
AN2X1 gate13802(.O (g13833), .I1 (g4546), .I2 (g10613));
AN3X1 gate13803(.O (I18819), .I1 (g13156), .I2 (g11450), .I3 (g11498));
AN2X1 gate13804(.O (g26362), .I1 (g19557), .I2 (g25538));
AN4X1 gate13805(.O (g27044), .I1 (g7766), .I2 (g5873), .I3 (g5881), .I4 (g26241));
AN2X1 gate13806(.O (g31470), .I1 (g29753), .I2 (g23398));
AN2X1 gate13807(.O (g23397), .I1 (g11154), .I2 (g20239));
AN3X1 gate13808(.O (g33470), .I1 (g32528), .I2 (I31046), .I3 (I31047));
AN2X1 gate13809(.O (g33915), .I1 (g33140), .I2 (g7846));
AN2X1 gate13810(.O (g32241), .I1 (g31244), .I2 (g20323));
AN2X1 gate13811(.O (g26165), .I1 (g11980), .I2 (g25153));
AN4X1 gate13812(.O (g17793), .I1 (g6772), .I2 (g11592), .I3 (g6789), .I4 (I18803));
AN4X1 gate13813(.O (g10998), .I1 (g8567), .I2 (g8509), .I3 (g8451), .I4 (g7650));
AN2X1 gate13814(.O (g18766), .I1 (g5495), .I2 (g17929));
AN2X1 gate13815(.O (g13048), .I1 (g8558), .I2 (g11043));
AN2X1 gate13816(.O (g23062), .I1 (g718), .I2 (g20248));
AN2X1 gate13817(.O (g27281), .I1 (g9830), .I2 (g26615));
AN3X1 gate13818(.O (g24861), .I1 (g3712), .I2 (g23582), .I3 (I24033));
AN2X1 gate13819(.O (g24573), .I1 (g17198), .I2 (g23716));
AN2X1 gate13820(.O (g34517), .I1 (g34290), .I2 (g19493));
AN2X1 gate13821(.O (g28148), .I1 (g27355), .I2 (g26093));
AN2X1 gate13822(.O (g14233), .I1 (g8639), .I2 (g11855));
AN2X1 gate13823(.O (g21933), .I1 (g5212), .I2 (g18997));
AN2X1 gate13824(.O (g27301), .I1 (g11992), .I2 (g26679));
AN4X1 gate13825(.O (I14225), .I1 (g8457), .I2 (g255), .I3 (g8406), .I4 (g262));
AN2X1 gate13826(.O (g27957), .I1 (g25947), .I2 (g15995));
AN2X1 gate13827(.O (g7804), .I1 (g2975), .I2 (g2970));
AN2X1 gate13828(.O (g25041), .I1 (g23261), .I2 (g20494));
AN2X1 gate13829(.O (g13221), .I1 (g6946), .I2 (g11425));
AN2X1 gate13830(.O (g27120), .I1 (g25878), .I2 (g22543));
AN4X1 gate13831(.O (g17690), .I1 (g11547), .I2 (g11592), .I3 (g11640), .I4 (I18671));
AN2X1 gate13832(.O (g29865), .I1 (g1802), .I2 (g29115));
AN2X1 gate13833(.O (g21851), .I1 (g3901), .I2 (g21070));
AN2X1 gate13834(.O (g21872), .I1 (g4098), .I2 (g19801));
AN2X1 gate13835(.O (g23872), .I1 (g19389), .I2 (g4157));
AN2X1 gate13836(.O (g15883), .I1 (g9180), .I2 (g14258));
AN2X1 gate13837(.O (g18360), .I1 (g1830), .I2 (g17955));
AN2X1 gate13838(.O (g31467), .I1 (g30162), .I2 (g27937));
AN2X1 gate13839(.O (g31494), .I1 (g29792), .I2 (g23435));
AN2X1 gate13840(.O (g28343), .I1 (g27380), .I2 (g19799));
AN3X1 gate13841(.O (I24527), .I1 (g9672), .I2 (g9264), .I3 (g5401));
AN2X1 gate13842(.O (g19655), .I1 (g2729), .I2 (g16966));
AN3X1 gate13843(.O (g33467), .I1 (g32505), .I2 (I31031), .I3 (I31032));
AN3X1 gate13844(.O (g33494), .I1 (g32700), .I2 (I31166), .I3 (I31167));
AN2X1 gate13845(.O (g24324), .I1 (g4540), .I2 (g22228));
AN3X1 gate13846(.O (g27146), .I1 (g26148), .I2 (g8187), .I3 (g1648));
AN2X1 gate13847(.O (g27645), .I1 (g26488), .I2 (g15344));
AN2X1 gate13848(.O (g26863), .I1 (g24974), .I2 (g24957));
AN2X1 gate13849(.O (g18447), .I1 (g2208), .I2 (g18008));
AN2X1 gate13850(.O (g30193), .I1 (g28650), .I2 (g23848));
AN2X1 gate13851(.O (g24777), .I1 (g11345), .I2 (g23066));
AN2X1 gate13852(.O (g27699), .I1 (g26396), .I2 (g20766));
AN2X1 gate13853(.O (g16653), .I1 (g8343), .I2 (g13850));
AN2X1 gate13854(.O (g18162), .I1 (g686), .I2 (g17433));
AN2X1 gate13855(.O (g25983), .I1 (g2476), .I2 (g25009));
AN2X1 gate13856(.O (g29610), .I1 (g28483), .I2 (g8026));
AN2X1 gate13857(.O (g30165), .I1 (g28619), .I2 (g23788));
AN2X1 gate13858(.O (g22129), .I1 (g6633), .I2 (g19277));
AN2X1 gate13859(.O (g34523), .I1 (g9162), .I2 (g34351));
AN2X1 gate13860(.O (g22002), .I1 (g5706), .I2 (g21562));
AN2X1 gate13861(.O (g22057), .I1 (g15159), .I2 (g21611));
AN2X1 gate13862(.O (g17317), .I1 (g1079), .I2 (g13124));
AN2X1 gate13863(.O (g22128), .I1 (g6629), .I2 (g19277));
AN2X1 gate13864(.O (g33352), .I1 (g32237), .I2 (g20712));
AN4X1 gate13865(.O (I31207), .I1 (g32754), .I2 (g32755), .I3 (g32756), .I4 (g32757));
AN2X1 gate13866(.O (g16636), .I1 (g5929), .I2 (g14768));
AN2X1 gate13867(.O (g18629), .I1 (g3680), .I2 (g17226));
AN2X1 gate13868(.O (g25142), .I1 (g4717), .I2 (g22885));
AN2X1 gate13869(.O (g18451), .I1 (g2295), .I2 (g15224));
AN2X1 gate13870(.O (g26347), .I1 (g262), .I2 (g24850));
AN2X1 gate13871(.O (g18472), .I1 (g2413), .I2 (g15224));
AN2X1 gate13872(.O (g32414), .I1 (g4944), .I2 (g30999));
AN2X1 gate13873(.O (g29188), .I1 (g27163), .I2 (g12762));
AN2X1 gate13874(.O (g33418), .I1 (g32372), .I2 (g21425));
AN2X1 gate13875(.O (g33822), .I1 (g33385), .I2 (g20157));
AN2X1 gate13876(.O (g18220), .I1 (g1002), .I2 (g16100));
AN2X1 gate13877(.O (g26253), .I1 (g2327), .I2 (g25435));
AN2X1 gate13878(.O (g30006), .I1 (g29032), .I2 (g9259));
AN2X1 gate13879(.O (g31266), .I1 (g30129), .I2 (g27742));
AN2X1 gate13880(.O (g31170), .I1 (g19128), .I2 (g29814));
AN2X1 gate13881(.O (g21452), .I1 (g16119), .I2 (g13624));
AN2X1 gate13882(.O (g18628), .I1 (g15095), .I2 (g17226));
AN2X1 gate13883(.O (g27427), .I1 (g26400), .I2 (g17575));
AN2X1 gate13884(.O (g34475), .I1 (g27450), .I2 (g34327));
AN2X1 gate13885(.O (g17057), .I1 (g446), .I2 (g13173));
AN2X1 gate13886(.O (g24140), .I1 (g17663), .I2 (g21654));
AN2X1 gate13887(.O (g22299), .I1 (g19999), .I2 (g21024));
AN2X1 gate13888(.O (g29686), .I1 (g2246), .I2 (g29057));
AN2X1 gate13889(.O (g24997), .I1 (g22929), .I2 (g10419));
AN2X1 gate13890(.O (g18246), .I1 (g1199), .I2 (g16431));
AN2X1 gate13891(.O (g21912), .I1 (g5052), .I2 (g21468));
AN2X1 gate13892(.O (g29383), .I1 (g28138), .I2 (g19412));
AN2X1 gate13893(.O (g30222), .I1 (g28701), .I2 (g23894));
AN2X1 gate13894(.O (g34863), .I1 (g16540), .I2 (g34833));
AN2X1 gate13895(.O (g28133), .I1 (g27367), .I2 (g23108));
AN2X1 gate13896(.O (g22298), .I1 (g19997), .I2 (g21012));
AN4X1 gate13897(.O (g26236), .I1 (g25357), .I2 (g6856), .I3 (g7586), .I4 (g7558));
AN2X1 gate13898(.O (g28229), .I1 (g27345), .I2 (g17213));
AN2X1 gate13899(.O (g19487), .I1 (g499), .I2 (g16680));
AN2X1 gate13900(.O (g29938), .I1 (g23552), .I2 (g28889));
AN2X1 gate13901(.O (g26351), .I1 (g239), .I2 (g24869));
AN2X1 gate13902(.O (g28228), .I1 (g27126), .I2 (g19636));
AN2X1 gate13903(.O (g25130), .I1 (g23358), .I2 (g20600));
AN2X1 gate13904(.O (g26821), .I1 (g24821), .I2 (g13103));
AN2X1 gate13905(.O (g27661), .I1 (g26576), .I2 (g15568));
AN4X1 gate13906(.O (I31241), .I1 (g30825), .I2 (g31838), .I3 (g32803), .I4 (g32804));
AN2X1 gate13907(.O (g27547), .I1 (g26549), .I2 (g17759));
AN2X1 gate13908(.O (g18591), .I1 (g2965), .I2 (g16349));
AN2X1 gate13909(.O (g31194), .I1 (g19128), .I2 (g29814));
AN2X1 gate13910(.O (g31167), .I1 (g10080), .I2 (g30076));
AN2X1 gate13911(.O (g18776), .I1 (g5813), .I2 (g18065));
AN2X1 gate13912(.O (g18785), .I1 (g5849), .I2 (g18065));
AN2X1 gate13913(.O (g15083), .I1 (g10362), .I2 (g12983));
AN2X1 gate13914(.O (g21756), .I1 (g3211), .I2 (g20785));
AN2X1 gate13915(.O (g18147), .I1 (g599), .I2 (g17533));
AN2X1 gate13916(.O (g25165), .I1 (g14062), .I2 (g23570));
AN2X1 gate13917(.O (g30253), .I1 (g28746), .I2 (g23943));
AN2X1 gate13918(.O (g16484), .I1 (g5244), .I2 (g14755));
AN2X1 gate13919(.O (g18754), .I1 (g5339), .I2 (g15595));
AN2X1 gate13920(.O (g31524), .I1 (g29897), .I2 (g20593));
AN3X1 gate13921(.O (g33524), .I1 (g32918), .I2 (I31316), .I3 (I31317));
AN2X1 gate13922(.O (g18355), .I1 (g1748), .I2 (g17955));
AN4X1 gate13923(.O (g26264), .I1 (g24688), .I2 (g8812), .I3 (g8778), .I4 (g10627));
AN2X1 gate13924(.O (g33836), .I1 (g33096), .I2 (g27020));
AN2X1 gate13925(.O (g21780), .I1 (g3391), .I2 (g20391));
AN2X1 gate13926(.O (g29875), .I1 (g28403), .I2 (g23337));
AN2X1 gate13927(.O (g32206), .I1 (g30609), .I2 (g25524));
AN2X1 gate13928(.O (g26516), .I1 (g24968), .I2 (g8876));
AN2X1 gate13929(.O (g13507), .I1 (g7023), .I2 (g12198));
AN2X1 gate13930(.O (g27481), .I1 (g26400), .I2 (g14630));
AN2X1 gate13931(.O (g30600), .I1 (g30287), .I2 (g18975));
AN2X1 gate13932(.O (g18825), .I1 (g6736), .I2 (g15680));
AN2X1 gate13933(.O (g18950), .I1 (g11193), .I2 (g16123));
AN2X1 gate13934(.O (g18370), .I1 (g1874), .I2 (g15171));
AN2X1 gate13935(.O (g31477), .I1 (g29763), .I2 (g23409));
AN2X1 gate13936(.O (g33401), .I1 (g32349), .I2 (g21381));
AN3X1 gate13937(.O (g33477), .I1 (g32577), .I2 (I31081), .I3 (I31082));
AN2X1 gate13938(.O (g20162), .I1 (g8737), .I2 (g16750));
AN2X1 gate13939(.O (g30236), .I1 (g28724), .I2 (g23916));
AN2X1 gate13940(.O (g14148), .I1 (g884), .I2 (g10632));
AN2X1 gate13941(.O (g29837), .I1 (g28369), .I2 (g20144));
AN2X1 gate13942(.O (g14097), .I1 (g878), .I2 (g10632));
AN2X1 gate13943(.O (g21820), .I1 (g3712), .I2 (g20453));
AN2X1 gate13944(.O (g11163), .I1 (g6727), .I2 (g10224));
AN3X1 gate13945(.O (I24067), .I1 (g3731), .I2 (g3736), .I3 (g8553));
AN2X1 gate13946(.O (g9906), .I1 (g996), .I2 (g1157));
AN2X1 gate13947(.O (g18151), .I1 (g617), .I2 (g17533));
AN2X1 gate13948(.O (g31118), .I1 (g29490), .I2 (g22906));
AN2X1 gate13949(.O (g18172), .I1 (g15058), .I2 (g17328));
AN2X1 gate13950(.O (g28627), .I1 (g27543), .I2 (g20574));
AN2X1 gate13951(.O (g32114), .I1 (g31624), .I2 (g29927));
AN4X1 gate13952(.O (g28959), .I1 (g17401), .I2 (g25194), .I3 (g26424), .I4 (g27440));
AN2X1 gate13953(.O (g30175), .I1 (g28629), .I2 (g23813));
AN2X1 gate13954(.O (g32082), .I1 (g4917), .I2 (g30673));
AN2X1 gate13955(.O (g33864), .I1 (g33274), .I2 (g20524));
AN2X1 gate13956(.O (g27127), .I1 (g25997), .I2 (g16582));
AN2X1 gate13957(.O (g21846), .I1 (g3897), .I2 (g21070));
AN2X1 gate13958(.O (g28112), .I1 (g27352), .I2 (g26162));
AN2X1 gate13959(.O (g32107), .I1 (g31624), .I2 (g29912));
AN2X1 gate13960(.O (g15653), .I1 (g3119), .I2 (g13530));
AN2X1 gate13961(.O (g24629), .I1 (g6163), .I2 (g23699));
AN2X1 gate13962(.O (g23396), .I1 (g20051), .I2 (g20229));
AN2X1 gate13963(.O (g18367), .I1 (g1783), .I2 (g17955));
AN2X1 gate13964(.O (g18394), .I1 (g1862), .I2 (g15171));
AN2X1 gate13965(.O (g31313), .I1 (g30160), .I2 (g27907));
AN2X1 gate13966(.O (g24451), .I1 (g3476), .I2 (g23112));
AN2X1 gate13967(.O (g21731), .I1 (g3029), .I2 (g20330));
AN2X1 gate13968(.O (g24220), .I1 (g255), .I2 (g22594));
AN2X1 gate13969(.O (g20628), .I1 (g1046), .I2 (g15789));
AN2X1 gate13970(.O (g27490), .I1 (g26576), .I2 (g17651));
AN2X1 gate13971(.O (g13541), .I1 (g7069), .I2 (g12308));
AN2X1 gate13972(.O (g30264), .I1 (g28774), .I2 (g23963));
AN2X1 gate13973(.O (g34063), .I1 (g33806), .I2 (g23121));
AN2X1 gate13974(.O (g13473), .I1 (g9797), .I2 (g11841));
AN2X1 gate13975(.O (g30137), .I1 (g28594), .I2 (g21181));
AN2X1 gate13976(.O (g19601), .I1 (g16198), .I2 (g11149));
AN2X1 gate13977(.O (g24628), .I1 (g5835), .I2 (g23666));
AN2X1 gate13978(.O (g32345), .I1 (g2138), .I2 (g31672));
AN2X1 gate13979(.O (g34137), .I1 (g33928), .I2 (g23802));
AN2X1 gate13980(.O (g31285), .I1 (g30134), .I2 (g27800));
AN2X1 gate13981(.O (g34516), .I1 (g34289), .I2 (g19492));
AN2X1 gate13982(.O (g27376), .I1 (g26549), .I2 (g17481));
AN2X1 gate13983(.O (g27385), .I1 (g26400), .I2 (g17497));
AN3X1 gate13984(.O (g33704), .I1 (g33176), .I2 (g10710), .I3 (g22319));
AN2X1 gate13985(.O (g29617), .I1 (g2024), .I2 (g28987));
AN2X1 gate13986(.O (g31305), .I1 (g29741), .I2 (g23354));
AN4X1 gate13987(.O (I24695), .I1 (g24050), .I2 (g24051), .I3 (g24052), .I4 (g24053));
AN3X1 gate13988(.O (I24018), .I1 (g8155), .I2 (g8390), .I3 (g3396));
AN2X1 gate13989(.O (g27103), .I1 (g25997), .I2 (g16509));
AN2X1 gate13990(.O (g33305), .I1 (g31935), .I2 (g17811));
AN2X1 gate13991(.O (g22831), .I1 (g19441), .I2 (g19629));
AN2X1 gate13992(.O (g23691), .I1 (g14731), .I2 (g20993));
AN2X1 gate13993(.O (g26542), .I1 (g13102), .I2 (g24376));
AN2X1 gate13994(.O (g34873), .I1 (g34830), .I2 (g20046));
AN2X1 gate13995(.O (g26021), .I1 (g9568), .I2 (g25035));
AN2X1 gate13996(.O (g18420), .I1 (g1996), .I2 (g15373));
AN2X1 gate13997(.O (g15852), .I1 (g13820), .I2 (g13223));
AN2X1 gate13998(.O (g27095), .I1 (g25997), .I2 (g16473));
AN2X1 gate13999(.O (g18319), .I1 (g1600), .I2 (g17873));
AN2X1 gate14000(.O (g33809), .I1 (g33432), .I2 (g30184));
AN2X1 gate14001(.O (g33900), .I1 (g33316), .I2 (g20913));
AN3X1 gate14002(.O (g33466), .I1 (g32498), .I2 (I31026), .I3 (I31027));
AN2X1 gate14003(.O (g16184), .I1 (g9285), .I2 (g14183));
AN2X1 gate14004(.O (g16805), .I1 (g7187), .I2 (g12972));
AN2X1 gate14005(.O (g21405), .I1 (g13377), .I2 (g15811));
AN2X1 gate14006(.O (g16674), .I1 (g6637), .I2 (g15014));
AN3X1 gate14007(.O (g29201), .I1 (g24081), .I2 (I27503), .I3 (I27504));
AN2X1 gate14008(.O (g32141), .I1 (g31639), .I2 (g29963));
AN2X1 gate14009(.O (g22316), .I1 (g2837), .I2 (g20270));
AN2X1 gate14010(.O (g18318), .I1 (g1604), .I2 (g17873));
AN2X1 gate14011(.O (g18446), .I1 (g2279), .I2 (g18008));
AN2X1 gate14012(.O (g33808), .I1 (g33109), .I2 (g22161));
AN2X1 gate14013(.O (g24785), .I1 (g7051), .I2 (g23645));
AN2X1 gate14014(.O (g18227), .I1 (g1052), .I2 (g16129));
AN3X1 gate14015(.O (g7777), .I1 (g723), .I2 (g822), .I3 (g817));
AN2X1 gate14016(.O (g27181), .I1 (g26026), .I2 (g16655));
AN2X1 gate14017(.O (g30209), .I1 (g28682), .I2 (g23876));
AN3X1 gate14018(.O (g22498), .I1 (g7753), .I2 (g7717), .I3 (g21334));
AN2X1 gate14019(.O (g33101), .I1 (g32398), .I2 (g18976));
AN2X1 gate14020(.O (g19791), .I1 (g14253), .I2 (g17189));
AN2X1 gate14021(.O (g24754), .I1 (g19604), .I2 (g23027));
AN2X1 gate14022(.O (g29595), .I1 (g28475), .I2 (g11833));
AN2X1 gate14023(.O (g29494), .I1 (g9073), .I2 (g28479));
AN2X1 gate14024(.O (g30208), .I1 (g28681), .I2 (g23875));
AN2X1 gate14025(.O (g16732), .I1 (g5555), .I2 (g14882));
AN2X1 gate14026(.O (g21929), .I1 (g5176), .I2 (g18997));
AN2X1 gate14027(.O (g32263), .I1 (g31631), .I2 (g30306));
AN2X1 gate14028(.O (g18540), .I1 (g2775), .I2 (g15277));
AN2X1 gate14029(.O (g10896), .I1 (g1205), .I2 (g8654));
AN2X1 gate14030(.O (g22056), .I1 (g6133), .I2 (g21611));
AN2X1 gate14031(.O (g26274), .I1 (g2130), .I2 (g25210));
AN2X1 gate14032(.O (g29623), .I1 (g28496), .I2 (g11563));
AN2X1 gate14033(.O (g32332), .I1 (g31325), .I2 (g23558));
AN4X1 gate14034(.O (I31206), .I1 (g31710), .I2 (g31832), .I3 (g32752), .I4 (g32753));
AN2X1 gate14035(.O (g21928), .I1 (g5170), .I2 (g18997));
AN2X1 gate14036(.O (g22080), .I1 (g6275), .I2 (g19210));
AN2X1 gate14037(.O (g25063), .I1 (g13078), .I2 (g22325));
AN3X1 gate14038(.O (g24858), .I1 (g3361), .I2 (g23223), .I3 (I24030));
AN2X1 gate14039(.O (g29782), .I1 (g28328), .I2 (g23245));
AN2X1 gate14040(.O (g18203), .I1 (g911), .I2 (g15938));
AN2X1 gate14041(.O (g26122), .I1 (g24557), .I2 (g19762));
AN2X1 gate14042(.O (g16761), .I1 (g7170), .I2 (g12947));
AN2X1 gate14043(.O (g29984), .I1 (g2567), .I2 (g28877));
AN2X1 gate14044(.O (g34542), .I1 (g34332), .I2 (g20089));
AN3X1 gate14045(.O (g22432), .I1 (g9354), .I2 (g7717), .I3 (g21187));
AN2X1 gate14046(.O (g12931), .I1 (g392), .I2 (g11048));
AN2X1 gate14047(.O (g29352), .I1 (g4950), .I2 (g28410));
AN2X1 gate14048(.O (g25873), .I1 (g24854), .I2 (g16197));
AN2X1 gate14049(.O (g30614), .I1 (g20154), .I2 (g29814));
AN3X1 gate14050(.O (I24597), .I1 (g5736), .I2 (g5742), .I3 (g9875));
AN4X1 gate14051(.O (I31082), .I1 (g32573), .I2 (g32574), .I3 (g32575), .I4 (g32576));
AN2X1 gate14052(.O (g18281), .I1 (g1373), .I2 (g16136));
AN2X1 gate14053(.O (g27520), .I1 (g26519), .I2 (g17714));
AN2X1 gate14054(.O (g21787), .I1 (g15091), .I2 (g20391));
AN2X1 gate14055(.O (g15115), .I1 (g2946), .I2 (g14454));
AN4X1 gate14056(.O (I31107), .I1 (g32610), .I2 (g32611), .I3 (g32612), .I4 (g32613));
AN3X1 gate14057(.O (g22342), .I1 (g9354), .I2 (g9285), .I3 (g21287));
AN2X1 gate14058(.O (g18301), .I1 (g1532), .I2 (g16489));
AN2X1 gate14059(.O (g30607), .I1 (g30291), .I2 (g18989));
AN2X1 gate14060(.O (g32049), .I1 (g10902), .I2 (g30735));
AN4X1 gate14061(.O (I24689), .I1 (g20841), .I2 (g24040), .I3 (g24041), .I4 (g24042));
AN2X1 gate14062(.O (g26292), .I1 (g2689), .I2 (g25228));
AN2X1 gate14063(.O (g33693), .I1 (g33145), .I2 (g13594));
AN2X1 gate14064(.O (g18377), .I1 (g1894), .I2 (g15171));
AN2X1 gate14065(.O (g19556), .I1 (g11932), .I2 (g16809));
AN2X1 gate14066(.O (g30073), .I1 (g1379), .I2 (g28194));
AN2X1 gate14067(.O (g22145), .I1 (g14555), .I2 (g18832));
AN2X1 gate14068(.O (g18120), .I1 (g457), .I2 (g17015));
AN2X1 gate14069(.O (g26153), .I1 (g24565), .I2 (g19780));
AN2X1 gate14070(.O (g18739), .I1 (g5008), .I2 (g16826));
AN2X1 gate14071(.O (g21302), .I1 (g956), .I2 (g15731));
AN2X1 gate14072(.O (g22031), .I1 (g5917), .I2 (g19147));
AN2X1 gate14073(.O (g27546), .I1 (g26549), .I2 (g17758));
AN2X1 gate14074(.O (g30274), .I1 (g28815), .I2 (g23983));
AN2X1 gate14075(.O (g31166), .I1 (g1816), .I2 (g30074));
AN2X1 gate14076(.O (g34073), .I1 (g8948), .I2 (g33823));
AN2X1 gate14077(.O (g10925), .I1 (g7858), .I2 (g956));
AN2X1 gate14078(.O (g16207), .I1 (g9839), .I2 (g14204));
AN2X1 gate14079(.O (g27211), .I1 (g25997), .I2 (g16716));
AN2X1 gate14080(.O (g32048), .I1 (g31498), .I2 (g13869));
AN4X1 gate14081(.O (g16539), .I1 (g11547), .I2 (g6782), .I3 (g6789), .I4 (I17741));
AN2X1 gate14082(.O (g21743), .I1 (g3100), .I2 (g20330));
AN2X1 gate14083(.O (g21827), .I1 (g3759), .I2 (g20453));
AN2X1 gate14084(.O (g11029), .I1 (g5782), .I2 (g9103));
AN2X1 gate14085(.O (g17753), .I1 (g13281), .I2 (g13175));
AN2X1 gate14086(.O (g18146), .I1 (g595), .I2 (g17533));
AN2X1 gate14087(.O (g18738), .I1 (g15142), .I2 (g16826));
AN2X1 gate14088(.O (g13029), .I1 (g8359), .I2 (g11030));
AN2X1 gate14089(.O (g15745), .I1 (g686), .I2 (g13223));
AN2X1 gate14090(.O (g18645), .I1 (g15100), .I2 (g17271));
AN2X1 gate14091(.O (g30122), .I1 (g28578), .I2 (g21054));
AN2X1 gate14092(.O (g24420), .I1 (g23997), .I2 (g18980));
AN2X1 gate14093(.O (g24319), .I1 (g4561), .I2 (g22228));
AN2X1 gate14094(.O (g29853), .I1 (g1862), .I2 (g29081));
AN2X1 gate14095(.O (g16538), .I1 (g6255), .I2 (g15005));
AN2X1 gate14096(.O (g17145), .I1 (g7469), .I2 (g13249));
AN2X1 gate14097(.O (g26635), .I1 (g25321), .I2 (g20617));
AN2X1 gate14098(.O (g11028), .I1 (g9730), .I2 (g5428));
AN2X1 gate14099(.O (g18699), .I1 (g4760), .I2 (g16816));
AN2X1 gate14100(.O (g34565), .I1 (g34374), .I2 (g17471));
AN2X1 gate14101(.O (g15813), .I1 (g3247), .I2 (g14069));
AN2X1 gate14102(.O (g31485), .I1 (g29776), .I2 (g23421));
AN2X1 gate14103(.O (g29589), .I1 (g2575), .I2 (g28977));
AN2X1 gate14104(.O (g33892), .I1 (g33312), .I2 (g20701));
AN2X1 gate14105(.O (g18290), .I1 (g1467), .I2 (g16449));
AN2X1 gate14106(.O (g17199), .I1 (g2236), .I2 (g13034));
AN2X1 gate14107(.O (g24318), .I1 (g4555), .I2 (g22228));
AN3X1 gate14108(.O (g33476), .I1 (g32570), .I2 (I31076), .I3 (I31077));
AN3X1 gate14109(.O (g33485), .I1 (g32635), .I2 (I31121), .I3 (I31122));
AN2X1 gate14110(.O (g21769), .I1 (g3247), .I2 (g20785));
AN2X1 gate14111(.O (g30034), .I1 (g29077), .I2 (g10541));
AN2X1 gate14112(.O (g22843), .I1 (g9429), .I2 (g20272));
AN2X1 gate14113(.O (g24227), .I1 (g890), .I2 (g22594));
AN2X1 gate14114(.O (g18698), .I1 (g15131), .I2 (g16777));
AN4X1 gate14115(.O (I31141), .I1 (g31376), .I2 (g31820), .I3 (g32659), .I4 (g32660));
AN3X1 gate14116(.O (g25453), .I1 (g5406), .I2 (g23789), .I3 (I24576));
AN2X1 gate14117(.O (g29588), .I1 (g2311), .I2 (g28942));
AN2X1 gate14118(.O (g29524), .I1 (g2004), .I2 (g28864));
AN2X1 gate14119(.O (g29836), .I1 (g28425), .I2 (g26841));
AN2X1 gate14120(.O (g21768), .I1 (g3243), .I2 (g20785));
AN2X1 gate14121(.O (g21803), .I1 (g3538), .I2 (g20924));
AN2X1 gate14122(.O (g28245), .I1 (g11367), .I2 (g27975));
AN2X1 gate14123(.O (g15805), .I1 (g3243), .I2 (g14041));
AN2X1 gate14124(.O (g28626), .I1 (g27542), .I2 (g20573));
AN2X1 gate14125(.O (g30153), .I1 (g28610), .I2 (g23768));
AN2X1 gate14126(.O (g28299), .I1 (g9716), .I2 (g27670));
AN4X1 gate14127(.O (g27700), .I1 (g22342), .I2 (g25182), .I3 (g26424), .I4 (g26148));
AN2X1 gate14128(.O (g22132), .I1 (g6645), .I2 (g19277));
AN2X1 gate14129(.O (g29477), .I1 (g14090), .I2 (g28441));
AN2X1 gate14130(.O (g32273), .I1 (g31255), .I2 (g20446));
AN2X1 gate14131(.O (g32106), .I1 (g31601), .I2 (g29911));
AN2X1 gate14132(.O (g18427), .I1 (g2181), .I2 (g18008));
AN2X1 gate14133(.O (g14681), .I1 (g4392), .I2 (g10476));
AN2X1 gate14134(.O (g19740), .I1 (g2783), .I2 (g15907));
AN2X1 gate14135(.O (g20203), .I1 (g6195), .I2 (g17789));
AN3X1 gate14136(.O (g33907), .I1 (g23088), .I2 (g33219), .I3 (g9104));
AN2X1 gate14137(.O (g18366), .I1 (g1854), .I2 (g17955));
AN4X1 gate14138(.O (I31332), .I1 (g32935), .I2 (g32936), .I3 (g32937), .I4 (g32938));
AN2X1 gate14139(.O (g21881), .I1 (g4064), .I2 (g19801));
AN2X1 gate14140(.O (g27658), .I1 (g22491), .I2 (g25786));
AN2X1 gate14141(.O (g18632), .I1 (g3698), .I2 (g17226));
AN2X1 gate14142(.O (g25905), .I1 (g24879), .I2 (g16311));
AN2X1 gate14143(.O (g17365), .I1 (g7650), .I2 (g13036));
AN2X1 gate14144(.O (g22161), .I1 (g13202), .I2 (g19071));
AN2X1 gate14145(.O (g33074), .I1 (g32387), .I2 (g18830));
AN2X1 gate14146(.O (g34136), .I1 (g33850), .I2 (g23293));
AN2X1 gate14147(.O (g33239), .I1 (g32117), .I2 (g19902));
AN2X1 gate14148(.O (g25530), .I1 (g23750), .I2 (g21414));
AN2X1 gate14149(.O (g27339), .I1 (g26400), .I2 (g17308));
AN2X1 gate14150(.O (g29749), .I1 (g28295), .I2 (g23214));
AN2X1 gate14151(.O (g29616), .I1 (g1974), .I2 (g29085));
AN3X1 gate14152(.O (g7511), .I1 (g2145), .I2 (g2138), .I3 (g2130));
AN2X1 gate14153(.O (g26711), .I1 (g25446), .I2 (g20713));
AN2X1 gate14154(.O (g31238), .I1 (g29583), .I2 (g20053));
AN2X1 gate14155(.O (g32234), .I1 (g31601), .I2 (g30292));
AN2X1 gate14156(.O (g25122), .I1 (g23374), .I2 (g20592));
AN2X1 gate14157(.O (g18403), .I1 (g2028), .I2 (g15373));
AN2X1 gate14158(.O (g18547), .I1 (g121), .I2 (g15277));
AN2X1 gate14159(.O (g25565), .I1 (g13013), .I2 (g22660));
AN2X1 gate14160(.O (g24301), .I1 (g6961), .I2 (g22228));
AN2X1 gate14161(.O (g28232), .I1 (g27732), .I2 (g23586));
AN2X1 gate14162(.O (g20739), .I1 (g16259), .I2 (g4674));
AN2X1 gate14163(.O (g13491), .I1 (g6999), .I2 (g12160));
AN2X1 gate14164(.O (g22087), .I1 (g6303), .I2 (g19210));
AN2X1 gate14165(.O (g30164), .I1 (g28618), .I2 (g23787));
AN2X1 gate14166(.O (g31941), .I1 (g1283), .I2 (g30825));
AN2X1 gate14167(.O (g33941), .I1 (g33380), .I2 (g21560));
AN2X1 gate14168(.O (g18226), .I1 (g15064), .I2 (g16129));
AN2X1 gate14169(.O (g21890), .I1 (g4125), .I2 (g19801));
AN2X1 gate14170(.O (g13604), .I1 (g4495), .I2 (g10487));
AN2X1 gate14171(.O (g31519), .I1 (g29864), .I2 (g23490));
AN2X1 gate14172(.O (g18715), .I1 (g4871), .I2 (g15915));
AN2X1 gate14173(.O (g27968), .I1 (g25958), .I2 (g19614));
AN2X1 gate14174(.O (g28697), .I1 (g27581), .I2 (g20669));
AN2X1 gate14175(.O (g31185), .I1 (g10114), .I2 (g30087));
AN2X1 gate14176(.O (g18481), .I1 (g2461), .I2 (g15426));
AN3X1 gate14177(.O (g33519), .I1 (g32881), .I2 (I31291), .I3 (I31292));
AN2X1 gate14178(.O (g29809), .I1 (g28362), .I2 (g23274));
AN3X1 gate14179(.O (g33675), .I1 (g33164), .I2 (g10727), .I3 (g22332));
AN2X1 gate14180(.O (g24645), .I1 (g22639), .I2 (g19709));
AN2X1 gate14181(.O (g28261), .I1 (g27878), .I2 (g23695));
AN2X1 gate14182(.O (g26606), .I1 (g1018), .I2 (g24510));
AN4X1 gate14183(.O (g28880), .I1 (g21434), .I2 (g26424), .I3 (g25438), .I4 (g27494));
AN2X1 gate14184(.O (g18551), .I1 (g2811), .I2 (g15277));
AN2X1 gate14185(.O (g22043), .I1 (g5965), .I2 (g19147));
AN2X1 gate14186(.O (g26303), .I1 (g2685), .I2 (g25439));
AN2X1 gate14187(.O (g31518), .I1 (g20041), .I2 (g29970));
AN2X1 gate14188(.O (g31154), .I1 (g19128), .I2 (g29814));
AN2X1 gate14189(.O (g18572), .I1 (g2864), .I2 (g16349));
AN3X1 gate14190(.O (g33518), .I1 (g32874), .I2 (I31286), .I3 (I31287));
AN2X1 gate14191(.O (g29808), .I1 (g28361), .I2 (g23273));
AN2X1 gate14192(.O (g21710), .I1 (g287), .I2 (g20283));
AN4X1 gate14193(.O (I31221), .I1 (g31327), .I2 (g31835), .I3 (g32773), .I4 (g32774));
AN2X1 gate14194(.O (g24290), .I1 (g4430), .I2 (g22550));
AN4X1 gate14195(.O (g29036), .I1 (g27163), .I2 (g12762), .I3 (g20875), .I4 (I27381));
AN2X1 gate14196(.O (g27411), .I1 (g26549), .I2 (g17528));
AN2X1 gate14197(.O (g34474), .I1 (g20083), .I2 (g34326));
AN2X1 gate14198(.O (g24698), .I1 (g22664), .I2 (g19761));
AN2X1 gate14199(.O (g21779), .I1 (g3385), .I2 (g20391));
AN2X1 gate14200(.O (g26750), .I1 (g24514), .I2 (g24474));
AN2X1 gate14201(.O (g12527), .I1 (g8680), .I2 (g667));
AN2X1 gate14202(.O (g23779), .I1 (g1105), .I2 (g19355));
AN2X1 gate14203(.O (g18127), .I1 (g499), .I2 (g16971));
AN2X1 gate14204(.O (g22069), .I1 (g6227), .I2 (g19210));
AN2X1 gate14205(.O (g25408), .I1 (g22682), .I2 (g9772));
AN2X1 gate14206(.O (g30109), .I1 (g28562), .I2 (g20912));
AN2X1 gate14207(.O (g26381), .I1 (g4456), .I2 (g25548));
AN2X1 gate14208(.O (g34109), .I1 (g33918), .I2 (g23708));
AN2X1 gate14209(.O (g29642), .I1 (g27954), .I2 (g28669));
AN2X1 gate14210(.O (g33883), .I1 (g33294), .I2 (g20589));
AN2X1 gate14211(.O (g21778), .I1 (g3355), .I2 (g20391));
AN2X1 gate14212(.O (g22068), .I1 (g6219), .I2 (g19210));
AN2X1 gate14213(.O (g26091), .I1 (g1691), .I2 (g25082));
AN2X1 gate14214(.O (g18490), .I1 (g2504), .I2 (g15426));
AN2X1 gate14215(.O (g30108), .I1 (g28561), .I2 (g20910));
AN2X1 gate14216(.O (g32163), .I1 (g3502), .I2 (g31170));
AN2X1 gate14217(.O (g32012), .I1 (g8297), .I2 (g31233));
AN3X1 gate14218(.O (g34108), .I1 (g22957), .I2 (g9104), .I3 (g33766));
AN2X1 gate14219(.O (g24427), .I1 (g4961), .I2 (g22919));
AN2X1 gate14220(.O (g21786), .I1 (g3436), .I2 (g20391));
AN2X1 gate14221(.O (g27503), .I1 (g26488), .I2 (g14668));
AN3X1 gate14222(.O (I24054), .I1 (g8443), .I2 (g8075), .I3 (g3747));
AN2X1 gate14223(.O (g30283), .I1 (g28851), .I2 (g23993));
AN4X1 gate14224(.O (I31106), .I1 (g30825), .I2 (g31814), .I3 (g32608), .I4 (g32609));
AN2X1 gate14225(.O (g18784), .I1 (g15155), .I2 (g18065));
AN2X1 gate14226(.O (g18376), .I1 (g1913), .I2 (g15171));
AN2X1 gate14227(.O (g18385), .I1 (g1959), .I2 (g15171));
AN2X1 gate14228(.O (g29733), .I1 (g2675), .I2 (g29157));
AN2X1 gate14229(.O (g18297), .I1 (g1478), .I2 (g16449));
AN2X1 gate14230(.O (g17810), .I1 (g1495), .I2 (g13246));
AN2X1 gate14231(.O (g18103), .I1 (g401), .I2 (g17015));
AN2X1 gate14232(.O (g10626), .I1 (g4057), .I2 (g7927));
AN2X1 gate14233(.O (g34492), .I1 (g34272), .I2 (g33430));
AN2X1 gate14234(.O (g13633), .I1 (g4567), .I2 (g10509));
AN2X1 gate14235(.O (g25164), .I1 (g16883), .I2 (g23569));
AN2X1 gate14236(.O (g21945), .I1 (g5248), .I2 (g18997));
AN2X1 gate14237(.O (g28499), .I1 (g27982), .I2 (g17762));
AN2X1 gate14238(.O (g18354), .I1 (g1792), .I2 (g17955));
AN2X1 gate14239(.O (g29874), .I1 (g28402), .I2 (g23336));
AN4X1 gate14240(.O (g27714), .I1 (g22384), .I2 (g25195), .I3 (g26424), .I4 (g26171));
AN2X1 gate14241(.O (g21826), .I1 (g3742), .I2 (g20453));
AN2X1 gate14242(.O (g21999), .I1 (g5723), .I2 (g21562));
AN2X1 gate14243(.O (g26390), .I1 (g4423), .I2 (g25554));
AN2X1 gate14244(.O (g31501), .I1 (g2047), .I2 (g29310));
AN2X1 gate14245(.O (g18824), .I1 (g6732), .I2 (g15680));
AN2X1 gate14246(.O (g27315), .I1 (g12022), .I2 (g26709));
AN3X1 gate14247(.O (g33501), .I1 (g32751), .I2 (I31201), .I3 (I31202));
AN2X1 gate14248(.O (g29630), .I1 (g28212), .I2 (g19781));
AN2X1 gate14249(.O (g24403), .I1 (g4894), .I2 (g22858));
AN2X1 gate14250(.O (g29693), .I1 (g28207), .I2 (g10233));
AN2X1 gate14251(.O (g30982), .I1 (g8895), .I2 (g29933));
AN2X1 gate14252(.O (g34750), .I1 (g34673), .I2 (g19542));
AN2X1 gate14253(.O (g16759), .I1 (g5587), .I2 (g14761));
AN2X1 gate14254(.O (g18181), .I1 (g772), .I2 (g17328));
AN2X1 gate14255(.O (g21998), .I1 (g5712), .I2 (g21562));
AN2X1 gate14256(.O (g18671), .I1 (g4628), .I2 (g15758));
AN2X1 gate14257(.O (g34381), .I1 (g34166), .I2 (g20594));
AN2X1 gate14258(.O (g23998), .I1 (g19631), .I2 (g10971));
AN3X1 gate14259(.O (g33728), .I1 (g22626), .I2 (g10851), .I3 (g33187));
AN2X1 gate14260(.O (g27202), .I1 (g25997), .I2 (g13876));
AN2X1 gate14261(.O (g19568), .I1 (g1467), .I2 (g15959));
AN2X1 gate14262(.O (g30091), .I1 (g28127), .I2 (g20716));
AN2X1 gate14263(.O (g32325), .I1 (g31316), .I2 (g23538));
AN2X1 gate14264(.O (g29665), .I1 (g2375), .I2 (g28696));
AN2X1 gate14265(.O (g16758), .I1 (g5220), .I2 (g14758));
AN3X1 gate14266(.O (g34091), .I1 (g22957), .I2 (g9104), .I3 (g33761));
AN2X1 gate14267(.O (g24226), .I1 (g446), .I2 (g22594));
AN2X1 gate14268(.O (g13832), .I1 (g8880), .I2 (g10612));
AN2X1 gate14269(.O (g28722), .I1 (g27955), .I2 (g20738));
AN4X1 gate14270(.O (g28924), .I1 (g17317), .I2 (g25183), .I3 (g26424), .I4 (g27416));
AN2X1 gate14271(.O (g30174), .I1 (g28628), .I2 (g23812));
AN4X1 gate14272(.O (g29008), .I1 (g27163), .I2 (g12730), .I3 (g20739), .I4 (I27364));
AN2X1 gate14273(.O (g12979), .I1 (g424), .I2 (g11048));
AN2X1 gate14274(.O (g24551), .I1 (g17148), .I2 (g23331));
AN2X1 gate14275(.O (g24572), .I1 (g5462), .I2 (g23393));
AN2X1 gate14276(.O (g33349), .I1 (g32233), .I2 (g20699));
AN2X1 gate14277(.O (g25108), .I1 (g23345), .I2 (g20576));
AN2X1 gate14278(.O (g21932), .I1 (g5204), .I2 (g18997));
AN2X1 gate14279(.O (g32121), .I1 (g31616), .I2 (g29942));
AN2X1 gate14280(.O (g18426), .I1 (g2177), .I2 (g18008));
AN2X1 gate14281(.O (g33906), .I1 (g33084), .I2 (g22311));
AN2X1 gate14282(.O (g13247), .I1 (g8964), .I2 (g11316));
AN2X1 gate14283(.O (g29555), .I1 (g29004), .I2 (g22498));
AN2X1 gate14284(.O (g21513), .I1 (g16196), .I2 (g10882));
AN2X1 gate14285(.O (g18190), .I1 (g822), .I2 (g17821));
AN2X1 gate14286(.O (g22010), .I1 (g5787), .I2 (g21562));
AN2X1 gate14287(.O (g23513), .I1 (g19430), .I2 (g13007));
AN2X1 gate14288(.O (g34390), .I1 (g34172), .I2 (g21069));
AN2X1 gate14289(.O (g10856), .I1 (g4269), .I2 (g8967));
AN2X1 gate14290(.O (g11045), .I1 (g5787), .I2 (g9883));
AN2X1 gate14291(.O (g15882), .I1 (g3554), .I2 (g13986));
AN2X1 gate14292(.O (g27384), .I1 (g26400), .I2 (g17496));
AN2X1 gate14293(.O (g29570), .I1 (g2763), .I2 (g28598));
AN2X1 gate14294(.O (g29712), .I1 (g2643), .I2 (g28726));
AN4X1 gate14295(.O (I24694), .I1 (g20982), .I2 (g24047), .I3 (g24048), .I4 (g24049));
AN2X1 gate14296(.O (g33304), .I1 (g32427), .I2 (g31971));
AN2X1 gate14297(.O (g14261), .I1 (g4507), .I2 (g10738));
AN2X1 gate14298(.O (g18520), .I1 (g2661), .I2 (g15509));
AN2X1 gate14299(.O (g21961), .I1 (g5424), .I2 (g21514));
AN2X1 gate14300(.O (g22079), .I1 (g6271), .I2 (g19210));
AN2X1 gate14301(.O (g27094), .I1 (g25997), .I2 (g16472));
AN2X1 gate14302(.O (g30192), .I1 (g28649), .I2 (g23847));
AN2X1 gate14303(.O (g31566), .I1 (g19050), .I2 (g29814));
AN2X1 gate14304(.O (g13324), .I1 (g854), .I2 (g11326));
AN2X1 gate14305(.O (g29907), .I1 (g2629), .I2 (g29177));
AN2X1 gate14306(.O (g32291), .I1 (g31268), .I2 (g20527));
AN2X1 gate14307(.O (g16804), .I1 (g5905), .I2 (g14813));
AN2X1 gate14308(.O (g21404), .I1 (g16069), .I2 (g13569));
AN2X1 gate14309(.O (g28199), .I1 (g27479), .I2 (g16684));
AN2X1 gate14310(.O (g22078), .I1 (g6267), .I2 (g19210));
AN2X1 gate14311(.O (g23404), .I1 (g20063), .I2 (g20247));
AN2X1 gate14312(.O (g32173), .I1 (g160), .I2 (g31134));
AN2X1 gate14313(.O (g18546), .I1 (g2795), .I2 (g15277));
AN2X1 gate14314(.O (g25982), .I1 (g2351), .I2 (g25008));
AN4X1 gate14315(.O (I31012), .I1 (g32473), .I2 (g32474), .I3 (g32475), .I4 (g32476));
AN2X1 gate14316(.O (g18211), .I1 (g15062), .I2 (g15979));
AN2X1 gate14317(.O (g21717), .I1 (g15051), .I2 (g21037));
AN2X1 gate14318(.O (g28198), .I1 (g26649), .I2 (g27492));
AN2X1 gate14319(.O (g24297), .I1 (g4455), .I2 (g22550));
AN2X1 gate14320(.O (g22086), .I1 (g6299), .I2 (g19210));
AN2X1 gate14321(.O (g25091), .I1 (g12830), .I2 (g23492));
AN2X1 gate14322(.O (g20095), .I1 (g8873), .I2 (g16632));
AN3X1 gate14323(.O (I24619), .I1 (g6423), .I2 (g6428), .I3 (g10014));
AN2X1 gate14324(.O (g29567), .I1 (g2357), .I2 (g28593));
AN2X1 gate14325(.O (g29594), .I1 (g28529), .I2 (g14192));
AN3X1 gate14326(.O (g12735), .I1 (g7121), .I2 (g3873), .I3 (g3881));
AN2X1 gate14327(.O (g31139), .I1 (g12221), .I2 (g30036));
AN2X1 gate14328(.O (g28528), .I1 (g27187), .I2 (g12730));
AN2X1 gate14329(.O (g28330), .I1 (g27238), .I2 (g19786));
AN2X1 gate14330(.O (g26252), .I1 (g2283), .I2 (g25309));
AN2X1 gate14331(.O (g11032), .I1 (g9354), .I2 (g7717));
AN2X1 gate14332(.O (g34483), .I1 (g34406), .I2 (g18938));
AN2X1 gate14333(.O (g18497), .I1 (g2541), .I2 (g15426));
AN2X1 gate14334(.O (g32029), .I1 (g31318), .I2 (g16482));
AN2X1 gate14335(.O (g24671), .I1 (g5481), .I2 (g23630));
AN2X1 gate14336(.O (g14831), .I1 (g1152), .I2 (g10909));
AN2X1 gate14337(.O (g22125), .I1 (g6617), .I2 (g19277));
AN3X1 gate14338(.O (g29382), .I1 (g26424), .I2 (g22763), .I3 (g28172));
AN2X1 gate14339(.O (g27526), .I1 (g26576), .I2 (g17721));
AN2X1 gate14340(.O (g34862), .I1 (g16540), .I2 (g34830));
AN2X1 gate14341(.O (g29519), .I1 (g2295), .I2 (g28840));
AN2X1 gate14342(.O (g32028), .I1 (g30569), .I2 (g29339));
AN2X1 gate14343(.O (g19578), .I1 (g16183), .I2 (g11130));
AN2X1 gate14344(.O (g33415), .I1 (g32368), .I2 (g21422));
AN2X1 gate14345(.O (g22158), .I1 (g13698), .I2 (g19609));
AN2X1 gate14346(.O (g14316), .I1 (g2370), .I2 (g11920));
AN2X1 gate14347(.O (g33333), .I1 (g32218), .I2 (g20612));
AN2X1 gate14348(.O (g18700), .I1 (g15132), .I2 (g16816));
AN4X1 gate14349(.O (g17817), .I1 (g11547), .I2 (g6782), .I3 (g11640), .I4 (I18819));
AN2X1 gate14350(.O (g18126), .I1 (g15054), .I2 (g16971));
AN2X1 gate14351(.O (g18659), .I1 (g4366), .I2 (g17183));
AN2X1 gate14352(.O (g18625), .I1 (g15092), .I2 (g17062));
AN2X1 gate14353(.O (g18987), .I1 (g182), .I2 (g16162));
AN2X1 gate14354(.O (g29518), .I1 (g28906), .I2 (g22384));
AN2X1 gate14355(.O (g18250), .I1 (g6821), .I2 (g16897));
AN2X1 gate14356(.O (g24931), .I1 (g23153), .I2 (g20178));
AN2X1 gate14357(.O (g15114), .I1 (g4239), .I2 (g14454));
AN2X1 gate14358(.O (g25192), .I1 (g20276), .I2 (g23648));
AN2X1 gate14359(.O (g26847), .I1 (g2873), .I2 (g24525));
AN2X1 gate14360(.O (g34948), .I1 (g16540), .I2 (g34935));
AN2X1 gate14361(.O (g18658), .I1 (g15121), .I2 (g17183));
AN2X1 gate14362(.O (g27457), .I1 (g26519), .I2 (g17606));
AN2X1 gate14363(.O (g26397), .I1 (g19475), .I2 (g25563));
AN2X1 gate14364(.O (g15082), .I1 (g2697), .I2 (g12983));
AN2X1 gate14365(.O (g23387), .I1 (g16506), .I2 (g20211));
AN2X1 gate14366(.O (g31963), .I1 (g30731), .I2 (g18895));
AN2X1 gate14367(.O (g29637), .I1 (g2533), .I2 (g29134));
AN2X1 gate14368(.O (g22680), .I1 (g19530), .I2 (g7781));
AN2X1 gate14369(.O (g34702), .I1 (g34537), .I2 (g20208));
AN2X1 gate14370(.O (g15107), .I1 (g4258), .I2 (g14454));
AN2X1 gate14371(.O (g23148), .I1 (g19128), .I2 (g9104));
AN2X1 gate14372(.O (g34757), .I1 (g34682), .I2 (g19635));
AN2X1 gate14373(.O (g17783), .I1 (g7851), .I2 (g13110));
AN2X1 gate14374(.O (g25522), .I1 (g6888), .I2 (g22544));
AN4X1 gate14375(.O (I31121), .I1 (g30614), .I2 (g31817), .I3 (g32629), .I4 (g32630));
AN2X1 gate14376(.O (g24190), .I1 (g329), .I2 (g22722));
AN2X1 gate14377(.O (g18339), .I1 (g1714), .I2 (g17873));
AN2X1 gate14378(.O (g18943), .I1 (g269), .I2 (g16099));
AN2X1 gate14379(.O (g29883), .I1 (g2465), .I2 (g29152));
AN2X1 gate14380(.O (g18296), .I1 (g1495), .I2 (g16449));
AN2X1 gate14381(.O (g21811), .I1 (g3582), .I2 (g20924));
AN2X1 gate14382(.O (g28225), .I1 (g27770), .I2 (g23400));
AN2X1 gate14383(.O (g23104), .I1 (g661), .I2 (g20248));
AN2X1 gate14384(.O (g23811), .I1 (g4087), .I2 (g19364));
AN2X1 gate14385(.O (g23646), .I1 (g16959), .I2 (g20737));
AN2X1 gate14386(.O (g18644), .I1 (g15098), .I2 (g17125));
AN4X1 gate14387(.O (g28471), .I1 (g27187), .I2 (g12762), .I3 (g21024), .I4 (I26960));
AN2X1 gate14388(.O (g16221), .I1 (g5791), .I2 (g14231));
AN2X1 gate14389(.O (g18338), .I1 (g1710), .I2 (g17873));
AN2X1 gate14390(.O (g30564), .I1 (g21358), .I2 (g29385));
AN2X1 gate14391(.O (g9967), .I1 (g1178), .I2 (g1157));
AN2X1 gate14392(.O (g28258), .I1 (g27182), .I2 (g19687));
AN2X1 gate14393(.O (g21971), .I1 (g5417), .I2 (g21514));
AN2X1 gate14394(.O (g34564), .I1 (g34373), .I2 (g17466));
AN2X1 gate14395(.O (g15849), .I1 (g3538), .I2 (g14136));
AN2X1 gate14396(.O (g31484), .I1 (g29775), .I2 (g23418));
AN2X1 gate14397(.O (g24546), .I1 (g22447), .I2 (g19523));
AN3X1 gate14398(.O (g33484), .I1 (g32628), .I2 (I31116), .I3 (I31117));
AN2X1 gate14399(.O (g16613), .I1 (g5925), .I2 (g14732));
AN4X1 gate14400(.O (I31291), .I1 (g31021), .I2 (g31847), .I3 (g32875), .I4 (g32876));
AN2X1 gate14401(.O (g15848), .I1 (g3259), .I2 (g13892));
AN2X1 gate14402(.O (g19275), .I1 (g7823), .I2 (g16044));
AN2X1 gate14403(.O (g31554), .I1 (g19050), .I2 (g29814));
AN2X1 gate14404(.O (g30673), .I1 (g20175), .I2 (g29814));
AN2X1 gate14405(.O (g27256), .I1 (g25937), .I2 (g19698));
AN2X1 gate14406(.O (g19746), .I1 (g9816), .I2 (g17147));
AN2X1 gate14407(.O (g28244), .I1 (g27926), .I2 (g26715));
AN2X1 gate14408(.O (g34183), .I1 (g33695), .I2 (g24385));
AN2X1 gate14409(.O (g18197), .I1 (g854), .I2 (g17821));
AN2X1 gate14410(.O (g22017), .I1 (g5763), .I2 (g21562));
AN2X1 gate14411(.O (g15652), .I1 (g174), .I2 (g13437));
AN2X1 gate14412(.O (g15804), .I1 (g3223), .I2 (g13889));
AN2X1 gate14413(.O (g34397), .I1 (g7673), .I2 (g34068));
AN2X1 gate14414(.O (g25949), .I1 (g24701), .I2 (g19559));
AN2X1 gate14415(.O (g27280), .I1 (g9825), .I2 (g26614));
AN2X1 gate14416(.O (g31312), .I1 (g30136), .I2 (g27858));
AN2X1 gate14417(.O (g29577), .I1 (g2441), .I2 (g28946));
AN2X1 gate14418(.O (g30062), .I1 (g13129), .I2 (g28174));
AN2X1 gate14419(.O (g27300), .I1 (g12370), .I2 (g26672));
AN2X1 gate14420(.O (g10736), .I1 (g4040), .I2 (g8751));
AN3X1 gate14421(.O (g10887), .I1 (g7812), .I2 (g6565), .I3 (g6573));
AN2X1 gate14422(.O (g31115), .I1 (g29487), .I2 (g22882));
AN2X1 gate14423(.O (g18411), .I1 (g2093), .I2 (g15373));
AN2X1 gate14424(.O (g25536), .I1 (g23770), .I2 (g21431));
AN2X1 gate14425(.O (g25040), .I1 (g12738), .I2 (g23443));
AN4X1 gate14426(.O (g26213), .I1 (g25357), .I2 (g11724), .I3 (g7586), .I4 (g7558));
AN2X1 gate14427(.O (g34509), .I1 (g34283), .I2 (g19473));
AN2X1 gate14428(.O (g21850), .I1 (g3893), .I2 (g21070));
AN2X1 gate14429(.O (g28602), .I1 (g27509), .I2 (g20515));
AN2X1 gate14430(.O (g23412), .I1 (g7297), .I2 (g21510));
AN2X1 gate14431(.O (g28657), .I1 (g27562), .I2 (g20606));
AN2X1 gate14432(.O (g25904), .I1 (g14001), .I2 (g24791));
AN3X1 gate14433(.O (g33921), .I1 (g33187), .I2 (g9104), .I3 (g19200));
AN2X1 gate14434(.O (g19684), .I1 (g2735), .I2 (g17297));
AN2X1 gate14435(.O (g34508), .I1 (g34282), .I2 (g19472));
AN2X1 gate14436(.O (g10528), .I1 (g1576), .I2 (g9051));
AN2X1 gate14437(.O (g34872), .I1 (g34827), .I2 (g19954));
AN3X1 gate14438(.O (I18740), .I1 (g13156), .I2 (g11450), .I3 (g11498));
AN2X1 gate14439(.O (g24700), .I1 (g645), .I2 (g23512));
AN4X1 gate14440(.O (g28970), .I1 (g17405), .I2 (g25196), .I3 (g26424), .I4 (g27445));
AN2X1 gate14441(.O (g24659), .I1 (g5134), .I2 (g23590));
AN4X1 gate14442(.O (g14528), .I1 (g12459), .I2 (g12306), .I3 (g12245), .I4 (I16646));
AN2X1 gate14443(.O (g26205), .I1 (g2098), .I2 (g25492));
AN2X1 gate14444(.O (g23229), .I1 (g18994), .I2 (g4521));
AN4X1 gate14445(.O (g16234), .I1 (g6772), .I2 (g6782), .I3 (g11640), .I4 (I17575));
AN2X1 gate14446(.O (g29349), .I1 (g4760), .I2 (g28391));
AN2X1 gate14447(.O (g22309), .I1 (g1478), .I2 (g19751));
AN2X1 gate14448(.O (g20658), .I1 (g1389), .I2 (g15800));
AN2X1 gate14449(.O (g18503), .I1 (g2563), .I2 (g15509));
AN2X1 gate14450(.O (g22023), .I1 (g5881), .I2 (g19147));
AN2X1 gate14451(.O (g26311), .I1 (g2527), .I2 (g25400));
AN2X1 gate14452(.O (g24658), .I1 (g22645), .I2 (g19732));
AN3X1 gate14453(.O (I24015), .I1 (g8334), .I2 (g7975), .I3 (g3045));
AN3X1 gate14454(.O (g10869), .I1 (g7766), .I2 (g5873), .I3 (g5881));
AN2X1 gate14455(.O (g22308), .I1 (g1135), .I2 (g19738));
AN2X1 gate14456(.O (g28171), .I1 (g27016), .I2 (g19385));
AN2X1 gate14457(.O (g33798), .I1 (g33227), .I2 (g20058));
AN2X1 gate14458(.O (g21716), .I1 (g301), .I2 (g20283));
AN2X1 gate14459(.O (g30213), .I1 (g28688), .I2 (g23880));
AN2X1 gate14460(.O (g24296), .I1 (g4382), .I2 (g22550));
AN2X1 gate14461(.O (g18581), .I1 (g2912), .I2 (g16349));
AN2X1 gate14462(.O (g18714), .I1 (g4864), .I2 (g15915));
AN2X1 gate14463(.O (g26051), .I1 (g24896), .I2 (g14169));
AN2X1 gate14464(.O (g18450), .I1 (g2299), .I2 (g15224));
AN2X1 gate14465(.O (g31184), .I1 (g1950), .I2 (g30085));
AN2X1 gate14466(.O (g34213), .I1 (g33766), .I2 (g22689));
AN2X1 gate14467(.O (g18315), .I1 (g1548), .I2 (g16931));
AN2X1 gate14468(.O (g33805), .I1 (g33232), .I2 (g20079));
AN3X1 gate14469(.O (g33674), .I1 (g33164), .I2 (g10710), .I3 (g22319));
AN2X1 gate14470(.O (g24644), .I1 (g11714), .I2 (g22903));
AN2X1 gate14471(.O (g29622), .I1 (g2579), .I2 (g29001));
AN2X1 gate14472(.O (g29566), .I1 (g2307), .I2 (g28907));
AN2X1 gate14473(.O (g18707), .I1 (g15134), .I2 (g16782));
AN2X1 gate14474(.O (g18819), .I1 (g6541), .I2 (g15483));
AN2X1 gate14475(.O (g18910), .I1 (g16227), .I2 (g16075));
AN2X1 gate14476(.O (g18202), .I1 (g907), .I2 (g15938));
AN2X1 gate14477(.O (g30047), .I1 (g29109), .I2 (g9407));
AN2X1 gate14478(.O (g18257), .I1 (g1205), .I2 (g16897));
AN2X1 gate14479(.O (g26780), .I1 (g4098), .I2 (g24437));
AN2X1 gate14480(.O (g30205), .I1 (g28671), .I2 (g23869));
AN2X1 gate14481(.O (g32191), .I1 (g27593), .I2 (g31376));
AN2X1 gate14482(.O (g18818), .I1 (g15165), .I2 (g15483));
AN2X1 gate14483(.O (g18496), .I1 (g2537), .I2 (g15426));
AN2X1 gate14484(.O (g34205), .I1 (g33729), .I2 (g24541));
AN2X1 gate14485(.O (g31934), .I1 (g31670), .I2 (g18827));
AN2X1 gate14486(.O (g18111), .I1 (g174), .I2 (g17015));
AN2X1 gate14487(.O (g21959), .I1 (g5413), .I2 (g21514));
AN2X1 gate14488(.O (g21925), .I1 (g5073), .I2 (g21468));
AN2X1 gate14489(.O (g26350), .I1 (g13087), .I2 (g25517));
AN2X1 gate14490(.O (g25872), .I1 (g3119), .I2 (g24655));
AN2X1 gate14491(.O (g28919), .I1 (g27663), .I2 (g21295));
AN2X1 gate14492(.O (g14708), .I1 (g74), .I2 (g12369));
AN3X1 gate14493(.O (I18762), .I1 (g13156), .I2 (g6767), .I3 (g11498));
AN4X1 gate14494(.O (g28458), .I1 (g27187), .I2 (g12730), .I3 (g20887), .I4 (I26948));
AN2X1 gate14495(.O (g24197), .I1 (g347), .I2 (g22722));
AN3X1 gate14496(.O (g24855), .I1 (g3050), .I2 (g23534), .I3 (I24027));
AN3X1 gate14497(.O (g27660), .I1 (g24688), .I2 (g26424), .I3 (g22763));
AN2X1 gate14498(.O (g16163), .I1 (g14254), .I2 (g14179));
AN2X1 gate14499(.O (g22752), .I1 (g15792), .I2 (g19612));
AN2X1 gate14500(.O (g15613), .I1 (g3490), .I2 (g13555));
AN2X1 gate14501(.O (g18590), .I1 (g2917), .I2 (g16349));
AN2X1 gate14502(.O (g21958), .I1 (g5396), .I2 (g21514));
AN2X1 gate14503(.O (g21378), .I1 (g7887), .I2 (g16090));
AN2X1 gate14504(.O (g23050), .I1 (g655), .I2 (g20248));
AN4X1 gate14505(.O (g28010), .I1 (g23032), .I2 (g26223), .I3 (g26424), .I4 (g25535));
AN2X1 gate14506(.O (g23958), .I1 (g9104), .I2 (g19200));
AN2X1 gate14507(.O (g24411), .I1 (g4584), .I2 (g22161));
AN2X1 gate14508(.O (g30051), .I1 (g28513), .I2 (g20604));
AN2X1 gate14509(.O (g26846), .I1 (g37), .I2 (g24524));
AN2X1 gate14510(.O (g18741), .I1 (g15143), .I2 (g17384));
AN2X1 gate14511(.O (g34072), .I1 (g33839), .I2 (g24872));
AN2X1 gate14512(.O (g23386), .I1 (g20034), .I2 (g20207));
AN2X1 gate14513(.O (g30592), .I1 (g30270), .I2 (g18929));
AN2X1 gate14514(.O (g18384), .I1 (g1945), .I2 (g15171));
AN2X1 gate14515(.O (g29636), .I1 (g2403), .I2 (g29097));
AN2X1 gate14516(.O (g21742), .I1 (g3050), .I2 (g20330));
AN2X1 gate14517(.O (g17752), .I1 (g7841), .I2 (g13174));
AN2X1 gate14518(.O (g27480), .I1 (g26400), .I2 (g17638));
AN2X1 gate14519(.O (g34756), .I1 (g34680), .I2 (g19618));
AN2X1 gate14520(.O (g23742), .I1 (g19128), .I2 (g9104));
AN2X1 gate14521(.O (g28599), .I1 (g27027), .I2 (g8922));
AN2X1 gate14522(.O (g21944), .I1 (g5244), .I2 (g18997));
AN2X1 gate14523(.O (g33400), .I1 (g32347), .I2 (g21380));
AN2X1 gate14524(.O (g29852), .I1 (g1772), .I2 (g29080));
AN2X1 gate14525(.O (g17643), .I1 (g9681), .I2 (g14599));
AN2X1 gate14526(.O (g15812), .I1 (g3227), .I2 (g13915));
AN4X1 gate14527(.O (g13319), .I1 (g4076), .I2 (g8812), .I3 (g10658), .I4 (g8757));
AN2X1 gate14528(.O (g27314), .I1 (g12436), .I2 (g26702));
AN2X1 gate14529(.O (g24503), .I1 (g22225), .I2 (g19409));
AN2X1 gate14530(.O (g27287), .I1 (g26545), .I2 (g23011));
AN2X1 gate14531(.O (g32045), .I1 (g31491), .I2 (g16187));
AN4X1 gate14532(.O (I24685), .I1 (g24036), .I2 (g24037), .I3 (g24038), .I4 (g24039));
AN2X1 gate14533(.O (g33329), .I1 (g32210), .I2 (g20585));
AN2X1 gate14534(.O (g31207), .I1 (g30252), .I2 (g20739));
AN2X1 gate14535(.O (g18150), .I1 (g604), .I2 (g17533));
AN2X1 gate14536(.O (g10657), .I1 (g8451), .I2 (g4064));
AN2X1 gate14537(.O (g18801), .I1 (g15160), .I2 (g15348));
AN2X1 gate14538(.O (g18735), .I1 (g4983), .I2 (g16826));
AN2X1 gate14539(.O (g25574), .I1 (I24709), .I2 (I24710));
AN2X1 gate14540(.O (g27085), .I1 (g25835), .I2 (g22494));
AN2X1 gate14541(.O (g32324), .I1 (g31315), .I2 (g23537));
AN2X1 gate14542(.O (g29664), .I1 (g2273), .I2 (g29060));
AN2X1 gate14543(.O (g33328), .I1 (g32209), .I2 (g20584));
AN2X1 gate14544(.O (g21802), .I1 (g3562), .I2 (g20924));
AN2X1 gate14545(.O (g22489), .I1 (g12954), .I2 (g19386));
AN2X1 gate14546(.O (g21857), .I1 (g3933), .I2 (g21070));
AN2X1 gate14547(.O (g23802), .I1 (g9104), .I2 (g19050));
AN2X1 gate14548(.O (g16535), .I1 (g5595), .I2 (g14848));
AN2X1 gate14549(.O (g20581), .I1 (g10801), .I2 (g15571));
AN2X1 gate14550(.O (g10970), .I1 (g854), .I2 (g9582));
AN2X1 gate14551(.O (g23857), .I1 (g19626), .I2 (g7908));
AN2X1 gate14552(.O (g13059), .I1 (g6900), .I2 (g11303));
AN2X1 gate14553(.O (g13025), .I1 (g8431), .I2 (g11026));
AN2X1 gate14554(.O (g30152), .I1 (g28609), .I2 (g23767));
AN2X1 gate14555(.O (g24581), .I1 (g5124), .I2 (g23590));
AN2X1 gate14556(.O (g24714), .I1 (g6173), .I2 (g23699));
AN2X1 gate14557(.O (g32098), .I1 (g4732), .I2 (g30614));
AN2X1 gate14558(.O (g24450), .I1 (g3129), .I2 (g23067));
AN2X1 gate14559(.O (g21730), .I1 (g3025), .I2 (g20330));
AN2X1 gate14560(.O (g24315), .I1 (g4521), .I2 (g22228));
AN2X1 gate14561(.O (g21793), .I1 (g3412), .I2 (g20391));
AN2X1 gate14562(.O (g32272), .I1 (g31639), .I2 (g30310));
AN2X1 gate14563(.O (g22525), .I1 (g13006), .I2 (g19411));
AN2X1 gate14564(.O (g28159), .I1 (g8553), .I2 (g27317));
AN4X1 gate14565(.O (I31262), .I1 (g32833), .I2 (g32834), .I3 (g32835), .I4 (g32836));
AN2X1 gate14566(.O (g10878), .I1 (g7858), .I2 (g1135));
AN2X1 gate14567(.O (g18196), .I1 (g703), .I2 (g17821));
AN2X1 gate14568(.O (g22016), .I1 (g5747), .I2 (g21562));
AN2X1 gate14569(.O (g28125), .I1 (g27381), .I2 (g26209));
AN2X1 gate14570(.O (g15795), .I1 (g3566), .I2 (g14130));
AN2X1 gate14571(.O (g18695), .I1 (g4737), .I2 (g16053));
AN2X1 gate14572(.O (g28532), .I1 (g27394), .I2 (g20265));
AN2X1 gate14573(.O (g34396), .I1 (g34194), .I2 (g21337));
AN3X1 gate14574(.O (I18568), .I1 (g13156), .I2 (g11450), .I3 (g11498));
AN2X1 gate14575(.O (g24707), .I1 (g13295), .I2 (g22997));
AN2X1 gate14576(.O (g30731), .I1 (g11374), .I2 (g29361));
AN2X1 gate14577(.O (g29576), .I1 (g2177), .I2 (g28903));
AN2X1 gate14578(.O (g29585), .I1 (g1756), .I2 (g28920));
AN2X1 gate14579(.O (g21765), .I1 (g3231), .I2 (g20785));
AN3X1 gate14580(.O (g28158), .I1 (g26424), .I2 (g22763), .I3 (g27037));
AN4X1 gate14581(.O (I27523), .I1 (g20857), .I2 (g24111), .I3 (g24112), .I4 (g24113));
AN2X1 gate14582(.O (g18526), .I1 (g2555), .I2 (g15509));
AN2X1 gate14583(.O (g27269), .I1 (g25943), .I2 (g19734));
AN2X1 gate14584(.O (g29554), .I1 (g28997), .I2 (g22472));
AN2X1 gate14585(.O (g23690), .I1 (g14726), .I2 (g20978));
AN2X1 gate14586(.O (g19372), .I1 (g686), .I2 (g16289));
AN2X1 gate14587(.O (g26020), .I1 (g9559), .I2 (g25034));
AN2X1 gate14588(.O (g33241), .I1 (g32173), .I2 (g23128));
AN2X1 gate14589(.O (g34413), .I1 (g34094), .I2 (g22670));
AN2X1 gate14590(.O (g17424), .I1 (g1426), .I2 (g13176));
AN2X1 gate14591(.O (g11044), .I1 (g5343), .I2 (g10124));
AN4X1 gate14592(.O (I31191), .I1 (g30735), .I2 (g31829), .I3 (g32731), .I4 (g32732));
AN2X1 gate14593(.O (g27341), .I1 (g10203), .I2 (g26788));
AN2X1 gate14594(.O (g10967), .I1 (g7880), .I2 (g1448));
AN2X1 gate14595(.O (g29609), .I1 (g28482), .I2 (g11861));
AN2X1 gate14596(.O (g27268), .I1 (g25942), .I2 (g19733));
AN2X1 gate14597(.O (g32032), .I1 (g31373), .I2 (g16515));
AN2X1 gate14598(.O (g25780), .I1 (g25532), .I2 (g25527));
AN2X1 gate14599(.O (g15507), .I1 (g10970), .I2 (g13305));
AN2X1 gate14600(.O (g32140), .I1 (g31609), .I2 (g29961));
AN2X1 gate14601(.O (g28144), .I1 (g4608), .I2 (g27020));
AN2X1 gate14602(.O (g18402), .I1 (g2047), .I2 (g15373));
AN2X1 gate14603(.O (g18457), .I1 (g2319), .I2 (g15224));
AN2X1 gate14604(.O (g24590), .I1 (g6154), .I2 (g23413));
AN2X1 gate14605(.O (g29608), .I1 (g28568), .I2 (g11385));
AN2X1 gate14606(.O (g27180), .I1 (g26026), .I2 (g16654));
AN2X1 gate14607(.O (g19516), .I1 (g7824), .I2 (g16097));
AN2X1 gate14608(.O (g20094), .I1 (g8872), .I2 (g16631));
AN2X1 gate14609(.O (g27335), .I1 (g12087), .I2 (g26776));
AN3X1 gate14610(.O (g33683), .I1 (g33149), .I2 (g10727), .I3 (g22332));
AN2X1 gate14611(.O (g13738), .I1 (g8880), .I2 (g10572));
AN2X1 gate14612(.O (g25152), .I1 (g23383), .I2 (g20626));
AN2X1 gate14613(.O (g22042), .I1 (g5961), .I2 (g19147));
AN2X1 gate14614(.O (g26302), .I1 (g2393), .I2 (g25349));
AN2X1 gate14615(.O (g26357), .I1 (g22547), .I2 (g25525));
AN2X1 gate14616(.O (g29799), .I1 (g28271), .I2 (g10233));
AN2X1 gate14617(.O (g30583), .I1 (g19666), .I2 (g29355));
AN2X1 gate14618(.O (g16760), .I1 (g5559), .I2 (g14764));
AN2X1 gate14619(.O (g27667), .I1 (g26361), .I2 (g20601));
AN4X1 gate14620(.O (I31247), .I1 (g32812), .I2 (g32813), .I3 (g32814), .I4 (g32815));
AN2X1 gate14621(.O (g18706), .I1 (g4785), .I2 (g16782));
AN2X1 gate14622(.O (g18597), .I1 (g2975), .I2 (g16349));
AN2X1 gate14623(.O (g27965), .I1 (g25834), .I2 (g13117));
AN2X1 gate14624(.O (g13290), .I1 (g3897), .I2 (g11534));
AN2X1 gate14625(.O (g29798), .I1 (g28348), .I2 (g23260));
AN2X1 gate14626(.O (g22124), .I1 (g6613), .I2 (g19277));
AN2X1 gate14627(.O (g27131), .I1 (g26055), .I2 (g16588));
AN2X1 gate14628(.O (g30046), .I1 (g29108), .I2 (g10564));
AN2X1 gate14629(.O (g18256), .I1 (g1242), .I2 (g16897));
AN2X1 gate14630(.O (g29973), .I1 (g28981), .I2 (g9206));
AN2X1 gate14631(.O (g18689), .I1 (g15129), .I2 (g16752));
AN2X1 gate14632(.O (g31991), .I1 (g4912), .I2 (g30673));
AN3X1 gate14633(.O (g33515), .I1 (g32853), .I2 (I31271), .I3 (I31272));
AN2X1 gate14634(.O (g33882), .I1 (g33293), .I2 (g20587));
AN2X1 gate14635(.O (g18280), .I1 (g1367), .I2 (g16136));
AN2X1 gate14636(.O (g29805), .I1 (g28357), .I2 (g23270));
AN2X1 gate14637(.O (g33414), .I1 (g32367), .I2 (g21421));
AN2X1 gate14638(.O (g22686), .I1 (g19335), .I2 (g19577));
AN2X1 gate14639(.O (g22939), .I1 (g9708), .I2 (g21062));
AN2X1 gate14640(.O (g18688), .I1 (g4704), .I2 (g16752));
AN2X1 gate14641(.O (g18624), .I1 (g3490), .I2 (g17062));
AN2X1 gate14642(.O (g32162), .I1 (g31002), .I2 (g23014));
AN2X1 gate14643(.O (g18300), .I1 (g1306), .I2 (g16489));
AN2X1 gate14644(.O (g24196), .I1 (g333), .I2 (g22722));
AN2X1 gate14645(.O (g33407), .I1 (g32357), .I2 (g21406));
AN2X1 gate14646(.O (g34113), .I1 (g33734), .I2 (g19744));
AN2X1 gate14647(.O (g27502), .I1 (g26488), .I2 (g17677));
AN4X1 gate14648(.O (I31251), .I1 (g31710), .I2 (g31840), .I3 (g32817), .I4 (g32818));
AN2X1 gate14649(.O (g11427), .I1 (g5706), .I2 (g7158));
AN2X1 gate14650(.O (g22030), .I1 (g5909), .I2 (g19147));
AN4X1 gate14651(.O (I31272), .I1 (g32849), .I2 (g32850), .I3 (g32851), .I4 (g32852));
AN2X1 gate14652(.O (g22938), .I1 (g19782), .I2 (g19739));
AN2X1 gate14653(.O (g27557), .I1 (g26549), .I2 (g17774));
AN2X1 gate14654(.O (g22093), .I1 (g6423), .I2 (g18833));
AN2X1 gate14655(.O (g23533), .I1 (g19436), .I2 (g13015));
AN2X1 gate14656(.O (g11366), .I1 (g5016), .I2 (g10338));
AN3X1 gate14657(.O (g27210), .I1 (g26218), .I2 (g8373), .I3 (g2476));
AN2X1 gate14658(.O (g21298), .I1 (g7697), .I2 (g15825));
AN2X1 gate14659(.O (g29732), .I1 (g2514), .I2 (g29131));
AN2X1 gate14660(.O (g28289), .I1 (g27734), .I2 (g26575));
AN2X1 gate14661(.O (g21775), .I1 (g3372), .I2 (g20391));
AN3X1 gate14662(.O (I16671), .I1 (g10185), .I2 (g12461), .I3 (g12415));
AN2X1 gate14663(.O (g13632), .I1 (g10232), .I2 (g12228));
AN2X1 gate14664(.O (g18157), .I1 (g15057), .I2 (g17433));
AN2X1 gate14665(.O (g23775), .I1 (g14872), .I2 (g21267));
AN2X1 gate14666(.O (g22065), .I1 (g6203), .I2 (g19210));
AN3X1 gate14667(.O (g34105), .I1 (g33778), .I2 (g9104), .I3 (g18957));
AN3X1 gate14668(.O (g28224), .I1 (g27163), .I2 (g22763), .I3 (g27064));
AN2X1 gate14669(.O (g34743), .I1 (g8951), .I2 (g34703));
AN3X1 gate14670(.O (I17585), .I1 (g14988), .I2 (g11450), .I3 (g11498));
AN2X1 gate14671(.O (g28571), .I1 (g27458), .I2 (g20435));
AN2X1 gate14672(.O (g24402), .I1 (g4749), .I2 (g22857));
AN2X1 gate14673(.O (g29761), .I1 (g28310), .I2 (g23228));
AN4X1 gate14674(.O (I31032), .I1 (g32501), .I2 (g32502), .I3 (g32503), .I4 (g32504));
AN2X1 gate14675(.O (g18231), .I1 (g1105), .I2 (g16326));
AN2X1 gate14676(.O (g21737), .I1 (g3068), .I2 (g20330));
AN2X1 gate14677(.O (g32246), .I1 (g31246), .I2 (g20326));
AN4X1 gate14678(.O (g27469), .I1 (g8046), .I2 (g26314), .I3 (g518), .I4 (g9077));
AN2X1 gate14679(.O (g22219), .I1 (g19953), .I2 (g20887));
AN2X1 gate14680(.O (g25928), .I1 (g25022), .I2 (g23436));
AN2X1 gate14681(.O (g8583), .I1 (g2917), .I2 (g2912));
AN2X1 gate14682(.O (g27286), .I1 (g6856), .I2 (g26634));
AN2X1 gate14683(.O (g33441), .I1 (g32251), .I2 (g29722));
AN2X1 gate14684(.O (g31206), .I1 (g30260), .I2 (g23890));
AN2X1 gate14685(.O (g10656), .I1 (g3782), .I2 (g7952));
AN4X1 gate14686(.O (g27039), .I1 (g7738), .I2 (g5527), .I3 (g5535), .I4 (g26223));
AN2X1 gate14687(.O (g22218), .I1 (g19951), .I2 (g20875));
AN2X1 gate14688(.O (g28495), .I1 (g27012), .I2 (g12465));
AN2X1 gate14689(.O (g32071), .I1 (g27236), .I2 (g31070));
AN4X1 gate14690(.O (I31061), .I1 (g30825), .I2 (g31806), .I3 (g32543), .I4 (g32544));
AN2X1 gate14691(.O (g21856), .I1 (g3929), .I2 (g21070));
AN3X1 gate14692(.O (g10823), .I1 (g7704), .I2 (g5180), .I3 (g5188));
AN2X1 gate14693(.O (g14295), .I1 (g1811), .I2 (g11894));
AN2X1 gate14694(.O (g21995), .I1 (g5611), .I2 (g19074));
AN2X1 gate14695(.O (g31759), .I1 (g21291), .I2 (g29385));
AN2X1 gate14696(.O (g23856), .I1 (g4116), .I2 (g19483));
AN2X1 gate14697(.O (g14680), .I1 (g12024), .I2 (g12053));
AN2X1 gate14698(.O (g33759), .I1 (g33123), .I2 (g22847));
AN3X1 gate14699(.O (g33725), .I1 (g22626), .I2 (g10851), .I3 (g33176));
AN2X1 gate14700(.O (g24001), .I1 (g19651), .I2 (g10951));
AN2X1 gate14701(.O (g21880), .I1 (g4135), .I2 (g19801));
AN2X1 gate14702(.O (g29329), .I1 (g7995), .I2 (g28353));
AN2X1 gate14703(.O (g25113), .I1 (g23346), .I2 (g20577));
AN2X1 gate14704(.O (g18511), .I1 (g2599), .I2 (g15509));
AN3X1 gate14705(.O (g29207), .I1 (g24131), .I2 (I27533), .I3 (I27534));
AN2X1 gate14706(.O (g25787), .I1 (g24792), .I2 (g20887));
AN2X1 gate14707(.O (g32147), .I1 (g31616), .I2 (g29980));
AN2X1 gate14708(.O (g18763), .I1 (g5481), .I2 (g17929));
AN2X1 gate14709(.O (g31758), .I1 (g30115), .I2 (g23945));
AN2X1 gate14710(.O (g33114), .I1 (g22139), .I2 (g31945));
AN2X1 gate14711(.O (g24706), .I1 (g15910), .I2 (g22996));
AN2X1 gate14712(.O (g26249), .I1 (g1858), .I2 (g25300));
AN2X1 gate14713(.O (g33758), .I1 (g33133), .I2 (g20269));
AN2X1 gate14714(.O (g22160), .I1 (g8005), .I2 (g19795));
AN2X1 gate14715(.O (g27601), .I1 (g26766), .I2 (g26737));
AN2X1 gate14716(.O (g33082), .I1 (g32389), .I2 (g18877));
AN2X1 gate14717(.O (g21512), .I1 (g16225), .I2 (g10881));
AN3X1 gate14718(.O (g29328), .I1 (g28553), .I2 (g6928), .I3 (g3990));
AN2X1 gate14719(.O (g27677), .I1 (g13021), .I2 (g25888));
AN2X1 gate14720(.O (g25357), .I1 (g23810), .I2 (g23786));
AN2X1 gate14721(.O (g29538), .I1 (g2563), .I2 (g28914));
AN2X1 gate14722(.O (g11127), .I1 (g6479), .I2 (g10022));
AN2X1 gate14723(.O (g24923), .I1 (g23129), .I2 (g20167));
AN2X1 gate14724(.O (g25105), .I1 (g13973), .I2 (g23505));
AN2X1 gate14725(.O (g10966), .I1 (g9226), .I2 (g7948));
AN2X1 gate14726(.O (g31744), .I1 (g30092), .I2 (g23902));
AN2X1 gate14727(.O (g24688), .I1 (g22681), .I2 (g22663));
AN2X1 gate14728(.O (g26204), .I1 (g1720), .I2 (g25275));
AN2X1 gate14729(.O (g24624), .I1 (g16524), .I2 (g22867));
AN2X1 gate14730(.O (g24300), .I1 (g15123), .I2 (g22228));
AN3X1 gate14731(.O (I24579), .I1 (g5731), .I2 (g5736), .I3 (g9875));
AN2X1 gate14732(.O (g26779), .I1 (g24497), .I2 (g23620));
AN2X1 gate14733(.O (g33345), .I1 (g32229), .I2 (g20671));
AN2X1 gate14734(.O (g32151), .I1 (g31639), .I2 (g29996));
AN2X1 gate14735(.O (g32172), .I1 (g2767), .I2 (g31608));
AN4X1 gate14736(.O (I31162), .I1 (g32689), .I2 (g32690), .I3 (g32691), .I4 (g32692));
AN2X1 gate14737(.O (g31940), .I1 (g943), .I2 (g30735));
AN2X1 gate14738(.O (g18456), .I1 (g2338), .I2 (g15224));
AN2X1 gate14739(.O (g33849), .I1 (g33262), .I2 (g20387));
AN2X1 gate14740(.O (g30027), .I1 (g29104), .I2 (g12550));
AN2X1 gate14741(.O (g33399), .I1 (g32346), .I2 (g21379));
AN2X1 gate14742(.O (g21831), .I1 (g3782), .I2 (g20453));
AN2X1 gate14743(.O (g26778), .I1 (g25501), .I2 (g20923));
AN2X1 gate14744(.O (g34662), .I1 (g34576), .I2 (g18931));
AN2X1 gate14745(.O (g16845), .I1 (g6593), .I2 (g15011));
AN2X1 gate14746(.O (g11956), .I1 (g2070), .I2 (g7411));
AN2X1 gate14747(.O (g18480), .I1 (g2437), .I2 (g15426));
OR2X1 gate14748(.O (g32367), .I1 (g29880), .I2 (g31309));
OR2X1 gate14749(.O (g34890), .I1 (g34863), .I2 (g21674));
OR2X1 gate14750(.O (g28668), .I1 (g27411), .I2 (g16617));
OR2X1 gate14751(.O (g34249), .I1 (g34110), .I2 (g21702));
OR2X1 gate14752(.O (g13095), .I1 (g11374), .I2 (g1287));
OR2X1 gate14753(.O (g30482), .I1 (g30230), .I2 (g21978));
OR2X1 gate14754(.O (g24231), .I1 (g22589), .I2 (g18201));
OR2X1 gate14755(.O (g13888), .I1 (g2941), .I2 (g11691));
OR2X1 gate14756(.O (g26945), .I1 (g26379), .I2 (g24283));
OR2X1 gate14757(.O (g30552), .I1 (g30283), .I2 (g22123));
OR2X1 gate14758(.O (g34003), .I1 (g33866), .I2 (g18452));
OR2X1 gate14759(.O (g23989), .I1 (g20581), .I2 (g17179));
OR2X1 gate14760(.O (g29235), .I1 (g28110), .I2 (g18260));
OR2X1 gate14761(.O (g28525), .I1 (g27284), .I2 (g26176));
OR2X1 gate14762(.O (g34204), .I1 (g33832), .I2 (g33833));
OR4X1 gate14763(.O (I28566), .I1 (g29201), .I2 (g29202), .I3 (g29203), .I4 (g28035));
OR2X1 gate14764(.O (g14309), .I1 (g10320), .I2 (g11048));
OR4X1 gate14765(.O (I30330), .I1 (g29385), .I2 (g31376), .I3 (g30735), .I4 (g30825));
OR2X1 gate14766(.O (g24854), .I1 (g21453), .I2 (g24002));
OR2X1 gate14767(.O (g30081), .I1 (g28454), .I2 (g11366));
OR2X1 gate14768(.O (g32227), .I1 (g31146), .I2 (g29648));
OR2X1 gate14769(.O (g33962), .I1 (g33822), .I2 (g18123));
OR2X1 gate14770(.O (g19575), .I1 (g15693), .I2 (g13042));
OR2X1 gate14771(.O (g27556), .I1 (g26097), .I2 (g24687));
OR2X1 gate14772(.O (g25662), .I1 (g24656), .I2 (g21787));
OR2X1 gate14773(.O (g28544), .I1 (g27300), .I2 (g26229));
OR2X1 gate14774(.O (g30356), .I1 (g30096), .I2 (g18365));
OR2X1 gate14775(.O (g27580), .I1 (g26159), .I2 (g24749));
OR2X1 gate14776(.O (g34647), .I1 (g34558), .I2 (g18820));
OR2X1 gate14777(.O (g26932), .I1 (g26684), .I2 (g18549));
OR4X1 gate14778(.O (I31859), .I1 (g33501), .I2 (g33502), .I3 (g33503), .I4 (g33504));
OR2X1 gate14779(.O (g33049), .I1 (g31966), .I2 (g21929));
OR2X1 gate14780(.O (g30380), .I1 (g30161), .I2 (g18492));
OR2X1 gate14781(.O (g34826), .I1 (g34742), .I2 (g34685));
OR3X1 gate14782(.O (g16926), .I1 (g14061), .I2 (g11804), .I3 (g11780));
OR3X1 gate14783(.O (I25736), .I1 (g12), .I2 (g22150), .I3 (g20277));
OR4X1 gate14784(.O (I31858), .I1 (g33497), .I2 (g33498), .I3 (g33499), .I4 (g33500));
OR2X1 gate14785(.O (g33048), .I1 (g31960), .I2 (g21928));
OR2X1 gate14786(.O (g7684), .I1 (g4072), .I2 (g4176));
OR2X1 gate14787(.O (g25710), .I1 (g25031), .I2 (g21961));
OR2X1 gate14788(.O (g28610), .I1 (g27347), .I2 (g16484));
OR2X1 gate14789(.O (g26897), .I1 (g26611), .I2 (g18176));
OR2X1 gate14790(.O (g34090), .I1 (g33676), .I2 (g33680));
OR2X1 gate14791(.O (g26961), .I1 (g26280), .I2 (g24306));
OR2X1 gate14792(.O (g28705), .I1 (g27460), .I2 (g16672));
OR2X1 gate14793(.O (g28042), .I1 (g24148), .I2 (g26879));
OR2X1 gate14794(.O (g30672), .I1 (g13737), .I2 (g29752));
OR2X1 gate14795(.O (g34233), .I1 (g32455), .I2 (g33951));
OR2X1 gate14796(.O (g13211), .I1 (g11294), .I2 (g7567));
OR2X1 gate14797(.O (g33004), .I1 (g32246), .I2 (g18431));
OR2X1 gate14798(.O (g31221), .I1 (g29494), .I2 (g28204));
OR3X1 gate14799(.O (g23198), .I1 (g20214), .I2 (g20199), .I3 (I22298));
OR4X1 gate14800(.O (I31844), .I1 (g33474), .I2 (g33475), .I3 (g33476), .I4 (g33477));
OR2X1 gate14801(.O (g27179), .I1 (g25816), .I2 (g24409));
OR2X1 gate14802(.O (g28188), .I1 (g22535), .I2 (g27108));
OR2X1 gate14803(.O (g33613), .I1 (g33248), .I2 (g18649));
OR2X1 gate14804(.O (g34331), .I1 (g27121), .I2 (g34072));
OR2X1 gate14805(.O (g30513), .I1 (g30200), .I2 (g22034));
OR2X1 gate14806(.O (g30449), .I1 (g29845), .I2 (g21858));
OR2X1 gate14807(.O (g33947), .I1 (g32438), .I2 (g33457));
OR2X1 gate14808(.O (g34449), .I1 (g34279), .I2 (g18662));
OR2X1 gate14809(.O (g25647), .I1 (g24725), .I2 (g21740));
OR2X1 gate14810(.O (g24243), .I1 (g22992), .I2 (g18254));
OR2X1 gate14811(.O (g33273), .I1 (g32122), .I2 (g29553));
OR2X1 gate14812(.O (g28030), .I1 (g24018), .I2 (g26874));
OR2X1 gate14813(.O (g33605), .I1 (g33352), .I2 (g18521));
OR2X1 gate14814(.O (g25945), .I1 (g24427), .I2 (g22307));
OR2X1 gate14815(.O (g28093), .I1 (g27981), .I2 (g21951));
OR2X1 gate14816(.O (g30448), .I1 (g29809), .I2 (g21857));
OR2X1 gate14817(.O (g34897), .I1 (g34861), .I2 (g21682));
OR2X1 gate14818(.O (g34448), .I1 (g34365), .I2 (g18553));
OR2X1 gate14819(.O (g30505), .I1 (g30168), .I2 (g22026));
OR2X1 gate14820(.O (g29114), .I1 (g27646), .I2 (g26602));
OR2X1 gate14821(.O (g30404), .I1 (g29758), .I2 (g21763));
OR2X1 gate14822(.O (g28065), .I1 (g27299), .I2 (g21792));
OR2X1 gate14823(.O (g27800), .I1 (g17321), .I2 (g26703));
OR2X1 gate14824(.O (g24269), .I1 (g23131), .I2 (g18613));
OR2X1 gate14825(.O (g34404), .I1 (g34182), .I2 (g25102));
OR3X1 gate14826(.O (g33951), .I1 (g33469), .I2 (I31838), .I3 (I31839));
OR2X1 gate14827(.O (g33972), .I1 (g33941), .I2 (g18335));
OR2X1 gate14828(.O (g24341), .I1 (g23564), .I2 (g18771));
OR2X1 gate14829(.O (g33033), .I1 (g32333), .I2 (g21843));
OR2X1 gate14830(.O (g24268), .I1 (g23025), .I2 (g18612));
OR2X1 gate14831(.O (g25651), .I1 (g24680), .I2 (g21744));
OR2X1 gate14832(.O (g25672), .I1 (g24647), .I2 (g21829));
OR2X1 gate14833(.O (g33234), .I1 (g32039), .I2 (g32043));
OR2X1 gate14834(.O (g34026), .I1 (g33715), .I2 (g18682));
OR2X1 gate14835(.O (g32427), .I1 (g8928), .I2 (g30583));
OR2X1 gate14836(.O (g13296), .I1 (g10626), .I2 (g10657));
OR2X1 gate14837(.O (g23087), .I1 (g19487), .I2 (g15852));
OR2X1 gate14838(.O (g29849), .I1 (g26049), .I2 (g28273));
OR2X1 gate14839(.O (g13969), .I1 (g11448), .I2 (g8913));
OR2X1 gate14840(.O (g26343), .I1 (g1514), .I2 (g24609));
OR2X1 gate14841(.O (g19522), .I1 (g17057), .I2 (g14180));
OR2X1 gate14842(.O (g29848), .I1 (g28260), .I2 (g26077));
OR2X1 gate14843(.O (g24335), .I1 (g22165), .I2 (g18678));
OR2X1 gate14844(.O (g26971), .I1 (g26325), .I2 (g24333));
OR2X1 gate14845(.O (g34723), .I1 (g34710), .I2 (g18139));
OR2X1 gate14846(.O (g30433), .I1 (g29899), .I2 (g21817));
OR2X1 gate14847(.O (g34149), .I1 (g33760), .I2 (g19674));
OR2X1 gate14848(.O (g30387), .I1 (g30151), .I2 (g18524));
OR2X1 gate14849(.O (g24965), .I1 (g22667), .I2 (g23825));
OR2X1 gate14850(.O (g32226), .I1 (g31145), .I2 (g29645));
OR2X1 gate14851(.O (g29263), .I1 (g28239), .I2 (g18617));
OR2X1 gate14852(.O (g34620), .I1 (g34529), .I2 (g18582));
OR2X1 gate14853(.O (g34148), .I1 (g33758), .I2 (g19656));
OR2X1 gate14854(.O (g25717), .I1 (g25106), .I2 (g21968));
OR2X1 gate14855(.O (g27543), .I1 (g26085), .I2 (g24670));
OR2X1 gate14856(.O (g30104), .I1 (g28478), .I2 (g11427));
OR2X1 gate14857(.O (g33012), .I1 (g32274), .I2 (g18483));
OR2X1 gate14858(.O (g19949), .I1 (g17671), .I2 (g14681));
OR2X1 gate14859(.O (g30343), .I1 (g29344), .I2 (g18278));
OR2X1 gate14860(.O (g34646), .I1 (g34557), .I2 (g18803));
OR2X1 gate14861(.O (g24557), .I1 (g22308), .I2 (g19207));
OR2X1 gate14862(.O (g24210), .I1 (g22900), .I2 (g18125));
OR2X1 gate14863(.O (g27569), .I1 (g26124), .I2 (g24721));
OR2X1 gate14864(.O (g34971), .I1 (g34869), .I2 (g34962));
OR2X1 gate14865(.O (g33541), .I1 (g33101), .I2 (g18223));
OR2X1 gate14866(.O (g31473), .I1 (g26180), .I2 (g29666));
OR2X1 gate14867(.O (g28075), .I1 (g27083), .I2 (g21877));
OR2X1 gate14868(.O (g30369), .I1 (g30066), .I2 (g18439));
OR2X1 gate14869(.O (g24443), .I1 (g23917), .I2 (g21378));
OR2X1 gate14870(.O (g19904), .I1 (g17636), .I2 (g14654));
OR2X1 gate14871(.O (g23171), .I1 (g19536), .I2 (g15903));
OR2X1 gate14872(.O (g24279), .I1 (g23218), .I2 (g15105));
OR2X1 gate14873(.O (g26896), .I1 (g26341), .I2 (g18171));
OR2X1 gate14874(.O (g34369), .I1 (g26279), .I2 (g34136));
OR2X1 gate14875(.O (g28595), .I1 (g27335), .I2 (g26290));
OR2X1 gate14876(.O (g14030), .I1 (g11037), .I2 (g11046));
OR2X1 gate14877(.O (g30368), .I1 (g30098), .I2 (g18435));
OR2X1 gate14878(.O (g24278), .I1 (g23201), .I2 (g18648));
OR2X1 gate14879(.O (g25723), .I1 (g25033), .I2 (g22006));
OR2X1 gate14880(.O (g28623), .I1 (g27361), .I2 (g16520));
OR2X1 gate14881(.O (g34368), .I1 (g26274), .I2 (g34135));
OR2X1 gate14882(.O (g33788), .I1 (g33122), .I2 (g32041));
OR2X1 gate14883(.O (g31325), .I1 (g29625), .I2 (g29639));
OR2X1 gate14884(.O (g32385), .I1 (g31480), .I2 (g29938));
OR2X1 gate14885(.O (g31920), .I1 (g31493), .I2 (g22045));
OR2X1 gate14886(.O (g32980), .I1 (g32254), .I2 (g18198));
OR2X1 gate14887(.O (g30412), .I1 (g29885), .I2 (g21771));
OR2X1 gate14888(.O (g33535), .I1 (g33233), .I2 (g21711));
OR2X1 gate14889(.O (g24468), .I1 (g10925), .I2 (g22400));
OR2X1 gate14890(.O (g32354), .I1 (g29854), .I2 (g31285));
OR2X1 gate14891(.O (g34850), .I1 (g34841), .I2 (g18185));
OR2X1 gate14892(.O (g34412), .I1 (g34187), .I2 (g25143));
OR2X1 gate14893(.O (g28419), .I1 (g27221), .I2 (g15884));
OR2X1 gate14894(.O (g27974), .I1 (g26544), .I2 (g25063));
OR2X1 gate14895(.O (g33946), .I1 (g32434), .I2 (g33456));
OR2X1 gate14896(.O (g25646), .I1 (g24706), .I2 (g21739));
OR2X1 gate14897(.O (g28418), .I1 (g27220), .I2 (g15882));
OR2X1 gate14898(.O (g20187), .I1 (g16202), .I2 (g13491));
OR2X1 gate14899(.O (g26959), .I1 (g26381), .I2 (g24299));
OR2X1 gate14900(.O (g26925), .I1 (g25939), .I2 (g18301));
OR2X1 gate14901(.O (g34011), .I1 (g33884), .I2 (g18479));
OR2X1 gate14902(.O (g26958), .I1 (g26395), .I2 (g24297));
OR2X1 gate14903(.O (g29273), .I1 (g28269), .I2 (g18639));
OR2X1 gate14904(.O (g31291), .I1 (g29581), .I2 (g29593));
OR4X1 gate14905(.O (g17570), .I1 (g14419), .I2 (g14397), .I3 (g11999), .I4 (I18495));
OR2X1 gate14906(.O (g33291), .I1 (g32154), .I2 (g13477));
OR2X1 gate14907(.O (g26386), .I1 (g24719), .I2 (g23023));
OR3X1 gate14908(.O (g32426), .I1 (g26105), .I2 (g26131), .I3 (g30613));
OR2X1 gate14909(.O (g28194), .I1 (g22540), .I2 (g27122));
OR2X1 gate14910(.O (g28589), .I1 (g27331), .I2 (g26285));
OR2X1 gate14911(.O (g26944), .I1 (g26130), .I2 (g18658));
OR2X1 gate14912(.O (g20169), .I1 (g16184), .I2 (g13460));
OR2X1 gate14913(.O (g27579), .I1 (g26157), .I2 (g24748));
OR2X1 gate14914(.O (g29234), .I1 (g28415), .I2 (g18239));
OR2X1 gate14915(.O (g30379), .I1 (g30089), .I2 (g18491));
OR2X1 gate14916(.O (g34627), .I1 (g34534), .I2 (g18644));
OR2X1 gate14917(.O (g27578), .I1 (g26155), .I2 (g24747));
OR4X1 gate14918(.O (g17594), .I1 (g14450), .I2 (g14420), .I3 (g12025), .I4 (I18543));
OR2X1 gate14919(.O (g28401), .I1 (g27212), .I2 (g15871));
OR2X1 gate14920(.O (g31760), .I1 (g30007), .I2 (g30027));
OR2X1 gate14921(.O (g34379), .I1 (g26312), .I2 (g34143));
OR2X1 gate14922(.O (g33029), .I1 (g32332), .I2 (g21798));
OR2X1 gate14923(.O (g32211), .I1 (g31124), .I2 (g29603));
OR2X1 gate14924(.O (g30378), .I1 (g30125), .I2 (g18487));
OR2X1 gate14925(.O (g21901), .I1 (g21251), .I2 (g15115));
OR2X1 gate14926(.O (g20217), .I1 (g16221), .I2 (g13523));
OR2X1 gate14927(.O (g33028), .I1 (g32325), .I2 (g21797));
OR2X1 gate14928(.O (g30386), .I1 (g30139), .I2 (g18523));
OR2X1 gate14929(.O (g24363), .I1 (g7831), .I2 (g22138));
OR2X1 gate14930(.O (g26793), .I1 (g24478), .I2 (g7520));
OR2X1 gate14931(.O (g28118), .I1 (g27821), .I2 (g26815));
OR3X1 gate14932(.O (g13526), .I1 (g209), .I2 (g10685), .I3 (g301));
OR2X1 gate14933(.O (g24478), .I1 (g11003), .I2 (g22450));
OR2X1 gate14934(.O (g34603), .I1 (g34561), .I2 (g15075));
OR2X1 gate14935(.O (g25716), .I1 (g25088), .I2 (g21967));
OR2X1 gate14936(.O (g28749), .I1 (g27523), .I2 (g16764));
OR2X1 gate14937(.O (g26690), .I1 (g10776), .I2 (g24433));
OR2X1 gate14938(.O (g25582), .I1 (g21662), .I2 (g24152));
OR2X1 gate14939(.O (g28748), .I1 (g27522), .I2 (g16763));
OR2X1 gate14940(.O (g28704), .I1 (g27459), .I2 (g16671));
OR2X1 gate14941(.O (g24580), .I1 (g22340), .I2 (g13096));
OR2X1 gate14942(.O (g31927), .I1 (g31500), .I2 (g22091));
OR2X1 gate14943(.O (g30429), .I1 (g29844), .I2 (g21813));
OR2X1 gate14944(.O (g28305), .I1 (g27103), .I2 (g15793));
OR2X1 gate14945(.O (g28053), .I1 (g27393), .I2 (g18168));
OR2X1 gate14946(.O (g32987), .I1 (g32311), .I2 (g18323));
OR2X1 gate14947(.O (g32250), .I1 (g30598), .I2 (g29351));
OR2X1 gate14948(.O (g34802), .I1 (g34757), .I2 (g18589));
OR2X1 gate14949(.O (g25627), .I1 (g24503), .I2 (g18247));
OR2X1 gate14950(.O (g30428), .I1 (g29807), .I2 (g21812));
OR2X1 gate14951(.O (g34730), .I1 (g34658), .I2 (g18271));
OR2X1 gate14952(.O (g34793), .I1 (g34744), .I2 (g18570));
OR4X1 gate14953(.O (I26643), .I1 (g27073), .I2 (g27058), .I3 (g27045), .I4 (g27040));
OR2X1 gate14954(.O (g13077), .I1 (g11330), .I2 (g943));
OR3X1 gate14955(.O (I18492), .I1 (g14538), .I2 (g14513), .I3 (g14446));
OR2X1 gate14956(.O (g28101), .I1 (g27691), .I2 (g22062));
OR2X1 gate14957(.O (g33240), .I1 (g32052), .I2 (g32068));
OR2X1 gate14958(.O (g13597), .I1 (g9247), .I2 (g11149));
OR2X1 gate14959(.O (g28560), .I1 (g27311), .I2 (g26249));
OR2X1 gate14960(.O (g31903), .I1 (g31374), .I2 (g21911));
OR2X1 gate14961(.O (g30549), .I1 (g30215), .I2 (g22120));
OR2X1 gate14962(.O (g25603), .I1 (g24698), .I2 (g18114));
OR2X1 gate14963(.O (g25742), .I1 (g25093), .I2 (g22057));
OR2X1 gate14964(.O (g31755), .I1 (g29991), .I2 (g30008));
OR2X1 gate14965(.O (g33604), .I1 (g33345), .I2 (g18520));
OR2X1 gate14966(.O (g30548), .I1 (g30204), .I2 (g22119));
OR2X1 gate14967(.O (g10589), .I1 (g7223), .I2 (g7201));
OR2X1 gate14968(.O (g29325), .I1 (g28813), .I2 (g27820));
OR2X1 gate14969(.O (g13300), .I1 (g10656), .I2 (g10676));
OR2X1 gate14970(.O (g31770), .I1 (g30034), .I2 (g30047));
OR2X1 gate14971(.O (g30504), .I1 (g30253), .I2 (g22025));
OR2X1 gate14972(.O (g28064), .I1 (g27298), .I2 (g21781));
OR2X1 gate14973(.O (g33563), .I1 (g33361), .I2 (g18383));
OR2X1 gate14974(.O (g33981), .I1 (g33856), .I2 (g18371));
OR2X1 gate14975(.O (g25681), .I1 (g24710), .I2 (g18636));
OR2X1 gate14976(.O (g28733), .I1 (g27507), .I2 (g16735));
OR2X1 gate14977(.O (g26299), .I1 (g24551), .I2 (g22665));
OR3X1 gate14978(.O (g30317), .I1 (g29208), .I2 (I28566), .I3 (I28567));
OR2X1 gate14979(.O (g25730), .I1 (g25107), .I2 (g22013));
OR2X1 gate14980(.O (g22304), .I1 (g21347), .I2 (g17693));
OR2X1 gate14981(.O (g14119), .I1 (g10776), .I2 (g8703));
OR2X1 gate14982(.O (g31767), .I1 (g30031), .I2 (g30043));
OR2X1 gate14983(.O (g33794), .I1 (g33126), .I2 (g32053));
OR2X1 gate14984(.O (g34002), .I1 (g33857), .I2 (g18451));
OR2X1 gate14985(.O (g33262), .I1 (g32112), .I2 (g29528));
OR2X1 gate14986(.O (g31899), .I1 (g31470), .I2 (g21907));
OR2X1 gate14987(.O (g34057), .I1 (g33911), .I2 (g33915));
OR2X1 gate14988(.O (g28665), .I1 (g27409), .I2 (g16614));
OR2X1 gate14989(.O (g30128), .I1 (g28495), .I2 (g11497));
OR2X1 gate14990(.O (g33990), .I1 (g33882), .I2 (g18399));
OR2X1 gate14991(.O (g24334), .I1 (g23991), .I2 (g18676));
OR2X1 gate14992(.O (g25690), .I1 (g24864), .I2 (g21889));
OR2X1 gate14993(.O (g26737), .I1 (g24460), .I2 (g10720));
OR2X1 gate14994(.O (g29291), .I1 (g28660), .I2 (g18767));
OR2X1 gate14995(.O (g31898), .I1 (g31707), .I2 (g21906));
OR2X1 gate14996(.O (g34626), .I1 (g34533), .I2 (g18627));
OR2X1 gate14997(.O (g30533), .I1 (g30203), .I2 (g22079));
OR2X1 gate14998(.O (g22653), .I1 (g18993), .I2 (g15654));
OR2X1 gate14999(.O (g30298), .I1 (g28245), .I2 (g27251));
OR3X1 gate15000(.O (g23687), .I1 (g21384), .I2 (g21363), .I3 (I22830));
OR2X1 gate15001(.O (g26880), .I1 (g26610), .I2 (g24186));
OR2X1 gate15002(.O (g24216), .I1 (g23416), .I2 (g18197));
OR2X1 gate15003(.O (g23374), .I1 (g19767), .I2 (g13514));
OR2X1 gate15004(.O (g32202), .I1 (g31069), .I2 (g13410));
OR2X1 gate15005(.O (g22636), .I1 (g18943), .I2 (g15611));
OR2X1 gate15006(.O (g26512), .I1 (g24786), .I2 (g23130));
OR2X1 gate15007(.O (g32257), .I1 (g31184), .I2 (g29708));
OR2X1 gate15008(.O (g13660), .I1 (g8183), .I2 (g12527));
OR2X1 gate15009(.O (g32979), .I1 (g32181), .I2 (g18177));
OR2X1 gate15010(.O (g29506), .I1 (g28148), .I2 (g25880));
OR2X1 gate15011(.O (g34232), .I1 (g33451), .I2 (g33944));
OR2X1 gate15012(.O (g32978), .I1 (g32197), .I2 (g18145));
OR2X1 gate15013(.O (g28074), .I1 (g27119), .I2 (g21876));
OR2X1 gate15014(.O (g33573), .I1 (g33343), .I2 (g18415));
OR2X1 gate15015(.O (g31247), .I1 (g29513), .I2 (g13324));
OR2X1 gate15016(.O (g28594), .I1 (g27334), .I2 (g26289));
OR2X1 gate15017(.O (g31926), .I1 (g31765), .I2 (g22090));
OR2X1 gate15018(.O (g32986), .I1 (g31996), .I2 (g18280));
OR2X1 gate15019(.O (g27253), .I1 (g24661), .I2 (g26052));
OR2X1 gate15020(.O (g33389), .I1 (g32272), .I2 (g29964));
OR2X1 gate15021(.O (g33045), .I1 (g32206), .I2 (g24328));
OR2X1 gate15022(.O (g22664), .I1 (g19139), .I2 (g15694));
OR2X1 gate15023(.O (g34856), .I1 (g34811), .I2 (g34743));
OR2X1 gate15024(.O (g25626), .I1 (g24499), .I2 (g18235));
OR2X1 gate15025(.O (g33612), .I1 (g33247), .I2 (g18633));
OR2X1 gate15026(.O (g34261), .I1 (g34074), .I2 (g18688));
OR2X1 gate15027(.O (g34880), .I1 (g34867), .I2 (g18153));
OR2X1 gate15028(.O (g8921), .I1 (I12902), .I2 (I12903));
OR2X1 gate15029(.O (g30512), .I1 (g30191), .I2 (g22033));
OR2X1 gate15030(.O (g33534), .I1 (g33186), .I2 (g21700));
OR2X1 gate15031(.O (g27236), .I1 (g24620), .I2 (g25974));
OR2X1 gate15032(.O (g32094), .I1 (g30612), .I2 (g29363));
OR2X1 gate15033(.O (g31251), .I1 (g25973), .I2 (g29527));
OR2X1 gate15034(.O (g22585), .I1 (g20915), .I2 (g21061));
OR2X1 gate15035(.O (g33251), .I1 (g32096), .I2 (g29509));
OR2X1 gate15036(.O (g24242), .I1 (g22834), .I2 (g18253));
OR2X1 gate15037(.O (g33272), .I1 (g32121), .I2 (g29551));
OR2X1 gate15038(.O (g28092), .I1 (g27666), .I2 (g21924));
OR4X1 gate15039(.O (I30124), .I1 (g31070), .I2 (g31154), .I3 (g30614), .I4 (g30673));
OR2X1 gate15040(.O (g28518), .I1 (g27281), .I2 (g26158));
OR2X1 gate15041(.O (g21893), .I1 (g20094), .I2 (g18655));
OR2X1 gate15042(.O (g29240), .I1 (g28655), .I2 (g18328));
OR2X1 gate15043(.O (g26080), .I1 (g19393), .I2 (g24502));
OR3X1 gate15044(.O (I12583), .I1 (g1157), .I2 (g1239), .I3 (g990));
OR2X1 gate15045(.O (g25737), .I1 (g25045), .I2 (g22052));
OR2X1 gate15046(.O (g26924), .I1 (g26153), .I2 (g18291));
OR2X1 gate15047(.O (g30445), .I1 (g29772), .I2 (g21854));
OR2X1 gate15048(.O (g33032), .I1 (g32326), .I2 (g21842));
OR2X1 gate15049(.O (g34445), .I1 (g34382), .I2 (g18548));
OR2X1 gate15050(.O (g30499), .I1 (g30261), .I2 (g21995));
OR2X1 gate15051(.O (g33997), .I1 (g33871), .I2 (g18427));
OR2X1 gate15052(.O (g25697), .I1 (g25086), .I2 (g21916));
OR4X1 gate15053(.O (g25856), .I1 (g25518), .I2 (g25510), .I3 (g25488), .I4 (g25462));
OR2X1 gate15054(.O (g30498), .I1 (g30251), .I2 (g21994));
OR2X1 gate15055(.O (g25261), .I1 (g23348), .I2 (g20193));
OR2X1 gate15056(.O (g33061), .I1 (g32334), .I2 (g22050));
OR2X1 gate15057(.O (g24265), .I1 (g22316), .I2 (g18560));
OR2X1 gate15058(.O (g26342), .I1 (g8407), .I2 (g24591));
OR2X1 gate15059(.O (g31766), .I1 (g30029), .I2 (g30042));
OR2X1 gate15060(.O (g31871), .I1 (g30596), .I2 (g18279));
OR2X1 gate15061(.O (g30611), .I1 (g13671), .I2 (g29743));
OR2X1 gate15062(.O (g24841), .I1 (g21420), .I2 (g23998));
OR2X1 gate15063(.O (g34611), .I1 (g34508), .I2 (g18565));
OR2X1 gate15064(.O (g23255), .I1 (g19655), .I2 (g16122));
OR2X1 gate15065(.O (g34722), .I1 (g34707), .I2 (g18137));
OR2X1 gate15066(.O (g26887), .I1 (g26542), .I2 (g24193));
OR2X1 gate15067(.O (g28729), .I1 (g27502), .I2 (g16732));
OR2X1 gate15068(.O (g28577), .I1 (g27326), .I2 (g26272));
OR2X1 gate15069(.O (g24510), .I1 (g22488), .I2 (g7567));
OR2X1 gate15070(.O (g30432), .I1 (g29888), .I2 (g21816));
OR2X1 gate15071(.O (g28728), .I1 (g27501), .I2 (g16730));
OR2X1 gate15072(.O (g29262), .I1 (g28327), .I2 (g18608));
OR2X1 gate15073(.O (g27542), .I1 (g16190), .I2 (g26094));
OR2X1 gate15074(.O (g27453), .I1 (g25976), .I2 (g24606));
OR2X1 gate15075(.O (g23383), .I1 (g19756), .I2 (g16222));
OR2X1 gate15076(.O (g24578), .I1 (g2882), .I2 (g23825));
OR2X1 gate15077(.O (g30461), .I1 (g30219), .I2 (g21932));
OR2X1 gate15078(.O (g30342), .I1 (g29330), .I2 (g18261));
OR2X1 gate15079(.O (g34461), .I1 (g34291), .I2 (g18681));
OR2X1 gate15080(.O (g26365), .I1 (g25504), .I2 (g25141));
OR3X1 gate15081(.O (I18452), .I1 (g14514), .I2 (g14448), .I3 (g14418));
OR2X1 gate15082(.O (g26960), .I1 (g26258), .I2 (g24304));
OR2X1 gate15083(.O (g34031), .I1 (g33735), .I2 (g18705));
OR2X1 gate15084(.O (g31472), .I1 (g29642), .I2 (g28352));
OR2X1 gate15085(.O (g28083), .I1 (g27249), .I2 (g18689));
OR2X1 gate15086(.O (g28348), .I1 (g27139), .I2 (g15823));
OR2X1 gate15087(.O (g34199), .I1 (g33820), .I2 (g33828));
OR2X1 gate15088(.O (g32280), .I1 (g24790), .I2 (g31225));
OR2X1 gate15089(.O (g9984), .I1 (g4300), .I2 (g4242));
OR2X1 gate15090(.O (g34887), .I1 (g34865), .I2 (g21670));
OR2X1 gate15091(.O (g31911), .I1 (g31784), .I2 (g21969));
OR2X1 gate15092(.O (g30529), .I1 (g30212), .I2 (g22075));
OR2X1 gate15093(.O (g33628), .I1 (g33071), .I2 (g32450));
OR2X1 gate15094(.O (g27274), .I1 (g15779), .I2 (g25915));
OR2X1 gate15095(.O (g31246), .I1 (g25965), .I2 (g29518));
OR2X1 gate15096(.O (g25611), .I1 (g24931), .I2 (g18128));
OR2X1 gate15097(.O (g19356), .I1 (g17784), .I2 (g14874));
OR2X1 gate15098(.O (g25722), .I1 (g25530), .I2 (g18768));
OR2X1 gate15099(.O (g28622), .I1 (g27360), .I2 (g16519));
OR2X1 gate15100(.O (g28566), .I1 (g27316), .I2 (g26254));
OR2X1 gate15101(.O (g30528), .I1 (g30202), .I2 (g22074));
OR2X1 gate15102(.O (g9483), .I1 (g1008), .I2 (g969));
OR2X1 gate15103(.O (g30393), .I1 (g29986), .I2 (g21748));
OR2X1 gate15104(.O (g27122), .I1 (g22537), .I2 (g25917));
OR2X1 gate15105(.O (g34843), .I1 (g33924), .I2 (g34782));
OR2X1 gate15106(.O (g34330), .I1 (g34069), .I2 (g33717));
OR2X1 gate15107(.O (g30365), .I1 (g30158), .I2 (g18412));
OR2X1 gate15108(.O (g24275), .I1 (g23474), .I2 (g18645));
OR2X1 gate15109(.O (g29247), .I1 (g28694), .I2 (g18410));
OR2X1 gate15110(.O (g31591), .I1 (g29358), .I2 (g29353));
OR2X1 gate15111(.O (g31785), .I1 (g30071), .I2 (g30082));
OR2X1 gate15112(.O (g33591), .I1 (g33082), .I2 (g18474));
OR2X1 gate15113(.O (g24430), .I1 (g23151), .I2 (g8234));
OR2X1 gate15114(.O (g24746), .I1 (g22588), .I2 (g19461));
OR2X1 gate15115(.O (g32231), .I1 (g30590), .I2 (g29346));
OR2X1 gate15116(.O (g25753), .I1 (g25165), .I2 (g22100));
OR2X1 gate15117(.O (g31754), .I1 (g29989), .I2 (g30006));
OR2X1 gate15118(.O (g28138), .I1 (g27964), .I2 (g27968));
OR2X1 gate15119(.O (g24237), .I1 (g22515), .I2 (g18242));
OR2X1 gate15120(.O (g33950), .I1 (g32450), .I2 (g33460));
OR2X1 gate15121(.O (g29777), .I1 (g28227), .I2 (g28234));
OR2X1 gate15122(.O (g24340), .I1 (g24016), .I2 (g18770));
OR2X1 gate15123(.O (g25650), .I1 (g24663), .I2 (g21743));
OR2X1 gate15124(.O (g25736), .I1 (g25536), .I2 (g18785));
OR2X1 gate15125(.O (g29251), .I1 (g28679), .I2 (g18464));
OR2X1 gate15126(.O (g29272), .I1 (g28346), .I2 (g18638));
OR2X1 gate15127(.O (g28636), .I1 (g27376), .I2 (g16538));
OR2X1 gate15128(.O (g19449), .I1 (g15567), .I2 (g12939));
OR2X1 gate15129(.O (g28852), .I1 (g27559), .I2 (g16871));
OR2X1 gate15130(.O (g34259), .I1 (g34066), .I2 (g18679));
OR2X1 gate15131(.O (g30471), .I1 (g30175), .I2 (g21942));
OR2X1 gate15132(.O (g33996), .I1 (g33862), .I2 (g18426));
OR2X1 gate15133(.O (g34708), .I1 (g33381), .I2 (g34572));
OR4X1 gate15134(.O (g26657), .I1 (g24908), .I2 (g24900), .I3 (g24887), .I4 (g24861));
OR2X1 gate15135(.O (g25696), .I1 (g25012), .I2 (g21915));
OR2X1 gate15136(.O (g26955), .I1 (g26391), .I2 (g24293));
OR2X1 gate15137(.O (g34258), .I1 (g34211), .I2 (g18675));
OR2X1 gate15138(.O (g24517), .I1 (g22158), .I2 (g18906));
OR2X1 gate15139(.O (g26879), .I1 (g25580), .I2 (g25581));
OR2X1 gate15140(.O (g26970), .I1 (g26308), .I2 (g24332));
OR2X1 gate15141(.O (g25764), .I1 (g25551), .I2 (g18819));
OR2X1 gate15142(.O (g28664), .I1 (g27408), .I2 (g16613));
OR2X1 gate15143(.O (g26878), .I1 (g25578), .I2 (g25579));
OR2X1 gate15144(.O (g16867), .I1 (g13493), .I2 (g11045));
OR2X1 gate15145(.O (g25960), .I1 (g24566), .I2 (g24678));
OR2X1 gate15146(.O (g34043), .I1 (g33903), .I2 (g33905));
OR2X1 gate15147(.O (g26886), .I1 (g26651), .I2 (g24192));
OR2X1 gate15148(.O (g25868), .I1 (g25450), .I2 (g23885));
OR2X1 gate15149(.O (g28576), .I1 (g27325), .I2 (g26271));
OR2X1 gate15150(.O (g31319), .I1 (g29612), .I2 (g28324));
OR2X1 gate15151(.O (g27575), .I1 (g26147), .I2 (g24731));
OR2X1 gate15152(.O (g26967), .I1 (g26350), .I2 (g24319));
OR2X1 gate15153(.O (g33318), .I1 (g31969), .I2 (g32434));
OR2X1 gate15154(.O (g34602), .I1 (g34489), .I2 (g18269));
OR2X1 gate15155(.O (g25709), .I1 (g25014), .I2 (g21960));
OR2X1 gate15156(.O (g30375), .I1 (g30149), .I2 (g18466));
OR2X1 gate15157(.O (g34657), .I1 (g33114), .I2 (g34497));
OR2X1 gate15158(.O (g28609), .I1 (g27346), .I2 (g16483));
OR2X1 gate15159(.O (g33227), .I1 (g32029), .I2 (g32031));
OR2X1 gate15160(.O (g9536), .I1 (g1351), .I2 (g1312));
OR2X1 gate15161(.O (g33059), .I1 (g31987), .I2 (g22021));
OR2X1 gate15162(.O (g33025), .I1 (g32162), .I2 (g21780));
OR2X1 gate15163(.O (g25708), .I1 (g25526), .I2 (g18751));
OR2X1 gate15164(.O (g34970), .I1 (g34868), .I2 (g34961));
OR4X1 gate15165(.O (I29986), .I1 (g31070), .I2 (g31194), .I3 (g30614), .I4 (g30673));
OR2X1 gate15166(.O (g23822), .I1 (g20218), .I2 (g16929));
OR2X1 gate15167(.O (g33540), .I1 (g33099), .I2 (g18207));
OR2X1 gate15168(.O (g27108), .I1 (g22522), .I2 (g25911));
OR2X1 gate15169(.O (g33058), .I1 (g31976), .I2 (g22020));
OR2X1 gate15170(.O (g30337), .I1 (g29334), .I2 (g18220));
OR2X1 gate15171(.O (g32243), .I1 (g31166), .I2 (g29683));
OR2X1 gate15172(.O (g26919), .I1 (g25951), .I2 (g18267));
OR2X1 gate15173(.O (g28052), .I1 (g27710), .I2 (g18167));
OR2X1 gate15174(.O (g27283), .I1 (g25922), .I2 (g25924));
OR2X1 gate15175(.O (g26918), .I1 (g25931), .I2 (g18243));
OR2X1 gate15176(.O (g28745), .I1 (g27519), .I2 (g16760));
OR2X1 gate15177(.O (g15968), .I1 (g13038), .I2 (g10677));
OR4X1 gate15178(.O (I31854), .I1 (g33492), .I2 (g33493), .I3 (g33494), .I4 (g33495));
OR2X1 gate15179(.O (g33044), .I1 (g32199), .I2 (g24327));
OR2X1 gate15180(.O (g34792), .I1 (g34750), .I2 (g18569));
OR2X1 gate15181(.O (g32268), .I1 (g24785), .I2 (g31219));
OR2X1 gate15182(.O (g23194), .I1 (g19564), .I2 (g19578));
OR2X1 gate15183(.O (g33281), .I1 (g32142), .I2 (g29576));
OR2X1 gate15184(.O (g31902), .I1 (g31744), .I2 (g21910));
OR2X1 gate15185(.O (g30459), .I1 (g29314), .I2 (g21926));
OR2X1 gate15186(.O (g30425), .I1 (g29770), .I2 (g21809));
OR3X1 gate15187(.O (g33957), .I1 (g33523), .I2 (I31868), .I3 (I31869));
OR2X1 gate15188(.O (g24347), .I1 (g23754), .I2 (g18790));
OR2X1 gate15189(.O (g34459), .I1 (g34415), .I2 (g18673));
OR2X1 gate15190(.O (g25602), .I1 (g24673), .I2 (g18113));
OR2X1 gate15191(.O (g12982), .I1 (g12220), .I2 (g9968));
OR2X1 gate15192(.O (g25657), .I1 (g24624), .I2 (g21782));
OR2X1 gate15193(.O (g24253), .I1 (g22525), .I2 (g18300));
OR2X1 gate15194(.O (g25774), .I1 (g25223), .I2 (g12043));
OR2X1 gate15195(.O (g29246), .I1 (g28710), .I2 (g18406));
OR2X1 gate15196(.O (g30458), .I1 (g30005), .I2 (g24330));
OR2X1 gate15197(.O (g34458), .I1 (g34396), .I2 (g18671));
OR2X1 gate15198(.O (g33562), .I1 (g33414), .I2 (g18379));
OR2X1 gate15199(.O (g34010), .I1 (g33872), .I2 (g18478));
OR2X1 gate15200(.O (g24236), .I1 (g22489), .I2 (g18241));
OR2X1 gate15201(.O (g25878), .I1 (g25503), .I2 (g23920));
OR2X1 gate15202(.O (g28732), .I1 (g27505), .I2 (g16734));
OR2X1 gate15203(.O (g33699), .I1 (g32409), .I2 (g33433));
OR2X1 gate15204(.O (g32993), .I1 (g32255), .I2 (g18352));
OR2X1 gate15205(.O (g30545), .I1 (g30268), .I2 (g22116));
OR2X1 gate15206(.O (g30444), .I1 (g29901), .I2 (g21853));
OR2X1 gate15207(.O (g29776), .I1 (g28225), .I2 (g22846));
OR3X1 gate15208(.O (g24952), .I1 (g21326), .I2 (g21340), .I3 (I24117));
OR2X1 gate15209(.O (g24351), .I1 (g23774), .I2 (g18807));
OR2X1 gate15210(.O (g33290), .I1 (g32149), .I2 (g29589));
OR2X1 gate15211(.O (g26901), .I1 (g26362), .I2 (g24218));
OR2X1 gate15212(.O (g34444), .I1 (g34389), .I2 (g18546));
OR2X1 gate15213(.O (g24821), .I1 (g21404), .I2 (g23990));
OR2X1 gate15214(.O (g29754), .I1 (g28215), .I2 (g28218));
OR2X1 gate15215(.O (g34599), .I1 (g34542), .I2 (g18149));
OR2X1 gate15216(.O (g32131), .I1 (g24495), .I2 (g30926));
OR2X1 gate15217(.O (g20063), .I1 (g15978), .I2 (g13313));
OR2X1 gate15218(.O (g34598), .I1 (g34541), .I2 (g18136));
OR2X1 gate15219(.O (g15910), .I1 (g13025), .I2 (g10654));
OR2X1 gate15220(.O (g24264), .I1 (g22310), .I2 (g18559));
OR2X1 gate15221(.O (g23276), .I1 (g19681), .I2 (g16161));
OR2X1 gate15222(.O (g27663), .I1 (g26323), .I2 (g24820));
OR2X1 gate15223(.O (g28400), .I1 (g27211), .I2 (g15870));
OR2X1 gate15224(.O (g32210), .I1 (g31123), .I2 (g29600));
OR2X1 gate15225(.O (g21900), .I1 (g20977), .I2 (g15114));
OR2X1 gate15226(.O (g16866), .I1 (g13492), .I2 (g11044));
OR2X1 gate15227(.O (g28329), .I1 (g27128), .I2 (g15813));
OR2X1 gate15228(.O (g30532), .I1 (g30193), .I2 (g22078));
OR2X1 gate15229(.O (g32279), .I1 (g31220), .I2 (g31224));
OR2X1 gate15230(.O (g34125), .I1 (g33724), .I2 (g33124));
OR2X1 gate15231(.O (g22652), .I1 (g18992), .I2 (g15653));
OR2X1 gate15232(.O (g13762), .I1 (g499), .I2 (g12527));
OR2X1 gate15233(.O (g34977), .I1 (g34873), .I2 (g34966));
OR2X1 gate15234(.O (g25010), .I1 (g23267), .I2 (g2932));
OR2X1 gate15235(.O (g31895), .I1 (g31505), .I2 (g24296));
OR2X1 gate15236(.O (g28328), .I1 (g27127), .I2 (g15812));
OR2X1 gate15237(.O (g33547), .I1 (g33349), .I2 (g18331));
OR2X1 gate15238(.O (g34158), .I1 (g33784), .I2 (g19740));
OR2X1 gate15239(.O (g24209), .I1 (g23415), .I2 (g18122));
OR2X1 gate15240(.O (g34783), .I1 (g33110), .I2 (g34667));
OR2X1 gate15241(.O (g28538), .I1 (g27294), .I2 (g26206));
OR2X1 gate15242(.O (g26966), .I1 (g26345), .I2 (g24318));
OR2X1 gate15243(.O (g25545), .I1 (g23551), .I2 (g20658));
OR2X1 gate15244(.O (g30561), .I1 (g30284), .I2 (g22132));
OR2X1 gate15245(.O (g7673), .I1 (g4153), .I2 (g4172));
OR2X1 gate15246(.O (g30353), .I1 (g30095), .I2 (g18355));
OR2X1 gate15247(.O (g24208), .I1 (g23404), .I2 (g18121));
OR2X1 gate15248(.O (g25599), .I1 (g24914), .I2 (g21721));
OR2X1 gate15249(.O (g34353), .I1 (g26088), .I2 (g34114));
OR2X1 gate15250(.O (g29319), .I1 (g28812), .I2 (g14453));
OR2X1 gate15251(.O (g25598), .I1 (g24904), .I2 (g21720));
OR2X1 gate15252(.O (g33551), .I1 (g33446), .I2 (g18342));
OR2X1 gate15253(.O (g33572), .I1 (g33339), .I2 (g18414));
OR2X1 gate15254(.O (g30336), .I1 (g29324), .I2 (g18203));
OR2X1 gate15255(.O (g29227), .I1 (g28456), .I2 (g18169));
OR2X1 gate15256(.O (g13543), .I1 (g10543), .I2 (g10565));
OR4X1 gate15257(.O (I31839), .I1 (g33465), .I2 (g33466), .I3 (g33467), .I4 (g33468));
OR4X1 gate15258(.O (I31838), .I1 (g33461), .I2 (g33462), .I3 (g33463), .I4 (g33464));
OR2X1 gate15259(.O (g28100), .I1 (g27690), .I2 (g22051));
OR2X1 gate15260(.O (g20905), .I1 (g7216), .I2 (g17264));
OR2X1 gate15261(.O (g34631), .I1 (g34562), .I2 (g15118));
OR2X1 gate15262(.O (g30364), .I1 (g30086), .I2 (g18411));
OR2X1 gate15263(.O (g34017), .I1 (g33880), .I2 (g18504));
OR2X1 gate15264(.O (g24274), .I1 (g23187), .I2 (g18631));
OR2X1 gate15265(.O (g13242), .I1 (g11336), .I2 (g7601));
OR3X1 gate15266(.O (g33956), .I1 (g33514), .I2 (I31863), .I3 (I31864));
OR2X1 gate15267(.O (g24346), .I1 (g23725), .I2 (g18789));
OR2X1 gate15268(.O (g33297), .I1 (g32157), .I2 (g29621));
OR2X1 gate15269(.O (g25656), .I1 (g24945), .I2 (g18609));
OR2X1 gate15270(.O (g31889), .I1 (g31118), .I2 (g21822));
OR2X1 gate15271(.O (g33980), .I1 (g33843), .I2 (g18370));
OR2X1 gate15272(.O (g24565), .I1 (g22309), .I2 (g19275));
OR2X1 gate15273(.O (g21892), .I1 (g19788), .I2 (g15104));
OR2X1 gate15274(.O (g25680), .I1 (g24794), .I2 (g21839));
OR3X1 gate15275(.O (g16876), .I1 (g14028), .I2 (g11773), .I3 (g11755));
OR2X1 gate15276(.O (g29281), .I1 (g28541), .I2 (g18743));
OR2X1 gate15277(.O (g31888), .I1 (g31067), .I2 (g21821));
OR2X1 gate15278(.O (g20034), .I1 (g15902), .I2 (g13299));
OR2X1 gate15279(.O (g29301), .I1 (g28686), .I2 (g18797));
OR2X1 gate15280(.O (g27509), .I1 (g26023), .I2 (g24640));
OR2X1 gate15281(.O (g34289), .I1 (g26847), .I2 (g34218));
OR2X1 gate15282(.O (g24641), .I1 (g22151), .I2 (g22159));
OR2X1 gate15283(.O (g34023), .I1 (g33796), .I2 (g24320));
OR2X1 gate15284(.O (g34288), .I1 (g26846), .I2 (g34217));
OR2X1 gate15285(.O (g32217), .I1 (g31129), .I2 (g29616));
OR2X1 gate15286(.O (g26954), .I1 (g26380), .I2 (g24292));
OR3X1 gate15287(.O (I18449), .I1 (g14512), .I2 (g14445), .I3 (g14415));
OR2X1 gate15288(.O (g31931), .I1 (g31494), .I2 (g22095));
OR2X1 gate15289(.O (g29290), .I1 (g28569), .I2 (g18764));
OR2X1 gate15290(.O (g25631), .I1 (g24554), .I2 (g18275));
OR2X1 gate15291(.O (g30495), .I1 (g30222), .I2 (g21991));
OR2X1 gate15292(.O (g32223), .I1 (g31142), .I2 (g29637));
OR2X1 gate15293(.O (g29366), .I1 (g13738), .I2 (g28439));
OR2X1 gate15294(.O (g27574), .I1 (g26145), .I2 (g24730));
OR2X1 gate15295(.O (g34976), .I1 (g34872), .I2 (g34965));
OR2X1 gate15296(.O (g26392), .I1 (g24745), .I2 (g23050));
OR2X1 gate15297(.O (g27205), .I1 (g25833), .I2 (g24421));
OR2X1 gate15298(.O (g33546), .I1 (g33402), .I2 (g18327));
OR2X1 gate15299(.O (g30374), .I1 (g30078), .I2 (g18465));
OR2X1 gate15300(.O (g16076), .I1 (g13081), .I2 (g10736));
OR2X1 gate15301(.O (g34374), .I1 (g26294), .I2 (g34139));
OR4X1 gate15302(.O (I30728), .I1 (g32345), .I2 (g32350), .I3 (g32056), .I4 (g32018));
OR2X1 gate15303(.O (g33024), .I1 (g32324), .I2 (g21752));
OR2X1 gate15304(.O (g34643), .I1 (g34554), .I2 (g18752));
OR2X1 gate15305(.O (g28435), .I1 (g27234), .I2 (g15967));
OR2X1 gate15306(.O (g28082), .I1 (g27369), .I2 (g24315));
OR2X1 gate15307(.O (g26893), .I1 (g26753), .I2 (g24199));
OR2X1 gate15308(.O (g29226), .I1 (g28455), .I2 (g18159));
OR2X1 gate15309(.O (g28744), .I1 (g27518), .I2 (g16759));
OR2X1 gate15310(.O (g34260), .I1 (g34113), .I2 (g18680));
OR2X1 gate15311(.O (g28345), .I1 (g27137), .I2 (g15821));
OR2X1 gate15312(.O (g29481), .I1 (g28117), .I2 (g28125));
OR2X1 gate15313(.O (g30392), .I1 (g30091), .I2 (g18558));
OR2X1 gate15314(.O (g30489), .I1 (g30250), .I2 (g21985));
OR2X1 gate15315(.O (g33625), .I1 (g33373), .I2 (g18809));
OR2X1 gate15316(.O (g32373), .I1 (g29894), .I2 (g31321));
OR2X1 gate15317(.O (g33987), .I1 (g33847), .I2 (g18396));
OR2X1 gate15318(.O (g31250), .I1 (g25972), .I2 (g29526));
OR2X1 gate15319(.O (g25687), .I1 (g24729), .I2 (g21882));
OR2X1 gate15320(.O (g30559), .I1 (g30269), .I2 (g22130));
OR2X1 gate15321(.O (g30525), .I1 (g30266), .I2 (g22071));
OR2X1 gate15322(.O (g30488), .I1 (g30197), .I2 (g21984));
OR2X1 gate15323(.O (g30424), .I1 (g29760), .I2 (g21808));
OR2X1 gate15324(.O (g25752), .I1 (g25079), .I2 (g22099));
OR2X1 gate15325(.O (g34016), .I1 (g33867), .I2 (g18503));
OR2X1 gate15326(.O (g30558), .I1 (g30258), .I2 (g22129));
OR2X1 gate15327(.O (g27152), .I1 (g24393), .I2 (g25817));
OR2X1 gate15328(.O (g33296), .I1 (g32156), .I2 (g29617));
OR2X1 gate15329(.O (g25643), .I1 (g24602), .I2 (g21736));
OR2X1 gate15330(.O (g29490), .I1 (g25832), .I2 (g28136));
OR2X1 gate15331(.O (g16839), .I1 (g13473), .I2 (g11035));
OR2X1 gate15332(.O (g28332), .I1 (g27130), .I2 (g15815));
OR2X1 gate15333(.O (g30544), .I1 (g30257), .I2 (g22115));
OR2X1 gate15334(.O (g33969), .I1 (g33864), .I2 (g18321));
OR2X1 gate15335(.O (g25669), .I1 (g24657), .I2 (g18624));
OR2X1 gate15336(.O (g28135), .I1 (g27959), .I2 (g27963));
OR2X1 gate15337(.O (g29297), .I1 (g28683), .I2 (g18784));
OR2X1 gate15338(.O (g33060), .I1 (g31992), .I2 (g22022));
OR2X1 gate15339(.O (g33968), .I1 (g33855), .I2 (g18320));
OR2X1 gate15340(.O (g26939), .I1 (g25907), .I2 (g21884));
OR2X1 gate15341(.O (g25668), .I1 (g24646), .I2 (g18623));
OR3X1 gate15342(.O (g33197), .I1 (g32342), .I2 (I30745), .I3 (I30746));
OR2X1 gate15343(.O (g28361), .I1 (g27153), .I2 (g15839));
OR2X1 gate15344(.O (g32216), .I1 (g31128), .I2 (g29615));
OR2X1 gate15345(.O (g27405), .I1 (g24572), .I2 (g25968));
OR2X1 gate15346(.O (g26938), .I1 (g26186), .I2 (g21883));
OR2X1 gate15347(.O (g31870), .I1 (g30607), .I2 (g18262));
OR3X1 gate15348(.O (I28147), .I1 (g2946), .I2 (g24561), .I3 (g28220));
OR2X1 gate15349(.O (g24840), .I1 (g21419), .I2 (g23996));
OR2X1 gate15350(.O (g34610), .I1 (g34507), .I2 (g18564));
OR2X1 gate15351(.O (g24390), .I1 (g23779), .I2 (g21285));
OR2X1 gate15352(.O (g30189), .I1 (g23401), .I2 (g28543));
OR2X1 gate15353(.O (g28049), .I1 (g27684), .I2 (g18164));
OR2X1 gate15354(.O (g34255), .I1 (g34120), .I2 (g24302));
OR2X1 gate15355(.O (g34189), .I1 (g33801), .I2 (g33808));
OR2X1 gate15356(.O (g30270), .I1 (g28624), .I2 (g27664));
OR2X1 gate15357(.O (g28048), .I1 (g27362), .I2 (g18163));
OR2X1 gate15358(.O (g20522), .I1 (g691), .I2 (g16893));
OR2X1 gate15359(.O (g26875), .I1 (g21652), .I2 (g25575));
OR2X1 gate15360(.O (g32117), .I1 (g24482), .I2 (g30914));
OR4X1 gate15361(.O (I23163), .I1 (g20982), .I2 (g21127), .I3 (g21193), .I4 (g21256));
OR2X1 gate15362(.O (g31894), .I1 (g30671), .I2 (g21870));
OR2X1 gate15363(.O (g31867), .I1 (g31238), .I2 (g18175));
OR2X1 gate15364(.O (g30460), .I1 (g30207), .I2 (g21931));
OR2X1 gate15365(.O (g30383), .I1 (g30138), .I2 (g18513));
OR2X1 gate15366(.O (g34460), .I1 (g34301), .I2 (g18677));
OR2X1 gate15367(.O (g30093), .I1 (g28467), .I2 (g11397));
OR2X1 gate15368(.O (g34030), .I1 (g33727), .I2 (g18704));
OR2X1 gate15369(.O (g25713), .I1 (g25147), .I2 (g21964));
OR2X1 gate15370(.O (g28613), .I1 (g27350), .I2 (g26310));
OR2X1 gate15371(.O (g33581), .I1 (g33333), .I2 (g18443));
OR2X1 gate15372(.O (g33714), .I1 (g32419), .I2 (g33450));
OR4X1 gate15373(.O (g29520), .I1 (g28291), .I2 (g28281), .I3 (g28264), .I4 (g28254));
OR2X1 gate15374(.O (g34267), .I1 (g34079), .I2 (g18728));
OR2X1 gate15375(.O (g34294), .I1 (g26855), .I2 (g34225));
OR2X1 gate15376(.O (g31315), .I1 (g29607), .I2 (g29623));
OR2X1 gate15377(.O (g33315), .I1 (g29665), .I2 (g32175));
OR2X1 gate15378(.O (g31910), .I1 (g31471), .I2 (g21957));
OR2X1 gate15379(.O (g13006), .I1 (g12284), .I2 (g10034));
OR2X1 gate15380(.O (g25610), .I1 (g24923), .I2 (g18127));
OR2X1 gate15381(.O (g31257), .I1 (g29531), .I2 (g28253));
OR2X1 gate15382(.O (g25705), .I1 (g25069), .I2 (g18744));
OR2X1 gate15383(.O (g28605), .I1 (g27341), .I2 (g26302));
OR2X1 gate15384(.O (g33257), .I1 (g32108), .I2 (g29519));
OR2X1 gate15385(.O (g32123), .I1 (g30915), .I2 (g30919));
OR2X1 gate15386(.O (g33979), .I1 (g33942), .I2 (g18361));
OR2X1 gate15387(.O (g33055), .I1 (g31986), .I2 (g21976));
OR2X1 gate15388(.O (g16187), .I1 (g8822), .I2 (g13486));
OR2X1 gate15389(.O (g25679), .I1 (g24728), .I2 (g21836));
OR2X1 gate15390(.O (g33070), .I1 (g32010), .I2 (g22114));
OR2X1 gate15391(.O (g33978), .I1 (g33892), .I2 (g18356));
OR2X1 gate15392(.O (g25678), .I1 (g24709), .I2 (g21835));
OR2X1 gate15393(.O (g26915), .I1 (g25900), .I2 (g18230));
OR2X1 gate15394(.O (g33590), .I1 (g33358), .I2 (g18470));
OR2X1 gate15395(.O (g15965), .I1 (g13035), .I2 (g10675));
OR2X1 gate15396(.O (g28371), .I1 (g27177), .I2 (g15847));
OR4X1 gate15397(.O (I30745), .I1 (g31777), .I2 (g32321), .I3 (g32069), .I4 (g32084));
OR2X1 gate15398(.O (g32230), .I1 (g30589), .I2 (g29345));
OR2X1 gate15399(.O (g33986), .I1 (g33639), .I2 (g18387));
OR2X1 gate15400(.O (g24252), .I1 (g22518), .I2 (g18299));
OR2X1 gate15401(.O (g25686), .I1 (g24712), .I2 (g21881));
OR2X1 gate15402(.O (g33384), .I1 (g32248), .I2 (g29943));
OR2X1 gate15403(.O (g33067), .I1 (g31989), .I2 (g22111));
OR2X1 gate15404(.O (g12768), .I1 (g7785), .I2 (g7202));
OR2X1 gate15405(.O (g29250), .I1 (g28695), .I2 (g18460));
OR2X1 gate15406(.O (g32992), .I1 (g32242), .I2 (g18351));
OR2X1 gate15407(.O (g32391), .I1 (g31502), .I2 (g29982));
OR2X1 gate15408(.O (g30455), .I1 (g30041), .I2 (g21864));
OR2X1 gate15409(.O (g34455), .I1 (g34284), .I2 (g18668));
OR3X1 gate15410(.O (g11372), .I1 (g490), .I2 (g482), .I3 (g8038));
OR2X1 gate15411(.O (g31877), .I1 (g31278), .I2 (g21732));
OR2X1 gate15412(.O (g30470), .I1 (g30165), .I2 (g21941));
OR2X1 gate15413(.O (g34617), .I1 (g34526), .I2 (g18579));
OR2X1 gate15414(.O (g22648), .I1 (g18987), .I2 (g15652));
OR3X1 gate15415(.O (I12611), .I1 (g1500), .I2 (g1582), .I3 (g1333));
OR2X1 gate15416(.O (g29296), .I1 (g28586), .I2 (g18781));
OR2X1 gate15417(.O (g33019), .I1 (g32339), .I2 (g18536));
OR2X1 gate15418(.O (g30201), .I1 (g23412), .I2 (g28557));
OR2X1 gate15419(.O (g33018), .I1 (g32312), .I2 (g18525));
OR4X1 gate15420(.O (I30761), .I1 (g32071), .I2 (g32167), .I3 (g32067), .I4 (g32082));
OR2X1 gate15421(.O (g30467), .I1 (g30185), .I2 (g21938));
OR2X1 gate15422(.O (g30494), .I1 (g30209), .I2 (g21990));
OR2X1 gate15423(.O (g34467), .I1 (g34341), .I2 (g18717));
OR2X1 gate15424(.O (g34494), .I1 (g26849), .I2 (g34413));
OR2X1 gate15425(.O (g29197), .I1 (g27187), .I2 (g27163));
OR2X1 gate15426(.O (g34623), .I1 (g34525), .I2 (g18585));
OR2X1 gate15427(.O (g34037), .I1 (g33803), .I2 (g18734));
OR4X1 gate15428(.O (I30400), .I1 (g31021), .I2 (g30937), .I3 (g31327), .I4 (g30614));
OR2X1 gate15429(.O (g27248), .I1 (g24880), .I2 (g25953));
OR2X1 gate15430(.O (g30984), .I1 (g29765), .I2 (g29755));
OR2X1 gate15431(.O (g27552), .I1 (g26092), .I2 (g24676));
OR2X1 gate15432(.O (g31917), .I1 (g31478), .I2 (g22003));
OR2X1 gate15433(.O (g30419), .I1 (g29759), .I2 (g21803));
OR2X1 gate15434(.O (g31866), .I1 (g31252), .I2 (g18142));
OR2X1 gate15435(.O (g30352), .I1 (g30094), .I2 (g18340));
OR2X1 gate15436(.O (g27779), .I1 (g17317), .I2 (g26694));
OR2X1 gate15437(.O (g25617), .I1 (g25466), .I2 (g18189));
OR2X1 gate15438(.O (g24213), .I1 (g23220), .I2 (g18186));
OR3X1 gate15439(.O (g23184), .I1 (g20198), .I2 (g20185), .I3 (I22280));
OR2X1 gate15440(.O (g28724), .I1 (g27491), .I2 (g16707));
OR2X1 gate15441(.O (g34352), .I1 (g26079), .I2 (g34109));
OR2X1 gate15442(.O (g28359), .I1 (g27151), .I2 (g15838));
OR2X1 gate15443(.O (g30418), .I1 (g29751), .I2 (g21802));
OR2X1 gate15444(.O (g32275), .I1 (g31210), .I2 (g29732));
OR2X1 gate15445(.O (g31001), .I1 (g29360), .I2 (g28151));
OR2X1 gate15446(.O (g28358), .I1 (g27149), .I2 (g15837));
OR2X1 gate15447(.O (g34266), .I1 (g34076), .I2 (g18719));
OR2X1 gate15448(.O (g33001), .I1 (g32282), .I2 (g18404));
OR2X1 gate15449(.O (g34170), .I1 (g33790), .I2 (g19855));
OR2X1 gate15450(.O (g24205), .I1 (g23006), .I2 (g18109));
OR2X1 gate15451(.O (g33706), .I1 (g32412), .I2 (g33440));
OR2X1 gate15452(.O (g33597), .I1 (g33344), .I2 (g18495));
OR2X1 gate15453(.O (g32237), .I1 (g31153), .I2 (g29667));
OR2X1 gate15454(.O (g31256), .I1 (g25983), .I2 (g29537));
OR2X1 gate15455(.O (g33256), .I1 (g32107), .I2 (g29517));
OR2X1 gate15456(.O (g25595), .I1 (g24835), .I2 (g21717));
OR2X1 gate15457(.O (g31923), .I1 (g31763), .I2 (g22048));
OR2X1 gate15458(.O (g32983), .I1 (g31990), .I2 (g18222));
OR2X1 gate15459(.O (g19879), .I1 (g15841), .I2 (g13265));
OR2X1 gate15460(.O (g28344), .I1 (g27136), .I2 (g15820));
OR2X1 gate15461(.O (g22832), .I1 (g19354), .I2 (g15722));
OR2X1 gate15462(.O (g33280), .I1 (g32141), .I2 (g29574));
OR2X1 gate15463(.O (g25623), .I1 (g24552), .I2 (g18219));
OR2X1 gate15464(.O (g20051), .I1 (g15936), .I2 (g13306));
OR2X1 gate15465(.O (g25037), .I1 (g23103), .I2 (g19911));
OR2X1 gate15466(.O (g33624), .I1 (g33371), .I2 (g18808));
OR2X1 gate15467(.O (g34167), .I1 (g33786), .I2 (g19768));
OR2X1 gate15468(.O (g34194), .I1 (g33811), .I2 (g33815));
OR4X1 gate15469(.O (g26616), .I1 (g24881), .I2 (g24855), .I3 (g24843), .I4 (g24822));
OR2X1 gate15470(.O (g19337), .I1 (g17770), .I2 (g17785));
OR2X1 gate15471(.O (g28682), .I1 (g27430), .I2 (g16635));
OR2X1 gate15472(.O (g29257), .I1 (g28228), .I2 (g18600));
OR4X1 gate15473(.O (I23755), .I1 (g22904), .I2 (g22927), .I3 (g22980), .I4 (g23444));
OR2X1 gate15474(.O (g30524), .I1 (g30255), .I2 (g22070));
OR2X1 gate15475(.O (g27233), .I1 (g25876), .I2 (g24451));
OR2X1 gate15476(.O (g16800), .I1 (g13436), .I2 (g11027));
OR2X1 gate15477(.O (g29496), .I1 (g28567), .I2 (g27615));
OR2X1 gate15478(.O (g27182), .I1 (g25818), .I2 (g24410));
OR2X1 gate15479(.O (g30401), .I1 (g29782), .I2 (g21760));
OR2X1 gate15480(.O (g30477), .I1 (g30239), .I2 (g21948));
OR2X1 gate15481(.O (g26305), .I1 (g24556), .I2 (g24564));
OR2X1 gate15482(.O (g24350), .I1 (g23755), .I2 (g18806));
OR2X1 gate15483(.O (g26809), .I1 (g24930), .I2 (g24939));
OR2X1 gate15484(.O (g33066), .I1 (g32341), .I2 (g22096));
OR2X1 gate15485(.O (g26900), .I1 (g26819), .I2 (g24217));
OR2X1 gate15486(.O (g33231), .I1 (g32032), .I2 (g32036));
OR2X1 gate15487(.O (g29741), .I1 (g28205), .I2 (g15883));
OR2X1 gate15488(.O (g32130), .I1 (g30921), .I2 (g30925));
OR2X1 gate15489(.O (g34022), .I1 (g33873), .I2 (g18538));
OR2X1 gate15490(.O (g28134), .I1 (g27958), .I2 (g27962));
OR2X1 gate15491(.O (g31876), .I1 (g31125), .I2 (g21731));
OR2X1 gate15492(.O (g31885), .I1 (g31017), .I2 (g21779));
OR2X1 gate15493(.O (g32362), .I1 (g29870), .I2 (g31301));
OR2X1 gate15494(.O (g34616), .I1 (g34519), .I2 (g18577));
OR2X1 gate15495(.O (g25589), .I1 (g21690), .I2 (g24159));
OR2X1 gate15496(.O (g29801), .I1 (g25987), .I2 (g28251));
OR2X1 gate15497(.O (g29735), .I1 (g28202), .I2 (g10898));
OR2X1 gate15498(.O (g25588), .I1 (g21686), .I2 (g24158));
OR2X1 gate15499(.O (g34305), .I1 (g25775), .I2 (g34050));
OR2X1 gate15500(.O (g25836), .I1 (g25368), .I2 (g23856));
OR2X1 gate15501(.O (g27026), .I1 (g26828), .I2 (g17726));
OR2X1 gate15502(.O (g34254), .I1 (g34116), .I2 (g24301));
OR2X1 gate15503(.O (g30466), .I1 (g30174), .I2 (g21937));
OR2X1 gate15504(.O (g34809), .I1 (g33677), .I2 (g34738));
OR2X1 gate15505(.O (g34900), .I1 (g34860), .I2 (g21686));
OR2X1 gate15506(.O (g26733), .I1 (g10776), .I2 (g24447));
OR2X1 gate15507(.O (g34466), .I1 (g34337), .I2 (g18716));
OR2X1 gate15508(.O (g34808), .I1 (g34765), .I2 (g18599));
OR2X1 gate15509(.O (g32222), .I1 (g31141), .I2 (g29636));
OR3X1 gate15510(.O (g23771), .I1 (g21432), .I2 (g21416), .I3 (I22912));
OR2X1 gate15511(.O (g26874), .I1 (I25612), .I2 (I25613));
OR2X1 gate15512(.O (g34036), .I1 (g33722), .I2 (g18715));
OR2X1 gate15513(.O (g30560), .I1 (g30278), .I2 (g22131));
OR2X1 gate15514(.O (g34101), .I1 (g33693), .I2 (g33700));
OR2X1 gate15515(.O (g31916), .I1 (g31756), .I2 (g22002));
OR2X1 gate15516(.O (g34642), .I1 (g34482), .I2 (g18725));
OR2X1 gate15517(.O (g25749), .I1 (g25094), .I2 (g18800));
OR2X1 gate15518(.O (g25616), .I1 (g25096), .I2 (g18172));
OR2X1 gate15519(.O (g28649), .I1 (g27390), .I2 (g16597));
OR2X1 gate15520(.O (g33550), .I1 (g33342), .I2 (g18338));
OR2X1 gate15521(.O (g32347), .I1 (g29839), .I2 (g31273));
OR2X1 gate15522(.O (g33314), .I1 (g29663), .I2 (g32174));
OR2X1 gate15523(.O (g31287), .I1 (g29578), .I2 (g28292));
OR2X1 gate15524(.O (g15800), .I1 (g10821), .I2 (g13242));
OR2X1 gate15525(.O (g32253), .I1 (g24771), .I2 (g31207));
OR2X1 gate15526(.O (g25748), .I1 (g25078), .I2 (g18799));
OR2X1 gate15527(.O (g33287), .I1 (g32146), .I2 (g29586));
OR2X1 gate15528(.O (g34064), .I1 (g33919), .I2 (g33922));
OR2X1 gate15529(.O (g30733), .I1 (g13807), .I2 (g29773));
OR2X1 gate15530(.O (g31307), .I1 (g29596), .I2 (g28311));
OR2X1 gate15531(.O (g33076), .I1 (g32336), .I2 (g32446));
OR2X1 gate15532(.O (g34733), .I1 (g34678), .I2 (g18651));
OR2X1 gate15533(.O (g26892), .I1 (g26719), .I2 (g24198));
OR2X1 gate15534(.O (g25704), .I1 (g25173), .I2 (g21925));
OR2X1 gate15535(.O (g22447), .I1 (g21464), .I2 (g12761));
OR2X1 gate15536(.O (g33596), .I1 (g33341), .I2 (g18494));
OR2X1 gate15537(.O (g33054), .I1 (g31975), .I2 (g21975));
OR2X1 gate15538(.O (g32236), .I1 (g31152), .I2 (g29664));
OR2X1 gate15539(.O (g8790), .I1 (I12782), .I2 (I12783));
OR2X1 gate15540(.O (g32351), .I1 (g29851), .I2 (g31281));
OR2X1 gate15541(.O (g32372), .I1 (g29884), .I2 (g31314));
OR2X1 gate15542(.O (g34630), .I1 (g34560), .I2 (g15117));
OR2X1 gate15543(.O (g34693), .I1 (g34513), .I2 (g34310));
OR2X1 gate15544(.O (g24282), .I1 (g23407), .I2 (g18657));
OR2X1 gate15545(.O (g26914), .I1 (g25949), .I2 (g18227));
OR2X1 gate15546(.O (g29706), .I1 (g28198), .I2 (g27208));
OR2X1 gate15547(.O (g8461), .I1 (g301), .I2 (g534));
OR2X1 gate15548(.O (g31269), .I1 (g26024), .I2 (g29569));
OR2X1 gate15549(.O (g34166), .I1 (g33785), .I2 (g19752));
OR2X1 gate15550(.O (g34009), .I1 (g33863), .I2 (g18477));
OR2X1 gate15551(.O (g19336), .I1 (g17769), .I2 (g14831));
OR2X1 gate15552(.O (g26907), .I1 (g26513), .I2 (g24224));
OR2X1 gate15553(.O (g29256), .I1 (g28597), .I2 (g18533));
OR2X1 gate15554(.O (g31773), .I1 (g30044), .I2 (g30056));
OR4X1 gate15555(.O (I30399), .I1 (g29385), .I2 (g31376), .I3 (g30735), .I4 (g30825));
OR2X1 gate15556(.O (g31268), .I1 (g29552), .I2 (g28266));
OR2X1 gate15557(.O (g32264), .I1 (g31187), .I2 (g29711));
OR2X1 gate15558(.O (g34008), .I1 (g33849), .I2 (g18476));
OR2X1 gate15559(.O (g29280), .I1 (g28530), .I2 (g18742));
OR2X1 gate15560(.O (g33268), .I1 (g32116), .I2 (g29538));
OR2X1 gate15561(.O (g30476), .I1 (g30229), .I2 (g21947));
OR2X1 gate15562(.O (g30485), .I1 (g30166), .I2 (g21981));
OR2X1 gate15563(.O (g29300), .I1 (g28666), .I2 (g18796));
OR2X1 gate15564(.O (g31670), .I1 (g29937), .I2 (g28573));
OR2X1 gate15565(.O (g8904), .I1 (g1779), .I2 (g1798));
OR4X1 gate15566(.O (I31863), .I1 (g33506), .I2 (g33507), .I3 (g33508), .I4 (g33509));
OR2X1 gate15567(.O (g30555), .I1 (g30227), .I2 (g22126));
OR2X1 gate15568(.O (g30454), .I1 (g29909), .I2 (g21863));
OR2X1 gate15569(.O (g34454), .I1 (g34414), .I2 (g18667));
OR2X1 gate15570(.O (g25733), .I1 (g25108), .I2 (g18778));
OR3X1 gate15571(.O (g13091), .I1 (g329), .I2 (g319), .I3 (g10796));
OR2X1 gate15572(.O (g22591), .I1 (g18893), .I2 (g18909));
OR2X1 gate15573(.O (g27133), .I1 (g25788), .I2 (g24392));
OR2X1 gate15574(.O (g28719), .I1 (g27485), .I2 (g16703));
OR4X1 gate15575(.O (g28191), .I1 (g27217), .I2 (g27210), .I3 (g27186), .I4 (g27162));
OR2X1 gate15576(.O (g31930), .I1 (g31769), .I2 (g22094));
OR2X1 gate15577(.O (g32209), .I1 (g31122), .I2 (g29599));
OR2X1 gate15578(.O (g33993), .I1 (g33646), .I2 (g18413));
OR2X1 gate15579(.O (g25630), .I1 (g24532), .I2 (g18263));
OR2X1 gate15580(.O (g28718), .I1 (g27483), .I2 (g16702));
OR2X1 gate15581(.O (g25693), .I1 (g24627), .I2 (g18707));
OR2X1 gate15582(.O (g29231), .I1 (g28301), .I2 (g18229));
OR2X1 gate15583(.O (g33694), .I1 (g32402), .I2 (g33429));
OR2X1 gate15584(.O (g32208), .I1 (g31120), .I2 (g29584));
OR2X1 gate15585(.O (g33965), .I1 (g33805), .I2 (g18179));
OR4X1 gate15586(.O (I12783), .I1 (g4204), .I2 (g4207), .I3 (g4210), .I4 (g4180));
OR2X1 gate15587(.O (g25665), .I1 (g24708), .I2 (g21790));
OR2X1 gate15588(.O (g34239), .I1 (g32845), .I2 (g33957));
OR2X1 gate15589(.O (g34238), .I1 (g32780), .I2 (g33956));
OR2X1 gate15590(.O (g23345), .I1 (g19735), .I2 (g16203));
OR2X1 gate15591(.O (g26883), .I1 (g26670), .I2 (g24189));
OR4X1 gate15592(.O (I23162), .I1 (g19919), .I2 (g19968), .I3 (g20014), .I4 (g20841));
OR2X1 gate15593(.O (g33619), .I1 (g33359), .I2 (g18758));
OR2X1 gate15594(.O (g33557), .I1 (g33331), .I2 (g18363));
OR2X1 gate15595(.O (g29763), .I1 (g28217), .I2 (g22762));
OR2X1 gate15596(.O (g30382), .I1 (g30137), .I2 (g18498));
OR2X1 gate15597(.O (g30519), .I1 (g30264), .I2 (g22040));
OR2X1 gate15598(.O (g33618), .I1 (g33353), .I2 (g18757));
OR2X1 gate15599(.O (g28389), .I1 (g27206), .I2 (g15860));
OR2X1 gate15600(.O (g30176), .I1 (g23392), .I2 (g28531));
OR2X1 gate15601(.O (g28045), .I1 (g27378), .I2 (g18141));
OR2X1 gate15602(.O (g30092), .I1 (g28466), .I2 (g16699));
OR2X1 gate15603(.O (g31279), .I1 (g29571), .I2 (g29579));
OR2X1 gate15604(.O (g24249), .I1 (g22624), .I2 (g18294));
OR2X1 gate15605(.O (g33279), .I1 (g32140), .I2 (g29573));
OR2X1 gate15606(.O (g25712), .I1 (g25126), .I2 (g21963));
OR2X1 gate15607(.O (g28099), .I1 (g27992), .I2 (g22043));
OR2X1 gate15608(.O (g30518), .I1 (g30254), .I2 (g22039));
OR3X1 gate15609(.O (I22280), .I1 (g20271), .I2 (g20150), .I3 (g20134));
OR2X1 gate15610(.O (g28388), .I1 (g27204), .I2 (g15859));
OR2X1 gate15611(.O (g16430), .I1 (g182), .I2 (g13657));
OR2X1 gate15612(.O (g28701), .I1 (g27455), .I2 (g16669));
OR2X1 gate15613(.O (g24248), .I1 (g22710), .I2 (g18286));
OR2X1 gate15614(.O (g33278), .I1 (g32139), .I2 (g29572));
OR2X1 gate15615(.O (g12925), .I1 (g8928), .I2 (g10511));
OR2X1 gate15616(.O (g28777), .I1 (g27539), .I2 (g16807));
OR2X1 gate15617(.O (g28534), .I1 (g27292), .I2 (g26204));
OR2X1 gate15618(.O (g28098), .I1 (g27683), .I2 (g22016));
OR2X1 gate15619(.O (g32346), .I1 (g29838), .I2 (g31272));
OR2X1 gate15620(.O (g34637), .I1 (g34478), .I2 (g18694));
OR2X1 gate15621(.O (g24204), .I1 (g22990), .I2 (g18108));
OR2X1 gate15622(.O (g33286), .I1 (g32145), .I2 (g29585));
OR2X1 gate15623(.O (g31468), .I1 (g29641), .I2 (g29656));
OR2X1 gate15624(.O (g31306), .I1 (g29595), .I2 (g29610));
OR4X1 gate15625(.O (I31873), .I1 (g33524), .I2 (g33525), .I3 (g33526), .I4 (g33527));
OR2X1 gate15626(.O (g33039), .I1 (g32187), .I2 (g24312));
OR2X1 gate15627(.O (g29480), .I1 (g28115), .I2 (g22172));
OR2X1 gate15628(.O (g27742), .I1 (g17292), .I2 (g26673));
OR2X1 gate15629(.O (g22318), .I1 (g21394), .I2 (g17783));
OR2X1 gate15630(.O (g25594), .I1 (g24772), .I2 (g21708));
OR2X1 gate15631(.O (g33038), .I1 (g32184), .I2 (g24311));
OR2X1 gate15632(.O (g29287), .I1 (g28555), .I2 (g18760));
OR2X1 gate15633(.O (g29307), .I1 (g28706), .I2 (g18814));
OR2X1 gate15634(.O (g28140), .I1 (I26643), .I2 (I26644));
OR2X1 gate15635(.O (g26349), .I1 (g24630), .I2 (g13409));
OR2X1 gate15636(.O (g33601), .I1 (g33422), .I2 (g18508));
OR2X1 gate15637(.O (g25941), .I1 (g24416), .I2 (g22219));
OR3X1 gate15638(.O (g33187), .I1 (g32014), .I2 (I30740), .I3 (I30741));
OR2X1 gate15639(.O (g33975), .I1 (g33860), .I2 (g18346));
OR2X1 gate15640(.O (g27429), .I1 (g25969), .I2 (g24589));
OR2X1 gate15641(.O (g26906), .I1 (g26423), .I2 (g24223));
OR2X1 gate15642(.O (g25675), .I1 (g24769), .I2 (g21832));
OR2X1 gate15643(.O (g29243), .I1 (g28657), .I2 (g18358));
OR2X1 gate15644(.O (g26348), .I1 (g8466), .I2 (g24609));
OR2X1 gate15645(.O (g30501), .I1 (g29327), .I2 (g22018));
OR2X1 gate15646(.O (g28061), .I1 (g27287), .I2 (g21735));
OR2X1 gate15647(.O (g34729), .I1 (g34666), .I2 (g18270));
OR2X1 gate15648(.O (g32408), .I1 (g31541), .I2 (g30073));
OR2X1 gate15649(.O (g30439), .I1 (g29761), .I2 (g21848));
OR2X1 gate15650(.O (g34728), .I1 (g34661), .I2 (g18214));
OR2X1 gate15651(.O (g34439), .I1 (g34344), .I2 (g18181));
OR2X1 gate15652(.O (g29269), .I1 (g28249), .I2 (g18634));
OR2X1 gate15653(.O (g25637), .I1 (g24618), .I2 (g18307));
OR2X1 gate15654(.O (g24233), .I1 (g22590), .I2 (g18236));
OR2X1 gate15655(.O (g25935), .I1 (g24402), .I2 (g22208));
OR2X1 gate15656(.O (g30438), .I1 (g29890), .I2 (g21847));
OR2X1 gate15657(.O (g19525), .I1 (g7696), .I2 (g16811));
OR2X1 gate15658(.O (g19488), .I1 (g16965), .I2 (g14148));
OR2X1 gate15659(.O (g34438), .I1 (g34348), .I2 (g18150));
OR2X1 gate15660(.O (g29268), .I1 (g28343), .I2 (g18625));
OR4X1 gate15661(.O (I25613), .I1 (g25571), .I2 (g25572), .I3 (g25573), .I4 (g25574));
OR2X1 gate15662(.O (g31884), .I1 (g31290), .I2 (g21778));
OR2X1 gate15663(.O (g33791), .I1 (g33379), .I2 (g32430));
OR2X1 gate15664(.O (g30349), .I1 (g30051), .I2 (g18333));
OR2X1 gate15665(.O (g34349), .I1 (g26019), .I2 (g34104));
OR3X1 gate15666(.O (g8417), .I1 (g1056), .I2 (g1116), .I3 (I12583));
OR2X1 gate15667(.O (g30348), .I1 (g30083), .I2 (g18329));
OR2X1 gate15668(.O (g22645), .I1 (g18982), .I2 (g15633));
OR2X1 gate15669(.O (g34906), .I1 (g34857), .I2 (g21694));
OR2X1 gate15670(.O (g29734), .I1 (g28201), .I2 (g15872));
OR2X1 gate15671(.O (g30304), .I1 (g28255), .I2 (g27259));
OR2X1 gate15672(.O (g33015), .I1 (g32343), .I2 (g18507));
OR2X1 gate15673(.O (g34622), .I1 (g34520), .I2 (g18584));
OR2X1 gate15674(.O (g25729), .I1 (g25091), .I2 (g22012));
OR4X1 gate15675(.O (g26636), .I1 (g24897), .I2 (g24884), .I3 (g24858), .I4 (g24846));
OR2X1 gate15676(.O (g28629), .I1 (g27371), .I2 (g16532));
OR2X1 gate15677(.O (g25577), .I1 (g24143), .I2 (g24144));
OR3X1 gate15678(.O (g28220), .I1 (g23495), .I2 (I26741), .I3 (I26742));
OR2X1 gate15679(.O (g25728), .I1 (g25076), .I2 (g22011));
OR2X1 gate15680(.O (g28628), .I1 (g27370), .I2 (g16531));
OR2X1 gate15681(.O (g33556), .I1 (g33329), .I2 (g18362));
OR2X1 gate15682(.O (g24212), .I1 (g23280), .I2 (g18155));
OR2X1 gate15683(.O (g26963), .I1 (g26306), .I2 (g24308));
OR2X1 gate15684(.O (g33580), .I1 (g33330), .I2 (g18442));
OR2X1 gate15685(.O (g29487), .I1 (g25815), .I2 (g28133));
OR2X1 gate15686(.O (g23795), .I1 (g20203), .I2 (g16884));
OR2X1 gate15687(.O (g28071), .I1 (g27085), .I2 (g21873));
OR2X1 gate15688(.O (g29502), .I1 (g28139), .I2 (g25871));
OR2X1 gate15689(.O (g27533), .I1 (g26078), .I2 (g24659));
OR4X1 gate15690(.O (I29351), .I1 (g29328), .I2 (g29323), .I3 (g29316), .I4 (g30316));
OR2X1 gate15691(.O (g28591), .I1 (g27332), .I2 (g26286));
OR2X1 gate15692(.O (g25906), .I1 (g25559), .I2 (g24014));
OR2X1 gate15693(.O (g28776), .I1 (g27538), .I2 (g13974));
OR2X1 gate15694(.O (g30415), .I1 (g29843), .I2 (g21799));
OR2X1 gate15695(.O (g30333), .I1 (g29834), .I2 (g21699));
OR2X1 gate15696(.O (g34636), .I1 (g34476), .I2 (g18693));
OR2X1 gate15697(.O (g22547), .I1 (g16855), .I2 (g20215));
OR2X1 gate15698(.O (g29279), .I1 (g28442), .I2 (g18741));
OR2X1 gate15699(.O (g31922), .I1 (g31525), .I2 (g22047));
OR2X1 gate15700(.O (g32982), .I1 (g31948), .I2 (g18208));
OR2X1 gate15701(.O (g33321), .I1 (g29712), .I2 (g32182));
OR2X1 gate15702(.O (g25622), .I1 (g24546), .I2 (g18217));
OR2X1 gate15703(.O (g29278), .I1 (g28626), .I2 (g18740));
OR2X1 gate15704(.O (g19267), .I1 (g17752), .I2 (g17768));
OR2X1 gate15705(.O (g22226), .I1 (g21333), .I2 (g17655));
OR2X1 gate15706(.O (g24433), .I1 (g10878), .I2 (g22400));
OR2X1 gate15707(.O (g20148), .I1 (g16128), .I2 (g13393));
OR2X1 gate15708(.O (g29286), .I1 (g28542), .I2 (g18759));
OR2X1 gate15709(.O (g27232), .I1 (g25874), .I2 (g24450));
OR2X1 gate15710(.O (g7404), .I1 (g933), .I2 (g939));
OR2X1 gate15711(.O (g29306), .I1 (g28689), .I2 (g18813));
OR4X1 gate15712(.O (g28172), .I1 (g27469), .I2 (g27440), .I3 (g27416), .I4 (g27395));
OR2X1 gate15713(.O (g33685), .I1 (g32396), .I2 (g33423));
OR2X1 gate15714(.O (g7764), .I1 (g2999), .I2 (g2932));
OR3X1 gate15715(.O (g33953), .I1 (g33487), .I2 (I31848), .I3 (I31849));
OR2X1 gate15716(.O (g24343), .I1 (g23724), .I2 (g18773));
OR2X1 gate15717(.O (g26921), .I1 (g25955), .I2 (g18285));
OR2X1 gate15718(.O (g25653), .I1 (g24664), .I2 (g18602));
OR2X1 gate15719(.O (g32390), .I1 (g31501), .I2 (g29979));
OR2X1 gate15720(.O (g27261), .I1 (g24544), .I2 (g25996));
OR2X1 gate15721(.O (g30484), .I1 (g30154), .I2 (g21980));
OR2X1 gate15722(.O (g30554), .I1 (g30216), .I2 (g22125));
OR2X1 gate15723(.O (g22490), .I1 (g21513), .I2 (g12795));
OR3X1 gate15724(.O (g13820), .I1 (g11184), .I2 (g9187), .I3 (g12527));
OR2X1 gate15725(.O (g26813), .I1 (g24940), .I2 (g24949));
OR4X1 gate15726(.O (g15727), .I1 (g13383), .I2 (g13345), .I3 (g13333), .I4 (g11010));
OR2X1 gate15727(.O (g25636), .I1 (g24507), .I2 (g18305));
OR2X1 gate15728(.O (g30609), .I1 (g13633), .I2 (g29742));
OR2X1 gate15729(.O (g34609), .I1 (g34503), .I2 (g18563));
OR2X1 gate15730(.O (g28420), .I1 (g27222), .I2 (g13290));
OR2X1 gate15731(.O (g30608), .I1 (g13604), .I2 (g29736));
OR2X1 gate15732(.O (g28319), .I1 (g27115), .I2 (g15807));
OR2X1 gate15733(.O (g30115), .I1 (g28489), .I2 (g11449));
OR2X1 gate15734(.O (g29143), .I1 (g27650), .I2 (g17146));
OR2X1 gate15735(.O (g34608), .I1 (g34568), .I2 (g15082));
OR4X1 gate15736(.O (g17490), .I1 (g14364), .I2 (g14337), .I3 (g11958), .I4 (I18421));
OR2X1 gate15737(.O (g26805), .I1 (g10776), .I2 (g24478));
OR2X1 gate15738(.O (g31762), .I1 (g30011), .I2 (g30030));
OR2X1 gate15739(.O (g23358), .I1 (g19746), .I2 (g16212));
OR4X1 gate15740(.O (I30760), .I1 (g31778), .I2 (g32295), .I3 (g32046), .I4 (g32050));
OR2X1 gate15741(.O (g31964), .I1 (g31654), .I2 (g14544));
OR2X1 gate15742(.O (g33964), .I1 (g33817), .I2 (g18146));
OR2X1 gate15743(.O (g25664), .I1 (g24681), .I2 (g21789));
OR2X1 gate15744(.O (g28059), .I1 (g27042), .I2 (g18276));
OR2X1 gate15745(.O (g29791), .I1 (g28233), .I2 (g22859));
OR2X1 gate15746(.O (g16021), .I1 (g13047), .I2 (g10706));
OR2X1 gate15747(.O (g26934), .I1 (g26845), .I2 (g18556));
OR2X1 gate15748(.O (g28058), .I1 (g27235), .I2 (g18268));
OR2X1 gate15749(.O (g29168), .I1 (g27658), .I2 (g26613));
OR2X1 gate15750(.O (g33587), .I1 (g33363), .I2 (g18463));
OR2X1 gate15751(.O (g24896), .I1 (g22863), .I2 (g19684));
OR2X1 gate15752(.O (g34799), .I1 (g34751), .I2 (g18578));
OR2X1 gate15753(.O (g25585), .I1 (g21674), .I2 (g24155));
OR2X1 gate15754(.O (g25576), .I1 (g24141), .I2 (g24142));
OR2X1 gate15755(.O (g29479), .I1 (g28113), .I2 (g28116));
OR2X1 gate15756(.O (g34798), .I1 (g34754), .I2 (g18575));
OR2X1 gate15757(.O (g31909), .I1 (g31750), .I2 (g21956));
OR2X1 gate15758(.O (g28044), .I1 (g27256), .I2 (g18130));
OR2X1 gate15759(.O (g33543), .I1 (g33106), .I2 (g18281));
OR2X1 gate15760(.O (g19595), .I1 (g17149), .I2 (g14218));
OR2X1 gate15761(.O (g29478), .I1 (g28111), .I2 (g22160));
OR2X1 gate15762(.O (g19467), .I1 (g16896), .I2 (g14097));
OR2X1 gate15763(.O (g25609), .I1 (g24915), .I2 (g18126));
OR2X1 gate15764(.O (g34805), .I1 (g34748), .I2 (g18594));
OR2X1 gate15765(.O (g31908), .I1 (g31519), .I2 (g21955));
OR2X1 gate15766(.O (g33000), .I1 (g32270), .I2 (g18403));
OR2X1 gate15767(.O (g29486), .I1 (g28537), .I2 (g27595));
OR2X1 gate15768(.O (g32252), .I1 (g31183), .I2 (g31206));
OR2X1 gate15769(.O (g25608), .I1 (g24643), .I2 (g18120));
OR2X1 gate15770(.O (g33569), .I1 (g33415), .I2 (g18402));
OR2X1 gate15771(.O (g30732), .I1 (g13778), .I2 (g29762));
OR2X1 gate15772(.O (g27271), .I1 (g24547), .I2 (g26053));
OR3X1 gate15773(.O (I18495), .I1 (g14539), .I2 (g14515), .I3 (g14449));
OR2X1 gate15774(.O (g34732), .I1 (g34686), .I2 (g18593));
OR2X1 gate15775(.O (g26329), .I1 (g8526), .I2 (g24609));
OR2X1 gate15776(.O (g33568), .I1 (g33409), .I2 (g18395));
OR2X1 gate15777(.O (g25745), .I1 (g25150), .I2 (g22060));
OR2X1 gate15778(.O (g29223), .I1 (g28341), .I2 (g18131));
OR2X1 gate15779(.O (g26328), .I1 (g1183), .I2 (g24591));
OR2X1 gate15780(.O (g28562), .I1 (g27313), .I2 (g26251));
OR2X1 gate15781(.O (g14844), .I1 (g10776), .I2 (g8703));
OR2X1 gate15782(.O (g34761), .I1 (g34679), .I2 (g34506));
OR2X1 gate15783(.O (g28699), .I1 (g27452), .I2 (g16667));
OR4X1 gate15784(.O (g27031), .I1 (g26213), .I2 (g26190), .I3 (g26166), .I4 (g26148));
OR2X1 gate15785(.O (g33123), .I1 (g31962), .I2 (g30577));
OR4X1 gate15786(.O (I30755), .I1 (g30564), .I2 (g32303), .I3 (g32049), .I4 (g32055));
OR2X1 gate15787(.O (g28698), .I1 (g27451), .I2 (g16666));
OR2X1 gate15788(.O (g31751), .I1 (g29975), .I2 (g29990));
OR2X1 gate15789(.O (g31772), .I1 (g30035), .I2 (g28654));
OR2X1 gate15790(.O (g30400), .I1 (g29766), .I2 (g21759));
OR2X1 gate15791(.O (g33974), .I1 (g33846), .I2 (g18345));
OR2X1 gate15792(.O (g30214), .I1 (g23424), .I2 (g28572));
OR2X1 gate15793(.O (g34013), .I1 (g33901), .I2 (g18488));
OR4X1 gate15794(.O (g25805), .I1 (g25453), .I2 (g25414), .I3 (g25374), .I4 (g25331));
OR2X1 gate15795(.O (g25674), .I1 (g24755), .I2 (g21831));
OR2X1 gate15796(.O (g31293), .I1 (g29582), .I2 (g28299));
OR2X1 gate15797(.O (g33293), .I1 (g32151), .I2 (g29602));
OR2X1 gate15798(.O (g30539), .I1 (g30267), .I2 (g22085));
OR2X1 gate15799(.O (g34207), .I1 (g33835), .I2 (g33304));
OR2X1 gate15800(.O (g22659), .I1 (g19062), .I2 (g15673));
OR2X1 gate15801(.O (g22625), .I1 (g18910), .I2 (g18933));
OR2X1 gate15802(.O (g25732), .I1 (g25201), .I2 (g22017));
OR2X1 gate15803(.O (g34005), .I1 (g33883), .I2 (g18454));
OR2X1 gate15804(.O (g28632), .I1 (g27373), .I2 (g16535));
OR2X1 gate15805(.O (g33265), .I1 (g32113), .I2 (g29530));
OR2X1 gate15806(.O (g30538), .I1 (g30256), .I2 (g22084));
OR2X1 gate15807(.O (g29373), .I1 (g13832), .I2 (g28453));
OR4X1 gate15808(.O (I30262), .I1 (g31672), .I2 (g31710), .I3 (g31021), .I4 (g30937));
OR2X1 gate15809(.O (g33992), .I1 (g33900), .I2 (g18408));
OR2X1 gate15810(.O (g25761), .I1 (g25152), .I2 (g18812));
OR2X1 gate15811(.O (g28661), .I1 (g27406), .I2 (g16611));
OR2X1 gate15812(.O (g28403), .I1 (g27214), .I2 (g13282));
OR2X1 gate15813(.O (g22644), .I1 (g18981), .I2 (g15632));
OR4X1 gate15814(.O (I12782), .I1 (g4188), .I2 (g4194), .I3 (g4197), .I4 (g4200));
OR2X1 gate15815(.O (g33579), .I1 (g33357), .I2 (g18437));
OR2X1 gate15816(.O (g14044), .I1 (g10776), .I2 (g8703));
OR2X1 gate15817(.O (g28715), .I1 (g27480), .I2 (g16700));
OR4X1 gate15818(.O (I30718), .I1 (g32348), .I2 (g32356), .I3 (g32097), .I4 (g32020));
OR2X1 gate15819(.O (g33578), .I1 (g33410), .I2 (g18433));
OR2X1 gate15820(.O (g31014), .I1 (g29367), .I2 (g28160));
OR2X1 gate15821(.O (g27225), .I1 (g2975), .I2 (g26364));
OR2X1 gate15822(.O (g33014), .I1 (g32305), .I2 (g18499));
OR2X1 gate15823(.O (g23770), .I1 (g20188), .I2 (g16868));
OR2X1 gate15824(.O (g26882), .I1 (g26650), .I2 (g24188));
OR2X1 gate15825(.O (g28551), .I1 (g27305), .I2 (g26234));
OR2X1 gate15826(.O (g31007), .I1 (g29364), .I2 (g28159));
OR2X1 gate15827(.O (g27258), .I1 (g25905), .I2 (g15749));
OR2X1 gate15828(.O (g34100), .I1 (g33690), .I2 (g33697));
OR2X1 gate15829(.O (g33586), .I1 (g33416), .I2 (g18459));
OR2X1 gate15830(.O (g33007), .I1 (g32331), .I2 (g18455));
OR2X1 gate15831(.O (g25539), .I1 (g23531), .I2 (g20628));
OR2X1 gate15832(.O (g13662), .I1 (g10896), .I2 (g10917));
OR2X1 gate15833(.O (g34235), .I1 (g32585), .I2 (g33953));
OR2X1 gate15834(.O (g27244), .I1 (g24652), .I2 (g25995));
OR2X1 gate15835(.O (g28490), .I1 (g27262), .I2 (g16185));
OR2X1 gate15836(.O (g33116), .I1 (g32403), .I2 (g32411));
OR2X1 gate15837(.O (g33615), .I1 (g33113), .I2 (g21871));
OR2X1 gate15838(.O (g23262), .I1 (g19661), .I2 (g16126));
OR2X1 gate15839(.O (g21899), .I1 (g20162), .I2 (g15113));
OR2X1 gate15840(.O (g30515), .I1 (g30223), .I2 (g22036));
OR2X1 gate15841(.O (g30414), .I1 (g30002), .I2 (g21794));
OR2X1 gate15842(.O (g28385), .I1 (g27201), .I2 (g15857));
OR2X1 gate15843(.O (g33041), .I1 (g32189), .I2 (g24323));
OR2X1 gate15844(.O (g28297), .I1 (g27096), .I2 (g15785));
OR2X1 gate15845(.O (g21898), .I1 (g20152), .I2 (g15112));
OR2X1 gate15846(.O (g34882), .I1 (g34876), .I2 (g18659));
OR2X1 gate15847(.O (g28103), .I1 (g27696), .I2 (g22097));
OR2X1 gate15848(.O (g24245), .I1 (g22849), .I2 (g18256));
OR2X1 gate15849(.O (g33275), .I1 (g32127), .I2 (g29564));
OR2X1 gate15850(.O (g28095), .I1 (g27674), .I2 (g21970));
OR2X1 gate15851(.O (g30407), .I1 (g29794), .I2 (g21766));
OR2X1 gate15852(.O (g34407), .I1 (g34185), .I2 (g25124));
OR2X1 gate15853(.O (g27970), .I1 (g26514), .I2 (g25050));
OR2X1 gate15854(.O (g31465), .I1 (g26156), .I2 (g29647));
OR2X1 gate15855(.O (g26759), .I1 (g24468), .I2 (g7511));
OR2X1 gate15856(.O (g26725), .I1 (g24457), .I2 (g10719));
OR2X1 gate15857(.O (g28671), .I1 (g27413), .I2 (g16619));
OR2X1 gate15858(.O (g33983), .I1 (g33877), .I2 (g18373));
OR2X1 gate15859(.O (g22707), .I1 (g20559), .I2 (g17156));
OR2X1 gate15860(.O (g33035), .I1 (g32019), .I2 (g21872));
OR2X1 gate15861(.O (g27886), .I1 (g14438), .I2 (g26759));
OR2X1 gate15862(.O (g25683), .I1 (g24669), .I2 (g18641));
OR2X1 gate15863(.O (g29242), .I1 (g28674), .I2 (g18354));
OR2X1 gate15864(.O (g26082), .I1 (g2898), .I2 (g24561));
OR2X1 gate15865(.O (g11380), .I1 (g8583), .I2 (g8530));
OR2X1 gate15866(.O (g30441), .I1 (g29787), .I2 (g21850));
OR2X1 gate15867(.O (g34441), .I1 (g34381), .I2 (g18540));
OR2X1 gate15868(.O (g24232), .I1 (g22686), .I2 (g18228));
OR2X1 gate15869(.O (g34206), .I1 (g33834), .I2 (g33836));
OR2X1 gate15870(.O (g26940), .I1 (g25908), .I2 (g21886));
OR4X1 gate15871(.O (I25612), .I1 (g25567), .I2 (g25568), .I3 (g25569), .I4 (g25570));
OR2X1 gate15872(.O (g34725), .I1 (g34700), .I2 (g18183));
OR2X1 gate15873(.O (g24261), .I1 (g22862), .I2 (g18314));
OR2X1 gate15874(.O (g29230), .I1 (g28107), .I2 (g18202));
OR2X1 gate15875(.O (g27458), .I1 (g24590), .I2 (g25989));
OR2X1 gate15876(.O (g29293), .I1 (g28570), .I2 (g18777));
OR2X1 gate15877(.O (g30114), .I1 (g28488), .I2 (g16761));
OR2X1 gate15878(.O (g30435), .I1 (g30025), .I2 (g21840));
OR2X1 gate15879(.O (g29265), .I1 (g28318), .I2 (g18620));
OR2X1 gate15880(.O (g28546), .I1 (g27302), .I2 (g26231));
OR2X1 gate15881(.O (g28089), .I1 (g27269), .I2 (g18731));
OR2X1 gate15882(.O (g23251), .I1 (g19637), .I2 (g16098));
OR2X1 gate15883(.O (g28211), .I1 (g27029), .I2 (g27034));
OR2X1 gate15884(.O (g34107), .I1 (g33710), .I2 (g33121));
OR2X1 gate15885(.O (g19555), .I1 (g15672), .I2 (g13030));
OR2X1 gate15886(.O (g28088), .I1 (g27264), .I2 (g18729));
OR2X1 gate15887(.O (g30345), .I1 (g29644), .I2 (g18302));
OR2X1 gate15888(.O (g30399), .I1 (g29757), .I2 (g21758));
OR2X1 gate15889(.O (g34849), .I1 (g34842), .I2 (g18154));
OR2X1 gate15890(.O (g34399), .I1 (g34178), .I2 (g25067));
OR2X1 gate15891(.O (g25584), .I1 (g21670), .I2 (g24154));
OR2X1 gate15892(.O (g28497), .I1 (g27267), .I2 (g16199));
OR2X1 gate15893(.O (g33006), .I1 (g32291), .I2 (g18447));
OR2X1 gate15894(.O (g30398), .I1 (g29749), .I2 (g21757));
OR2X1 gate15895(.O (g26962), .I1 (g26295), .I2 (g24307));
OR2X1 gate15896(.O (g26361), .I1 (g24674), .I2 (g22991));
OR2X1 gate15897(.O (g23997), .I1 (g20602), .I2 (g17191));
OR2X1 gate15898(.O (g30141), .I1 (g28499), .I2 (g16844));
OR2X1 gate15899(.O (g34804), .I1 (g34740), .I2 (g18591));
OR2X1 gate15900(.O (g28700), .I1 (g27454), .I2 (g16668));
OR2X1 gate15901(.O (g25759), .I1 (g25166), .I2 (g22106));
OR2X1 gate15902(.O (g28659), .I1 (g27404), .I2 (g16610));
OR2X1 gate15903(.O (g25725), .I1 (g25127), .I2 (g22008));
OR2X1 gate15904(.O (g28625), .I1 (g27363), .I2 (g26324));
OR2X1 gate15905(.O (g14888), .I1 (g10776), .I2 (g8703));
OR2X1 gate15906(.O (g32357), .I1 (g29865), .I2 (g31296));
OR2X1 gate15907(.O (g27159), .I1 (g25814), .I2 (g12953));
OR2X1 gate15908(.O (g27532), .I1 (g16176), .I2 (g26084));
OR2X1 gate15909(.O (g25758), .I1 (g25151), .I2 (g22105));
OR2X1 gate15910(.O (g34263), .I1 (g34078), .I2 (g18699));
OR2X1 gate15911(.O (g34332), .I1 (g34071), .I2 (g33723));
OR2X1 gate15912(.O (g33703), .I1 (g32410), .I2 (g33434));
OR2X1 gate15913(.O (g28296), .I1 (g27095), .I2 (g15784));
OR2X1 gate15914(.O (g31253), .I1 (g25980), .I2 (g29533));
OR2X1 gate15915(.O (g27561), .I1 (g26100), .I2 (g24702));
OR2X1 gate15916(.O (g33253), .I1 (g32103), .I2 (g29511));
OR2X1 gate15917(.O (g25744), .I1 (g25129), .I2 (g22059));
OR2X1 gate15918(.O (g28644), .I1 (g27387), .I2 (g16593));
OR2X1 gate15919(.O (g30406), .I1 (g29783), .I2 (g21765));
OR2X1 gate15920(.O (g24432), .I1 (g23900), .I2 (g21361));
OR2X1 gate15921(.O (g30361), .I1 (g30109), .I2 (g18391));
OR2X1 gate15922(.O (g34406), .I1 (g34184), .I2 (g25123));
OR2X1 gate15923(.O (g24271), .I1 (g23451), .I2 (g18628));
OR2X1 gate15924(.O (g33600), .I1 (g33418), .I2 (g18501));
OR2X1 gate15925(.O (g25940), .I1 (g24415), .I2 (g22218));
OR2X1 gate15926(.O (g31781), .I1 (g30058), .I2 (g30069));
OR3X1 gate15927(.O (g23162), .I1 (g20184), .I2 (g20170), .I3 (I22267));
OR2X1 gate15928(.O (g33236), .I1 (g32044), .I2 (g32045));
OR2X1 gate15929(.O (g30500), .I1 (g29326), .I2 (g21996));
OR2X1 gate15930(.O (g29275), .I1 (g28165), .I2 (g21868));
OR2X1 gate15931(.O (g28060), .I1 (g27616), .I2 (g18532));
OR3X1 gate15932(.O (g33952), .I1 (g33478), .I2 (I31843), .I3 (I31844));
OR2X1 gate15933(.O (g24342), .I1 (g23691), .I2 (g18772));
OR2X1 gate15934(.O (g25652), .I1 (g24777), .I2 (g21747));
OR2X1 gate15935(.O (g26947), .I1 (g26394), .I2 (g24285));
OR2X1 gate15936(.O (g8905), .I1 (g2204), .I2 (g2223));
OR2X1 gate15937(.O (g29237), .I1 (g28185), .I2 (g18289));
OR2X1 gate15938(.O (g28527), .I1 (g27286), .I2 (g26182));
OR2X1 gate15939(.O (g33063), .I1 (g31988), .I2 (g22066));
OR2X1 gate15940(.O (g34004), .I1 (g33879), .I2 (g18453));
OR2X1 gate15941(.O (g26951), .I1 (g26390), .I2 (g24289));
OR2X1 gate15942(.O (g26972), .I1 (g26780), .I2 (g25229));
OR2X1 gate15943(.O (g31873), .I1 (g31270), .I2 (g21728));
OR2X1 gate15944(.O (g19501), .I1 (g16986), .I2 (g14168));
OR2X1 gate15945(.O (g34613), .I1 (g34515), .I2 (g18567));
OR2X1 gate15946(.O (g32249), .I1 (g31169), .I2 (g29687));
OR2X1 gate15947(.O (g30605), .I1 (g29529), .I2 (g29520));
OR2X1 gate15948(.O (g27289), .I1 (g25925), .I2 (g25927));
OR2X1 gate15949(.O (g34273), .I1 (g27765), .I2 (g34203));
OR2X1 gate15950(.O (g34605), .I1 (g34566), .I2 (g15077));
OR2X1 gate15951(.O (g18879), .I1 (g17365), .I2 (g14423));
OR2X1 gate15952(.O (g28581), .I1 (g27329), .I2 (g26276));
OR2X1 gate15953(.O (g27224), .I1 (g25870), .I2 (g15678));
OR2X1 gate15954(.O (g30463), .I1 (g30140), .I2 (g21934));
OR2X1 gate15955(.O (g27571), .I1 (g26127), .I2 (g24723));
OR2X1 gate15956(.O (g28707), .I1 (g27461), .I2 (g16673));
OR2X1 gate15957(.O (g34463), .I1 (g34338), .I2 (g18686));
OR2X1 gate15958(.O (g23825), .I1 (g20705), .I2 (g20781));
OR2X1 gate15959(.O (g30371), .I1 (g30099), .I2 (g18445));
OR2X1 gate15960(.O (g28818), .I1 (g27549), .I2 (g13998));
OR2X1 gate15961(.O (g34033), .I1 (g33821), .I2 (g18708));
OR2X1 gate15962(.O (g34234), .I1 (g32520), .I2 (g33952));
OR2X1 gate15963(.O (g28055), .I1 (g27560), .I2 (g18190));
OR2X1 gate15964(.O (g33542), .I1 (g33102), .I2 (g18265));
OR2X1 gate15965(.O (g33021), .I1 (g32302), .I2 (g21749));
OR2X1 gate15966(.O (g24259), .I1 (g23008), .I2 (g18312));
OR2X1 gate15967(.O (g28070), .I1 (g27050), .I2 (g21867));
OR2X1 gate15968(.O (g31913), .I1 (g31485), .I2 (g21999));
OR2X1 gate15969(.O (g18994), .I1 (g16303), .I2 (g13632));
OR2X1 gate15970(.O (g24471), .I1 (g10999), .I2 (g22450));
OR2X1 gate15971(.O (g34795), .I1 (g34753), .I2 (g18572));
OR2X1 gate15972(.O (g25613), .I1 (g25181), .I2 (g18140));
OR2X1 gate15973(.O (g24258), .I1 (g22851), .I2 (g18311));
OR2X1 gate15974(.O (g33614), .I1 (g33249), .I2 (g18650));
OR4X1 gate15975(.O (g17511), .I1 (g14396), .I2 (g14365), .I3 (g11976), .I4 (I18452));
OR2X1 gate15976(.O (g32999), .I1 (g32337), .I2 (g18401));
OR2X1 gate15977(.O (g33607), .I1 (g33091), .I2 (g18526));
OR2X1 gate15978(.O (g31905), .I1 (g31746), .I2 (g21952));
OR2X1 gate15979(.O (g31320), .I1 (g26125), .I2 (g29632));
OR2X1 gate15980(.O (g30514), .I1 (g30211), .I2 (g22035));
OR2X1 gate15981(.O (g32380), .I1 (g29907), .I2 (g31467));
OR2X1 gate15982(.O (g31274), .I1 (g29565), .I2 (g28280));
OR2X1 gate15983(.O (g25605), .I1 (g24743), .I2 (g18116));
OR2X1 gate15984(.O (g29222), .I1 (g28252), .I2 (g18105));
OR2X1 gate15985(.O (g24244), .I1 (g23349), .I2 (g18255));
OR2X1 gate15986(.O (g33274), .I1 (g32126), .I2 (g29563));
OR2X1 gate15987(.O (g30507), .I1 (g30190), .I2 (g22028));
OR2X1 gate15988(.O (g32998), .I1 (g32300), .I2 (g18393));
OR2X1 gate15989(.O (g28094), .I1 (g27673), .I2 (g21959));
OR2X1 gate15990(.O (g28067), .I1 (g27309), .I2 (g21827));
OR2X1 gate15991(.O (g33593), .I1 (g33417), .I2 (g18482));
OR2X1 gate15992(.O (g26789), .I1 (g10776), .I2 (g24471));
OR2X1 gate15993(.O (g32233), .I1 (g31150), .I2 (g29661));
OR2X1 gate15994(.O (g12954), .I1 (g12186), .I2 (g9906));
OR2X1 gate15995(.O (g23319), .I1 (g19717), .I2 (g16193));
OR2X1 gate15996(.O (g30421), .I1 (g29784), .I2 (g21805));
OR2X1 gate15997(.O (g33565), .I1 (g33338), .I2 (g18389));
OR2X1 gate15998(.O (g34421), .I1 (g27686), .I2 (g34198));
OR2X1 gate15999(.O (g26359), .I1 (g24651), .I2 (g22939));
OR2X1 gate16000(.O (g28735), .I1 (g27510), .I2 (g16737));
OR2X1 gate16001(.O (g23318), .I1 (g19716), .I2 (g16192));
OR2X1 gate16002(.O (g30163), .I1 (g23381), .I2 (g28523));
OR2X1 gate16003(.O (g33034), .I1 (g32340), .I2 (g21844));
OR2X1 gate16004(.O (g26920), .I1 (g25865), .I2 (g18283));
OR2X1 gate16005(.O (g34012), .I1 (g33886), .I2 (g18480));
OR2X1 gate16006(.O (g29253), .I1 (g28697), .I2 (g18490));
OR2X1 gate16007(.O (g24879), .I1 (g21465), .I2 (g24009));
OR2X1 gate16008(.O (g33292), .I1 (g32150), .I2 (g29601));
OR2X1 gate16009(.O (g26946), .I1 (g26389), .I2 (g24284));
OR2X1 gate16010(.O (g30541), .I1 (g30281), .I2 (g22087));
OR2X1 gate16011(.O (g30473), .I1 (g30196), .I2 (g21944));
OR2X1 gate16012(.O (g24337), .I1 (g23540), .I2 (g18754));
OR2X1 gate16013(.O (g27489), .I1 (g24608), .I2 (g26022));
OR2X1 gate16014(.O (g29236), .I1 (g28313), .I2 (g18287));
OR2X1 gate16015(.O (g28526), .I1 (g27285), .I2 (g26178));
OR2X1 gate16016(.O (g26344), .I1 (g2927), .I2 (g25010));
OR2X1 gate16017(.O (g27016), .I1 (g26821), .I2 (g14585));
OR2X1 gate16018(.O (g30359), .I1 (g30075), .I2 (g18385));
OR2X1 gate16019(.O (g34724), .I1 (g34702), .I2 (g18152));
OR2X1 gate16020(.O (g28402), .I1 (g27213), .I2 (g15873));
OR2X1 gate16021(.O (g30535), .I1 (g30225), .I2 (g22081));
OR2X1 gate16022(.O (g30434), .I1 (g30024), .I2 (g21818));
OR2X1 gate16023(.O (g19576), .I1 (g17138), .I2 (g14202));
OR2X1 gate16024(.O (g30358), .I1 (g30108), .I2 (g18381));
OR2X1 gate16025(.O (g34535), .I1 (g34309), .I2 (g34073));
OR2X1 gate16026(.O (g29264), .I1 (g28248), .I2 (g18618));
OR2X1 gate16027(.O (g29790), .I1 (g25975), .I2 (g28242));
OR2X1 gate16028(.O (g16928), .I1 (g13525), .I2 (g11127));
OR2X1 gate16029(.O (g27544), .I1 (g26087), .I2 (g24671));
OR3X1 gate16030(.O (g33164), .I1 (g32203), .I2 (I30727), .I3 (I30728));
OR2X1 gate16031(.O (g17268), .I1 (g9220), .I2 (g14387));
OR2X1 gate16032(.O (g24919), .I1 (g21606), .I2 (g22143));
OR2X1 gate16033(.O (g30344), .I1 (g29630), .I2 (g18298));
OR2X1 gate16034(.O (g31891), .I1 (g31305), .I2 (g21824));
OR2X1 gate16035(.O (g28077), .I1 (g27120), .I2 (g21879));
OR2X1 gate16036(.O (g33891), .I1 (g33264), .I2 (g33269));
OR2X1 gate16037(.O (g31474), .I1 (g29668), .I2 (g13583));
OR2X1 gate16038(.O (g33575), .I1 (g33086), .I2 (g18420));
OR2X1 gate16039(.O (g24444), .I1 (g10890), .I2 (g22400));
OR2X1 gate16040(.O (g30291), .I1 (g28672), .I2 (g27685));
OR2X1 gate16041(.O (g25789), .I1 (g25285), .I2 (g14543));
OR2X1 gate16042(.O (g32387), .I1 (g31489), .I2 (g29952));
OR2X1 gate16043(.O (g25724), .I1 (g25043), .I2 (g22007));
OR2X1 gate16044(.O (g28688), .I1 (g27435), .I2 (g16639));
OR2X1 gate16045(.O (g33537), .I1 (g33244), .I2 (g21716));
OR2X1 gate16046(.O (g22487), .I1 (g21512), .I2 (g12794));
OR2X1 gate16047(.O (g28102), .I1 (g27995), .I2 (g22089));
OR2X1 gate16048(.O (g33283), .I1 (g31995), .I2 (g30318));
OR2X1 gate16049(.O (g27383), .I1 (g24569), .I2 (g25961));
OR2X1 gate16050(.O (g33606), .I1 (g33369), .I2 (g18522));
OR2X1 gate16051(.O (g31303), .I1 (g29592), .I2 (g29606));
OR2X1 gate16052(.O (g33303), .I1 (g32159), .I2 (g29638));
OR2X1 gate16053(.O (g34029), .I1 (g33798), .I2 (g18703));
OR2X1 gate16054(.O (g26927), .I1 (g26711), .I2 (g18539));
OR2X1 gate16055(.O (g30506), .I1 (g30179), .I2 (g22027));
OR2X1 gate16056(.O (g28066), .I1 (g27553), .I2 (g21819));
OR2X1 gate16057(.O (g21895), .I1 (g20135), .I2 (g15108));
OR2X1 gate16058(.O (g34028), .I1 (g33720), .I2 (g18684));
OR2X1 gate16059(.O (g32368), .I1 (g29881), .I2 (g31310));
OR2X1 gate16060(.O (g33982), .I1 (g33865), .I2 (g18372));
OR2X1 gate16061(.O (g25682), .I1 (g24658), .I2 (g18640));
OR2X1 gate16062(.O (g29274), .I1 (g28360), .I2 (g18642));
OR2X1 gate16063(.O (g24561), .I1 (I23755), .I2 (I23756));
OR2X1 gate16064(.O (g24353), .I1 (g23682), .I2 (g18822));
OR2X1 gate16065(.O (g26903), .I1 (g26388), .I2 (g24220));
OR2X1 gate16066(.O (g35000), .I1 (g34953), .I2 (g34999));
OR2X1 gate16067(.O (g11737), .I1 (g8359), .I2 (g8292));
OR2X1 gate16068(.O (g9012), .I1 (g2047), .I2 (g2066));
OR2X1 gate16069(.O (g26755), .I1 (g10776), .I2 (g24457));
OR2X1 gate16070(.O (g28511), .I1 (g27272), .I2 (g16208));
OR2X1 gate16071(.O (g32229), .I1 (g31148), .I2 (g29652));
OR2X1 gate16072(.O (g26770), .I1 (g24471), .I2 (g10732));
OR2X1 gate16073(.O (g24336), .I1 (g24012), .I2 (g18753));
OR2X1 gate16074(.O (g27837), .I1 (g17401), .I2 (g26725));
OR2X1 gate16075(.O (g33390), .I1 (g32276), .I2 (g29968));
OR2X1 gate16076(.O (g32228), .I1 (g31147), .I2 (g29651));
OR2X1 gate16077(.O (g25760), .I1 (g25238), .I2 (g22109));
OR2X1 gate16078(.O (g29292), .I1 (g28556), .I2 (g18776));
OR2X1 gate16079(.O (g34649), .I1 (g33111), .I2 (g34492));
OR2X1 gate16080(.O (g34240), .I1 (g32910), .I2 (g33958));
OR2X1 gate16081(.O (g30491), .I1 (g30178), .I2 (g21987));
OR2X1 gate16082(.O (g34903), .I1 (g34859), .I2 (g21690));
OR2X1 gate16083(.O (g23297), .I1 (g19692), .I2 (g16178));
OR2X1 gate16084(.O (g34604), .I1 (g34563), .I2 (g15076));
OR2X1 gate16085(.O (g26899), .I1 (g26844), .I2 (g18199));
OR2X1 gate16086(.O (g30563), .I1 (g29347), .I2 (g22134));
OR2X1 gate16087(.O (g26898), .I1 (g26387), .I2 (g18194));
OR2X1 gate16088(.O (g28085), .I1 (g27263), .I2 (g18700));
OR2X1 gate16089(.O (g28076), .I1 (g27098), .I2 (g21878));
OR2X1 gate16090(.O (g28721), .I1 (g27488), .I2 (g16705));
OR2X1 gate16091(.O (g28596), .I1 (g27336), .I2 (g26291));
OR2X1 gate16092(.O (g28054), .I1 (g27723), .I2 (g18170));
OR2X1 gate16093(.O (g33553), .I1 (g33403), .I2 (g18350));
OR2X1 gate16094(.O (g15803), .I1 (g12924), .I2 (g10528));
OR2X1 gate16095(.O (g22217), .I1 (g21302), .I2 (g17617));
OR2X1 gate16096(.O (g33949), .I1 (g32446), .I2 (g33459));
OR2X1 gate16097(.O (g31326), .I1 (g29627), .I2 (g29640));
OR2X1 gate16098(.O (g32386), .I1 (g31488), .I2 (g29949));
OR2X1 gate16099(.O (g30395), .I1 (g29841), .I2 (g21754));
OR2X1 gate16100(.O (g34794), .I1 (g34746), .I2 (g18571));
OR2X1 gate16101(.O (g25649), .I1 (g24654), .I2 (g21742));
OR4X1 gate16102(.O (I26644), .I1 (g27057), .I2 (g27044), .I3 (g27039), .I4 (g27032));
OR4X1 gate16103(.O (g27037), .I1 (g26236), .I2 (g26218), .I3 (g26195), .I4 (g26171));
OR2X1 gate16104(.O (g34262), .I1 (g34075), .I2 (g18697));
OR2X1 gate16105(.O (g33536), .I1 (g33241), .I2 (g21715));
OR2X1 gate16106(.O (g33040), .I1 (g32164), .I2 (g24313));
OR2X1 gate16107(.O (g33948), .I1 (g32442), .I2 (g33458));
OR2X1 gate16108(.O (g25648), .I1 (g24644), .I2 (g21741));
OR2X1 gate16109(.O (g28773), .I1 (g27535), .I2 (g16803));
OR2X1 gate16110(.O (g31757), .I1 (g29992), .I2 (g30010));
OR2X1 gate16111(.O (g31904), .I1 (g31780), .I2 (g21923));
OR2X1 gate16112(.O (g34633), .I1 (g34481), .I2 (g18690));
OR2X1 gate16113(.O (g25604), .I1 (g24717), .I2 (g18115));
OR2X1 gate16114(.O (g25755), .I1 (g25192), .I2 (g22102));
OR2X1 gate16115(.O (g33621), .I1 (g33365), .I2 (g18775));
OR2X1 gate16116(.O (g34719), .I1 (g34701), .I2 (g18133));
OR2X1 gate16117(.O (g28180), .I1 (g20242), .I2 (g27511));
OR2X1 gate16118(.O (g28670), .I1 (g27412), .I2 (g16618));
OR2X1 gate16119(.O (g26926), .I1 (g26633), .I2 (g18531));
OR2X1 gate16120(.O (g32429), .I1 (g30318), .I2 (g31794));
OR2X1 gate16121(.O (g30521), .I1 (g29331), .I2 (g22042));
OR2X1 gate16122(.O (g14511), .I1 (g10685), .I2 (g546));
OR2X1 gate16123(.O (g33564), .I1 (g33332), .I2 (g18388));
OR2X1 gate16124(.O (g26099), .I1 (g24506), .I2 (g22538));
OR2X1 gate16125(.O (g29283), .I1 (g28627), .I2 (g18746));
OR2X1 gate16126(.O (g28734), .I1 (g27508), .I2 (g16736));
OR2X1 gate16127(.O (g28335), .I1 (g27132), .I2 (g15818));
OR2X1 gate16128(.O (g29303), .I1 (g28703), .I2 (g18801));
OR2X1 gate16129(.O (g24374), .I1 (g19345), .I2 (g24004));
OR2X1 gate16130(.O (g30440), .I1 (g29771), .I2 (g21849));
OR2X1 gate16131(.O (g34440), .I1 (g34364), .I2 (g24226));
OR2X1 gate16132(.O (g25767), .I1 (g25207), .I2 (g12015));
OR2X1 gate16133(.O (g28667), .I1 (g27410), .I2 (g16616));
OR2X1 gate16134(.O (g33062), .I1 (g31977), .I2 (g22065));
OR2X1 gate16135(.O (g22531), .I1 (g20773), .I2 (g20922));
OR2X1 gate16136(.O (g27589), .I1 (g26177), .I2 (g24763));
OR2X1 gate16137(.O (g16448), .I1 (g13287), .I2 (g10934));
OR2X1 gate16138(.O (g30389), .I1 (g29969), .I2 (g18554));
OR2X1 gate16139(.O (g24260), .I1 (g23373), .I2 (g18313));
OR2X1 gate16140(.O (g27524), .I1 (g26050), .I2 (g24649));
OR2X1 gate16141(.O (g25633), .I1 (g24420), .I2 (g18282));
OR2X1 gate16142(.O (g31872), .I1 (g31524), .I2 (g18535));
OR2X1 gate16143(.O (g24842), .I1 (g7804), .I2 (g22669));
OR2X1 gate16144(.O (g30388), .I1 (g30023), .I2 (g18534));
OR2X1 gate16145(.O (g34612), .I1 (g34514), .I2 (g18566));
OR2X1 gate16146(.O (g25719), .I1 (g25089), .I2 (g18761));
OR2X1 gate16147(.O (g28619), .I1 (g27358), .I2 (g16517));
OR2X1 gate16148(.O (g34099), .I1 (g33684), .I2 (g33689));
OR2X1 gate16149(.O (g30534), .I1 (g30213), .I2 (g22080));
OR2X1 gate16150(.O (g19441), .I1 (g15507), .I2 (g12931));
OR2X1 gate16151(.O (g25718), .I1 (g25187), .I2 (g21971));
OR2X1 gate16152(.O (g28618), .I1 (g27357), .I2 (g16516));
OR2X1 gate16153(.O (g34251), .I1 (g34157), .I2 (g18147));
OR2X1 gate16154(.O (g28279), .I1 (g27087), .I2 (g25909));
OR2X1 gate16155(.O (g26766), .I1 (g10776), .I2 (g24460));
OR2X1 gate16156(.O (g30462), .I1 (g30228), .I2 (g21933));
OR2X1 gate16157(.O (g23296), .I1 (g19691), .I2 (g16177));
OR2X1 gate16158(.O (g34462), .I1 (g34334), .I2 (g18685));
OR2X1 gate16159(.O (g28286), .I1 (g27090), .I2 (g15757));
OR2X1 gate16160(.O (g32245), .I1 (g31167), .I2 (g29684));
OR2X1 gate16161(.O (g34032), .I1 (g33816), .I2 (g18706));
OR2X1 gate16162(.O (g28306), .I1 (g27104), .I2 (g15794));
OR2X1 gate16163(.O (g33574), .I1 (g33362), .I2 (g18416));
OR2X1 gate16164(.O (g33047), .I1 (g31944), .I2 (g21927));
OR4X1 gate16165(.O (I26741), .I1 (g22881), .I2 (g22905), .I3 (g22928), .I4 (g27402));
OR2X1 gate16166(.O (g31912), .I1 (g31752), .I2 (g21998));
OR2X1 gate16167(.O (g31311), .I1 (g26103), .I2 (g29618));
OR2X1 gate16168(.O (g23197), .I1 (g19571), .I2 (g15966));
OR2X1 gate16169(.O (g25612), .I1 (g24941), .I2 (g18132));
OR2X1 gate16170(.O (g28815), .I1 (g27546), .I2 (g16842));
OR2X1 gate16171(.O (g29483), .I1 (g25801), .I2 (g28130));
OR2X1 gate16172(.O (g16811), .I1 (g8690), .I2 (g13914));
OR2X1 gate16173(.O (g25701), .I1 (g25054), .I2 (g21920));
OR4X1 gate16174(.O (I30055), .I1 (g31070), .I2 (g31170), .I3 (g30614), .I4 (g30673));
OR2X1 gate16175(.O (g24705), .I1 (g2890), .I2 (g23267));
OR2X1 gate16176(.O (g33051), .I1 (g32316), .I2 (g21958));
OR2X1 gate16177(.O (g24255), .I1 (g22835), .I2 (g18308));
OR2X1 gate16178(.O (g33592), .I1 (g33412), .I2 (g18475));
OR2X1 gate16179(.O (g30360), .I1 (g30145), .I2 (g18386));
OR2X1 gate16180(.O (g24270), .I1 (g23165), .I2 (g18614));
OR2X1 gate16181(.O (g26911), .I1 (g26612), .I2 (g24230));
OR4X1 gate16182(.O (I30741), .I1 (g32085), .I2 (g32030), .I3 (g32224), .I4 (g32013));
OR2X1 gate16183(.O (g30447), .I1 (g29798), .I2 (g21856));
OR2X1 gate16184(.O (g21894), .I1 (g20112), .I2 (g15107));
OR2X1 gate16185(.O (g34447), .I1 (g34363), .I2 (g18552));
OR2X1 gate16186(.O (g32995), .I1 (g32330), .I2 (g18375));
OR2X1 gate16187(.O (g24460), .I1 (g10967), .I2 (g22450));
OR2X1 gate16188(.O (g29904), .I1 (g28312), .I2 (g26146));
OR2X1 gate16189(.O (g13657), .I1 (g7251), .I2 (g10616));
OR2X1 gate16190(.O (g29252), .I1 (g28712), .I2 (g18486));
OR2X1 gate16191(.O (g28884), .I1 (g27568), .I2 (g16885));
OR2X1 gate16192(.O (g26785), .I1 (g10776), .I2 (g24468));
OR2X1 gate16193(.O (g24267), .I1 (g23439), .I2 (g18611));
OR2X1 gate16194(.O (g30451), .I1 (g29877), .I2 (g21860));
OR2X1 gate16195(.O (g30472), .I1 (g30186), .I2 (g21943));
OR4X1 gate16196(.O (I30735), .I1 (g32369), .I2 (g32376), .I3 (g32089), .I4 (g32035));
OR2X1 gate16197(.O (g34629), .I1 (g34495), .I2 (g18654));
OR4X1 gate16198(.O (g17569), .I1 (g14416), .I2 (g14394), .I3 (g11995), .I4 (I18492));
OR2X1 gate16199(.O (g34451), .I1 (g34393), .I2 (g18664));
OR2X1 gate16200(.O (g34628), .I1 (g34493), .I2 (g18653));
OR2X1 gate16201(.O (g34911), .I1 (g34909), .I2 (g18188));
OR2X1 gate16202(.O (g26950), .I1 (g26357), .I2 (g24288));
OR2X1 gate16203(.O (g22751), .I1 (g19333), .I2 (g15716));
OR3X1 gate16204(.O (g27008), .I1 (g26866), .I2 (g21370), .I3 (I25736));
OR2X1 gate16205(.O (g22639), .I1 (g18950), .I2 (g15612));
OR2X1 gate16206(.O (g27555), .I1 (g26095), .I2 (g24686));
OR2X1 gate16207(.O (g28580), .I1 (g27328), .I2 (g26275));
OR2X1 gate16208(.O (g29508), .I1 (g28152), .I2 (g27041));
OR3X1 gate16209(.O (g8476), .I1 (g1399), .I2 (g1459), .I3 (I12611));
OR2X1 gate16210(.O (g20160), .I1 (g16163), .I2 (g13415));
OR2X1 gate16211(.O (g30355), .I1 (g30131), .I2 (g18360));
OR2X1 gate16212(.O (g27570), .I1 (g26126), .I2 (g24722));
OR2X1 gate16213(.O (g31929), .I1 (g31540), .I2 (g22093));
OR2X1 gate16214(.O (g32989), .I1 (g32241), .I2 (g18326));
OR2X1 gate16215(.O (g30370), .I1 (g30135), .I2 (g18440));
OR2X1 gate16216(.O (g25629), .I1 (g24962), .I2 (g18258));
OR2X1 gate16217(.O (g27907), .I1 (g17424), .I2 (g26770));
OR2X1 gate16218(.O (g16959), .I1 (g13542), .I2 (g11142));
OR2X1 gate16219(.O (g31020), .I1 (g29375), .I2 (g28164));
OR2X1 gate16220(.O (g31928), .I1 (g31517), .I2 (g22092));
OR2X1 gate16221(.O (g14187), .I1 (g8871), .I2 (g11771));
OR2X1 gate16222(.O (g32988), .I1 (g32232), .I2 (g18325));
OR2X1 gate16223(.O (g28084), .I1 (g27254), .I2 (g18698));
OR2X1 gate16224(.O (g33020), .I1 (g32160), .I2 (g21734));
OR2X1 gate16225(.O (g33583), .I1 (g33074), .I2 (g18448));
OR2X1 gate16226(.O (g25628), .I1 (g24600), .I2 (g18249));
OR2X1 gate16227(.O (g25911), .I1 (g22514), .I2 (g24510));
OR2X1 gate16228(.O (g27239), .I1 (g25881), .I2 (g24465));
OR2X1 gate16229(.O (g19605), .I1 (g15707), .I2 (g13063));
OR2X1 gate16230(.O (g33046), .I1 (g32308), .I2 (g21912));
OR2X1 gate16231(.O (g32271), .I1 (g31209), .I2 (g29731));
OR2X1 gate16232(.O (g34172), .I1 (g33795), .I2 (g19914));
OR4X1 gate16233(.O (g28179), .I1 (g27494), .I2 (g27474), .I3 (g27445), .I4 (g27421));
OR2X1 gate16234(.O (g27567), .I1 (g26121), .I2 (g24714));
OR2X1 gate16235(.O (g27238), .I1 (g25879), .I2 (g24464));
OR4X1 gate16236(.O (g17510), .I1 (g14393), .I2 (g14362), .I3 (g11972), .I4 (I18449));
OR2X1 gate16237(.O (g30394), .I1 (g29805), .I2 (g21753));
OR2X1 gate16238(.O (g30367), .I1 (g30133), .I2 (g18418));
OR2X1 gate16239(.O (g24201), .I1 (g22848), .I2 (g18104));
OR2X1 gate16240(.O (g24277), .I1 (g23188), .I2 (g18647));
OR2X1 gate16241(.O (g25591), .I1 (g24642), .I2 (g21705));
OR2X1 gate16242(.O (g33282), .I1 (g32143), .I2 (g29577));
OR4X1 gate16243(.O (g28186), .I1 (g27209), .I2 (g27185), .I3 (g27161), .I4 (g27146));
OR2X1 gate16244(.O (g28685), .I1 (g27433), .I2 (g16637));
OR2X1 gate16245(.O (g31302), .I1 (g29590), .I2 (g28302));
OR2X1 gate16246(.O (g28373), .I1 (g27180), .I2 (g15849));
OR2X1 gate16247(.O (g25754), .I1 (g25179), .I2 (g22101));
OR2X1 gate16248(.O (g30420), .I1 (g29769), .I2 (g21804));
OR2X1 gate16249(.O (g28417), .I1 (g27219), .I2 (g15881));
OR2X1 gate16250(.O (g24782), .I1 (g23857), .I2 (g23872));
OR2X1 gate16251(.O (g30446), .I1 (g29788), .I2 (g21855));
OR2X1 gate16252(.O (g34446), .I1 (g34390), .I2 (g18550));
OR2X1 gate16253(.O (g34318), .I1 (g25850), .I2 (g34063));
OR2X1 gate16254(.O (g28334), .I1 (g27131), .I2 (g15817));
OR2X1 gate16255(.O (g29756), .I1 (g22717), .I2 (g28223));
OR2X1 gate16256(.O (g24352), .I1 (g22157), .I2 (g18821));
OR2X1 gate16257(.O (g26902), .I1 (g26378), .I2 (g24219));
OR2X1 gate16258(.O (g26957), .I1 (g26517), .I2 (g24295));
OR2X1 gate16259(.O (g34025), .I1 (g33927), .I2 (g18672));
OR2X1 gate16260(.O (g31768), .I1 (g30033), .I2 (g30045));
OR2X1 gate16261(.O (g26377), .I1 (g24700), .I2 (g23007));
OR2X1 gate16262(.O (g30540), .I1 (g30275), .I2 (g22086));
OR2X1 gate16263(.O (g13295), .I1 (g10625), .I2 (g10655));
OR2X1 gate16264(.O (g15582), .I1 (g8977), .I2 (g12925));
OR2X1 gate16265(.O (g24266), .I1 (g22329), .I2 (g18561));
OR2X1 gate16266(.O (g32132), .I1 (g31487), .I2 (g31479));
OR2X1 gate16267(.O (g9535), .I1 (g209), .I2 (g538));
OR2X1 gate16268(.O (g31881), .I1 (g31018), .I2 (g21775));
OR2X1 gate16269(.O (g28216), .I1 (g27036), .I2 (g27043));
OR2X1 gate16270(.O (g24853), .I1 (g21452), .I2 (g24001));
OR2X1 gate16271(.O (g22684), .I1 (g19206), .I2 (g15703));
OR2X1 gate16272(.O (g32259), .I1 (g31185), .I2 (g29709));
OR2X1 gate16273(.O (g30377), .I1 (g30124), .I2 (g18472));
OR2X1 gate16274(.O (g32225), .I1 (g30576), .I2 (g29336));
OR2X1 gate16275(.O (g34957), .I1 (g34948), .I2 (g21662));
OR2X1 gate16276(.O (g34377), .I1 (g26304), .I2 (g34141));
OR2X1 gate16277(.O (g33027), .I1 (g32314), .I2 (g21796));
OR3X1 gate16278(.O (I22912), .I1 (g21555), .I2 (g21364), .I3 (g21357));
OR2X1 gate16279(.O (g31890), .I1 (g31143), .I2 (g21823));
OR2X1 gate16280(.O (g24401), .I1 (g23811), .I2 (g21298));
OR2X1 gate16281(.O (g30562), .I1 (g30289), .I2 (g22133));
OR2X1 gate16282(.O (g31249), .I1 (g25971), .I2 (g29523));
OR2X1 gate16283(.O (g19359), .I1 (g17786), .I2 (g14875));
OR2X1 gate16284(.O (g34645), .I1 (g34556), .I2 (g18786));
OR2X1 gate16285(.O (g19535), .I1 (g15651), .I2 (g13020));
OR2X1 gate16286(.O (g31248), .I1 (g25970), .I2 (g29522));
OR2X1 gate16287(.O (g28747), .I1 (g27521), .I2 (g13942));
OR2X1 gate16288(.O (g34290), .I1 (g26848), .I2 (g34219));
OR2X1 gate16289(.O (g33552), .I1 (g33400), .I2 (g18343));
OR2X1 gate16290(.O (g13289), .I1 (g10619), .I2 (g10624));
OR2X1 gate16291(.O (g33003), .I1 (g32323), .I2 (g18429));
OR3X1 gate16292(.O (g33204), .I1 (g32317), .I2 (I30750), .I3 (I30751));
OR2X1 gate16293(.O (g26895), .I1 (g26783), .I2 (g18148));
OR2X1 gate16294(.O (g31779), .I1 (g30050), .I2 (g28673));
OR4X1 gate16295(.O (I31843), .I1 (g33470), .I2 (g33471), .I3 (g33472), .I4 (g33473));
OR2X1 gate16296(.O (g10800), .I1 (g7517), .I2 (g952));
OR2X1 gate16297(.O (g19344), .I1 (g17771), .I2 (g14832));
OR2X1 gate16298(.O (g27566), .I1 (g26119), .I2 (g24713));
OR2X1 gate16299(.O (g28814), .I1 (g27545), .I2 (g16841));
OR2X1 gate16300(.O (g30427), .I1 (g29796), .I2 (g21811));
OR2X1 gate16301(.O (g20276), .I1 (g16243), .I2 (g13566));
OR2X1 gate16302(.O (g29583), .I1 (g28182), .I2 (g27099));
OR2X1 gate16303(.O (g32375), .I1 (g29896), .I2 (g31324));
OR2X1 gate16304(.O (g14936), .I1 (g10776), .I2 (g8703));
OR2X1 gate16305(.O (g30366), .I1 (g30122), .I2 (g18417));
OR4X1 gate16306(.O (I30054), .I1 (g29385), .I2 (g31376), .I3 (g30735), .I4 (g30825));
OR2X1 gate16307(.O (g24276), .I1 (g23083), .I2 (g18646));
OR2X1 gate16308(.O (g28751), .I1 (g27526), .I2 (g16766));
OR2X1 gate16309(.O (g28772), .I1 (g27534), .I2 (g16802));
OR2X1 gate16310(.O (g34366), .I1 (g26257), .I2 (g34133));
OR4X1 gate16311(.O (I31869), .I1 (g33519), .I2 (g33520), .I3 (g33521), .I4 (g33522));
OR2X1 gate16312(.O (g34632), .I1 (g34565), .I2 (g15119));
OR2X1 gate16313(.O (g25739), .I1 (g25149), .I2 (g22054));
OR2X1 gate16314(.O (g24254), .I1 (g23265), .I2 (g18306));
OR4X1 gate16315(.O (I31868), .I1 (g33515), .I2 (g33516), .I3 (g33517), .I4 (g33518));
OR2X1 gate16316(.O (g28230), .I1 (g27669), .I2 (g14261));
OR2X1 gate16317(.O (g33945), .I1 (g32430), .I2 (g33455));
OR2X1 gate16318(.O (g25738), .I1 (g25059), .I2 (g22053));
OR2X1 gate16319(.O (g25645), .I1 (g24679), .I2 (g21738));
OR2X1 gate16320(.O (g30547), .I1 (g30194), .I2 (g22118));
OR2X1 gate16321(.O (g30403), .I1 (g29750), .I2 (g21762));
OR2X1 gate16322(.O (g33999), .I1 (g33893), .I2 (g18436));
OR2X1 gate16323(.O (g33380), .I1 (g32234), .I2 (g29926));
OR2X1 gate16324(.O (g25699), .I1 (g25125), .I2 (g21918));
OR2X1 gate16325(.O (g34403), .I1 (g34180), .I2 (g25085));
OR2X1 gate16326(.O (g29282), .I1 (g28617), .I2 (g18745));
OR2X1 gate16327(.O (g28416), .I1 (g27218), .I2 (g15880));
OR2X1 gate16328(.O (g16261), .I1 (g7898), .I2 (g13469));
OR2X1 gate16329(.O (g32994), .I1 (g32290), .I2 (g18367));
OR2X1 gate16330(.O (g33998), .I1 (g33878), .I2 (g18428));
OR2X1 gate16331(.O (g29302), .I1 (g28601), .I2 (g18798));
OR2X1 gate16332(.O (g25698), .I1 (g25104), .I2 (g21917));
OR2X1 gate16333(.O (g29105), .I1 (g27645), .I2 (g17134));
OR2X1 gate16334(.O (g30481), .I1 (g30221), .I2 (g21977));
OR2X1 gate16335(.O (g7932), .I1 (g4072), .I2 (g4153));
OR2X1 gate16336(.O (g26956), .I1 (g26487), .I2 (g24294));
OR2X1 gate16337(.O (g30551), .I1 (g30235), .I2 (g22122));
OR4X1 gate16338(.O (I30734), .I1 (g31790), .I2 (g32191), .I3 (g32086), .I4 (g32095));
OR2X1 gate16339(.O (g26889), .I1 (g26689), .I2 (g24195));
OR2X1 gate16340(.O (g31932), .I1 (g31792), .I2 (g22107));
OR2X1 gate16341(.O (g26888), .I1 (g26671), .I2 (g24194));
OR3X1 gate16342(.O (g23721), .I1 (g21401), .I2 (g21385), .I3 (I22852));
OR2X1 gate16343(.O (g25632), .I1 (g24558), .I2 (g18277));
OR2X1 gate16344(.O (g28578), .I1 (g27327), .I2 (g26273));
OR2X1 gate16345(.O (g30127), .I1 (g28494), .I2 (g16805));
OR2X1 gate16346(.O (g29768), .I1 (g22760), .I2 (g28229));
OR2X1 gate16347(.O (g34127), .I1 (g33657), .I2 (g32438));
OR2X1 gate16348(.O (g31897), .I1 (g31237), .I2 (g24322));
OR2X1 gate16349(.O (g30490), .I1 (g30167), .I2 (g21986));
OR2X1 gate16350(.O (g33961), .I1 (g33789), .I2 (g21712));
OR2X1 gate16351(.O (g25661), .I1 (g24754), .I2 (g21786));
OR2X1 gate16352(.O (g27484), .I1 (g25988), .I2 (g24628));
OR2X1 gate16353(.O (g30376), .I1 (g30112), .I2 (g18471));
OR2X1 gate16354(.O (g30385), .I1 (g30172), .I2 (g18518));
OR2X1 gate16355(.O (g26931), .I1 (g26778), .I2 (g18547));
OR2X1 gate16356(.O (g30103), .I1 (g28477), .I2 (g16731));
OR2X1 gate16357(.O (g34376), .I1 (g26301), .I2 (g34140));
OR2X1 gate16358(.O (g34297), .I1 (g26858), .I2 (g34228));
OR2X1 gate16359(.O (g34103), .I1 (g33701), .I2 (g33707));
OR2X1 gate16360(.O (g33026), .I1 (g32307), .I2 (g21795));
OR2X1 gate16361(.O (g30354), .I1 (g30064), .I2 (g18359));
OR2X1 gate16362(.O (g22516), .I1 (g21559), .I2 (g12817));
OR2X1 gate16363(.O (g34980), .I1 (g34969), .I2 (g18587));
OR3X1 gate16364(.O (g33212), .I1 (g32328), .I2 (I30755), .I3 (I30756));
OR2X1 gate16365(.O (g25715), .I1 (g25071), .I2 (g21966));
OR2X1 gate16366(.O (g8679), .I1 (g222), .I2 (g199));
OR2X1 gate16367(.O (g34095), .I1 (g33681), .I2 (g33687));
OR2X1 gate16368(.O (g30824), .I1 (g13833), .I2 (g29789));
OR2X1 gate16369(.O (g28720), .I1 (g27486), .I2 (g16704));
OR2X1 gate16370(.O (g28041), .I1 (g24145), .I2 (g26878));
OR2X1 gate16371(.O (g17264), .I1 (g7118), .I2 (g14309));
OR2X1 gate16372(.O (g28430), .I1 (g27229), .I2 (g15914));
OR2X1 gate16373(.O (g32125), .I1 (g30918), .I2 (g29376));
OR2X1 gate16374(.O (g28746), .I1 (g27520), .I2 (g16762));
OR2X1 gate16375(.O (g32977), .I1 (g32169), .I2 (g21710));
OR2X1 gate16376(.O (g19604), .I1 (g15704), .I2 (g13059));
OR4X1 gate16377(.O (I30469), .I1 (g31672), .I2 (g31710), .I3 (g31021), .I4 (g30937));
OR2X1 gate16378(.O (g29249), .I1 (g28658), .I2 (g18438));
OR2X1 gate16379(.O (g26089), .I1 (g24501), .I2 (g22534));
OR2X1 gate16380(.O (g24907), .I1 (g21558), .I2 (g24015));
OR4X1 gate16381(.O (I30468), .I1 (g29385), .I2 (g31376), .I3 (g30735), .I4 (g30825));
OR2X1 gate16382(.O (g29482), .I1 (g28524), .I2 (g27588));
OR2X1 gate16383(.O (g34931), .I1 (g2984), .I2 (g34912));
OR2X1 gate16384(.O (g29248), .I1 (g28677), .I2 (g18434));
OR3X1 gate16385(.O (g33149), .I1 (g32204), .I2 (I30717), .I3 (I30718));
OR2X1 gate16386(.O (g30426), .I1 (g29785), .I2 (g21810));
OR2X1 gate16387(.O (g32353), .I1 (g29853), .I2 (g31283));
OR2X1 gate16388(.O (g33387), .I1 (g32263), .I2 (g29954));
OR2X1 gate16389(.O (g24239), .I1 (g22752), .I2 (g18250));
OR2X1 gate16390(.O (g9055), .I1 (g2606), .I2 (g2625));
OR2X1 gate16391(.O (g28684), .I1 (g27432), .I2 (g16636));
OR2X1 gate16392(.O (g32144), .I1 (g30927), .I2 (g30930));
OR2X1 gate16393(.O (g33620), .I1 (g33360), .I2 (g18774));
OR2X1 gate16394(.O (g34190), .I1 (g33802), .I2 (g33810));
OR2X1 gate16395(.O (g24238), .I1 (g23254), .I2 (g18248));
OR2X1 gate16396(.O (g30520), .I1 (g30272), .I2 (g22041));
OR2X1 gate16397(.O (g28517), .I1 (g27280), .I2 (g26154));
OR2X1 gate16398(.O (g30546), .I1 (g30277), .I2 (g22117));
OR2X1 gate16399(.O (g33971), .I1 (g33890), .I2 (g18330));
OR2X1 gate16400(.O (g29786), .I1 (g22843), .I2 (g28240));
OR2X1 gate16401(.O (g25671), .I1 (g24637), .I2 (g21828));
OR2X1 gate16402(.O (g34024), .I1 (g33807), .I2 (g24331));
OR2X1 gate16403(.O (g13938), .I1 (g11213), .I2 (g11191));
OR2X1 gate16404(.O (g24518), .I1 (g22517), .I2 (g7601));
OR2X1 gate16405(.O (g22530), .I1 (g16751), .I2 (g20171));
OR2X1 gate16406(.O (g28362), .I1 (g27154), .I2 (g15840));
OR2X1 gate16407(.O (g30497), .I1 (g30242), .I2 (g21993));
OR2X1 gate16408(.O (g24935), .I1 (g22937), .I2 (g19749));
OR4X1 gate16409(.O (I12903), .I1 (g4222), .I2 (g4219), .I3 (g4216), .I4 (g4213));
OR2X1 gate16410(.O (g29233), .I1 (g28171), .I2 (g18234));
OR2X1 gate16411(.O (g26969), .I1 (g26313), .I2 (g24329));
OR3X1 gate16412(.O (I18421), .I1 (g14447), .I2 (g14417), .I3 (g14395));
OR2X1 gate16413(.O (g32289), .I1 (g24796), .I2 (g31230));
OR2X1 gate16414(.O (g22641), .I1 (g18974), .I2 (g15631));
OR2X1 gate16415(.O (g34625), .I1 (g34532), .I2 (g18610));
OR2X1 gate16416(.O (g26968), .I1 (g26307), .I2 (g24321));
OR4X1 gate16417(.O (g17464), .I1 (g14334), .I2 (g14313), .I3 (g11935), .I4 (I18385));
OR2X1 gate16418(.O (g31896), .I1 (g31242), .I2 (g24305));
OR2X1 gate16419(.O (g34250), .I1 (g34111), .I2 (g21713));
OR2X1 gate16420(.O (g32288), .I1 (g31226), .I2 (g31229));
OR2X1 gate16421(.O (g28727), .I1 (g27500), .I2 (g16729));
OR2X1 gate16422(.O (g16258), .I1 (g13247), .I2 (g10856));
OR2X1 gate16423(.O (g33011), .I1 (g32338), .I2 (g18481));
OR2X1 gate16424(.O (g30339), .I1 (g29629), .I2 (g18244));
OR2X1 gate16425(.O (g24215), .I1 (g23484), .I2 (g18196));
OR2X1 gate16426(.O (g24577), .I1 (g2856), .I2 (g22531));
OR2X1 gate16427(.O (g30338), .I1 (g29613), .I2 (g18240));
OR2X1 gate16428(.O (g34644), .I1 (g34555), .I2 (g18769));
OR2X1 gate16429(.O (g33582), .I1 (g33351), .I2 (g18444));
OR2X1 gate16430(.O (g19534), .I1 (g15650), .I2 (g13019));
OR2X1 gate16431(.O (g27241), .I1 (g24584), .I2 (g25984));
OR2X1 gate16432(.O (g28347), .I1 (g27138), .I2 (g15822));
OR2X1 gate16433(.O (g29717), .I1 (g28200), .I2 (g10883));
OR2X1 gate16434(.O (g33310), .I1 (g29631), .I2 (g32165));
OR2X1 gate16435(.O (g26894), .I1 (g25979), .I2 (g18129));
OR2X1 gate16436(.O (g33627), .I1 (g33376), .I2 (g18826));
OR2X1 gate16437(.O (g31925), .I1 (g31789), .I2 (g22061));
OR2X1 gate16438(.O (g32976), .I1 (g32207), .I2 (g21704));
OR2X1 gate16439(.O (g32985), .I1 (g31963), .I2 (g18266));
OR2X1 gate16440(.O (g24349), .I1 (g23646), .I2 (g18805));
OR2X1 gate16441(.O (g16810), .I1 (g13461), .I2 (g11032));
OR2X1 gate16442(.O (g25700), .I1 (g25040), .I2 (g21919));
OR2X1 gate16443(.O (g28600), .I1 (g27339), .I2 (g16427));
OR2X1 gate16444(.O (g25659), .I1 (g24707), .I2 (g21784));
OR2X1 gate16445(.O (g25625), .I1 (g24553), .I2 (g18226));
OR2X1 gate16446(.O (g20083), .I1 (g2902), .I2 (g17058));
OR2X1 gate16447(.O (g30527), .I1 (g30192), .I2 (g22073));
OR2X1 gate16448(.O (g30411), .I1 (g29872), .I2 (g21770));
OR2X1 gate16449(.O (g33050), .I1 (g31974), .I2 (g21930));
OR2X1 gate16450(.O (g32374), .I1 (g29895), .I2 (g31323));
OR3X1 gate16451(.O (g33958), .I1 (g33532), .I2 (I31873), .I3 (I31874));
OR2X1 gate16452(.O (g24348), .I1 (g22149), .I2 (g18804));
OR2X1 gate16453(.O (g34411), .I1 (g34186), .I2 (g25142));
OR2X1 gate16454(.O (g16970), .I1 (g13567), .I2 (g11163));
OR2X1 gate16455(.O (g25658), .I1 (g24635), .I2 (g21783));
OR2X1 gate16456(.O (g28372), .I1 (g27178), .I2 (g15848));
OR2X1 gate16457(.O (g23217), .I1 (g19588), .I2 (g16023));
OR2X1 gate16458(.O (g33386), .I1 (g32258), .I2 (g29951));
OR2X1 gate16459(.O (g26910), .I1 (g26571), .I2 (g24228));
OR2X1 gate16460(.O (g33603), .I1 (g33372), .I2 (g18515));
OR2X1 gate16461(.O (g25943), .I1 (g24423), .I2 (g22299));
OR4X1 gate16462(.O (I30740), .I1 (g31776), .I2 (g32188), .I3 (g32083), .I4 (g32087));
OR2X1 gate16463(.O (g13623), .I1 (g482), .I2 (g12527));
OR2X1 gate16464(.O (g25644), .I1 (g24622), .I2 (g21737));
OR2X1 gate16465(.O (g30503), .I1 (g30243), .I2 (g22024));
OR2X1 gate16466(.O (g28063), .I1 (g27541), .I2 (g21773));
OR2X1 gate16467(.O (g34894), .I1 (g34862), .I2 (g21678));
OR2X1 gate16468(.O (g29148), .I1 (g27651), .I2 (g26606));
OR2X1 gate16469(.O (g32392), .I1 (g31513), .I2 (g30000));
OR2X1 gate16470(.O (g27515), .I1 (g26051), .I2 (g13431));
OR2X1 gate16471(.O (g30450), .I1 (g29861), .I2 (g21859));
OR2X1 gate16472(.O (g24653), .I1 (g2848), .I2 (g22585));
OR2X1 gate16473(.O (g34450), .I1 (g34281), .I2 (g18663));
OR2X1 gate16474(.O (g13155), .I1 (g11496), .I2 (g11546));
OR2X1 gate16475(.O (g31793), .I1 (g28031), .I2 (g30317));
OR2X1 gate16476(.O (g34819), .I1 (g34741), .I2 (g34684));
OR2X1 gate16477(.O (g34257), .I1 (g34226), .I2 (g18674));
OR2X1 gate16478(.O (g28209), .I1 (g27223), .I2 (g27141));
OR2X1 gate16479(.O (g30496), .I1 (g30231), .I2 (g21992));
OR2X1 gate16480(.O (g8956), .I1 (g1913), .I2 (g1932));
OR2X1 gate16481(.O (g34979), .I1 (g34875), .I2 (g34968));
OR2X1 gate16482(.O (g34055), .I1 (g33909), .I2 (g33910));
OR2X1 gate16483(.O (g33549), .I1 (g33328), .I2 (g18337));
OR2X1 gate16484(.O (g28208), .I1 (g27025), .I2 (g27028));
OR2X1 gate16485(.O (g26877), .I1 (g21658), .I2 (g25577));
OR2X1 gate16486(.O (g34978), .I1 (g34874), .I2 (g34967));
OR2X1 gate16487(.O (g33548), .I1 (g33327), .I2 (g18336));
OR2X1 gate16488(.O (g27584), .I1 (g26165), .I2 (g24758));
OR2X1 gate16489(.O (g25867), .I1 (g25449), .I2 (g23884));
OR2X1 gate16490(.O (g25894), .I1 (g24817), .I2 (g23229));
OR2X1 gate16491(.O (g30384), .I1 (g30101), .I2 (g18517));
OR2X1 gate16492(.O (g31317), .I1 (g29611), .I2 (g29626));
OR2X1 gate16493(.O (g33317), .I1 (g29688), .I2 (g32179));
OR2X1 gate16494(.O (g29229), .I1 (g28532), .I2 (g18191));
OR2X1 gate16495(.O (g25714), .I1 (g25056), .I2 (g21965));
OR2X1 gate16496(.O (g28614), .I1 (g27351), .I2 (g26311));
OR2X1 gate16497(.O (g25707), .I1 (g25041), .I2 (g18749));
OR2X1 gate16498(.O (g25819), .I1 (g25323), .I2 (g23836));
OR2X1 gate16499(.O (g28607), .I1 (g27342), .I2 (g26303));
OR2X1 gate16500(.O (g29228), .I1 (g28426), .I2 (g18173));
OR2X1 gate16501(.O (g25910), .I1 (g25565), .I2 (g22142));
OR2X1 gate16502(.O (g28320), .I1 (g27116), .I2 (g15808));
OR2X1 gate16503(.O (g31002), .I1 (g29362), .I2 (g28154));
OR2X1 gate16504(.O (g28073), .I1 (g27097), .I2 (g21875));
OR2X1 gate16505(.O (g33002), .I1 (g32304), .I2 (g18419));
OR2X1 gate16506(.O (g33057), .I1 (g31968), .I2 (g22019));
OR2X1 gate16507(.O (g34801), .I1 (g34756), .I2 (g18588));
OR2X1 gate16508(.O (g34735), .I1 (g34709), .I2 (g15116));
OR2X1 gate16509(.O (g32124), .I1 (g24488), .I2 (g30920));
OR2X1 gate16510(.O (g29716), .I1 (g28199), .I2 (g15856));
OR2X1 gate16511(.O (g24200), .I1 (g22831), .I2 (g18103));
OR2X1 gate16512(.O (g31245), .I1 (g25964), .I2 (g29516));
OR2X1 gate16513(.O (g34019), .I1 (g33889), .I2 (g18506));
OR2X1 gate16514(.O (g26917), .I1 (g26122), .I2 (g18233));
OR2X1 gate16515(.O (g15792), .I1 (g12920), .I2 (g10501));
OR3X1 gate16516(.O (g26866), .I1 (g20204), .I2 (g20242), .I3 (g24363));
OR2X1 gate16517(.O (g28565), .I1 (g27315), .I2 (g26253));
OR2X1 gate16518(.O (g33626), .I1 (g33374), .I2 (g18825));
OR2X1 gate16519(.O (g33323), .I1 (g31936), .I2 (g32442));
OR2X1 gate16520(.O (g34695), .I1 (g34523), .I2 (g34322));
OR2X1 gate16521(.O (g25590), .I1 (g21694), .I2 (g24160));
OR2X1 gate16522(.O (g34018), .I1 (g33887), .I2 (g18505));
OR2X1 gate16523(.O (g30526), .I1 (g30181), .I2 (g22072));
OR2X1 gate16524(.O (g32267), .I1 (g31208), .I2 (g31218));
OR2X1 gate16525(.O (g32294), .I1 (g31231), .I2 (g31232));
OR2X1 gate16526(.O (g33298), .I1 (g32158), .I2 (g29622));
OR2X1 gate16527(.O (g25741), .I1 (g25178), .I2 (g22056));
OR2X1 gate16528(.O (g28641), .I1 (g27385), .I2 (g16591));
OR2X1 gate16529(.O (g31775), .I1 (g30048), .I2 (g30059));
OR4X1 gate16530(.O (I30123), .I1 (g29385), .I2 (g31376), .I3 (g30735), .I4 (g30825));
OR2X1 gate16531(.O (g8957), .I1 (g2338), .I2 (g2357));
OR2X1 gate16532(.O (g24799), .I1 (g23901), .I2 (g23921));
OR2X1 gate16533(.O (g30402), .I1 (g29871), .I2 (g21761));
OR2X1 gate16534(.O (g24813), .I1 (g22685), .I2 (g19594));
OR4X1 gate16535(.O (I30751), .I1 (g32042), .I2 (g32161), .I3 (g31943), .I4 (g31959));
OR2X1 gate16536(.O (g30457), .I1 (g29369), .I2 (g21885));
OR2X1 gate16537(.O (g34402), .I1 (g34179), .I2 (g25084));
OR2X1 gate16538(.O (g34457), .I1 (g34394), .I2 (g18670));
OR2X1 gate16539(.O (g26923), .I1 (g25923), .I2 (g18290));
OR2X1 gate16540(.O (g32219), .I1 (g31131), .I2 (g29620));
OR2X1 gate16541(.O (g33232), .I1 (g32034), .I2 (g30936));
OR2X1 gate16542(.O (g25735), .I1 (g25077), .I2 (g18783));
OR2X1 gate16543(.O (g25877), .I1 (g25502), .I2 (g23919));
OR2X1 gate16544(.O (g28635), .I1 (g27375), .I2 (g16537));
OR2X1 gate16545(.O (g32218), .I1 (g31130), .I2 (g29619));
OR2X1 gate16546(.O (g27135), .I1 (g24387), .I2 (g25803));
OR2X1 gate16547(.O (g33995), .I1 (g33848), .I2 (g18425));
OR2X1 gate16548(.O (g34001), .I1 (g33844), .I2 (g18450));
OR2X1 gate16549(.O (g33261), .I1 (g32111), .I2 (g29525));
OR2X1 gate16550(.O (g25695), .I1 (g24998), .I2 (g21914));
OR2X1 gate16551(.O (g31880), .I1 (g31280), .I2 (g21774));
OR2X1 gate16552(.O (g30597), .I1 (g13564), .I2 (g29693));
OR2X1 gate16553(.O (g34256), .I1 (g34173), .I2 (g24303));
OR2X1 gate16554(.O (g29802), .I1 (g28243), .I2 (g22871));
OR2X1 gate16555(.O (g34280), .I1 (g26833), .I2 (g34213));
OR2X1 gate16556(.O (g29730), .I1 (g28150), .I2 (g28141));
OR2X1 gate16557(.O (g30300), .I1 (g28246), .I2 (g27252));
OR2X1 gate16558(.O (g29793), .I1 (g28237), .I2 (g27247));
OR2X1 gate16559(.O (g34624), .I1 (g34509), .I2 (g18592));
OR2X1 gate16560(.O (g34300), .I1 (g26864), .I2 (g34230));
OR2X1 gate16561(.O (g15125), .I1 (g10363), .I2 (g13605));
OR2X1 gate16562(.O (g26876), .I1 (g21655), .I2 (g25576));
OR2X1 gate16563(.O (g26885), .I1 (g26541), .I2 (g24191));
OR3X1 gate16564(.O (g23751), .I1 (g21415), .I2 (g21402), .I3 (I22880));
OR2X1 gate16565(.O (g25917), .I1 (g22524), .I2 (g24518));
OR2X1 gate16566(.O (g32277), .I1 (g31211), .I2 (g29733));
OR2X1 gate16567(.O (g24214), .I1 (g23471), .I2 (g18195));
OR2X1 gate16568(.O (g31316), .I1 (g29609), .I2 (g29624));
OR2X1 gate16569(.O (g33316), .I1 (g29685), .I2 (g32178));
OR2X1 gate16570(.O (g22634), .I1 (g18934), .I2 (g15590));
OR2X1 gate16571(.O (g24207), .I1 (g23396), .I2 (g18119));
OR2X1 gate16572(.O (g22872), .I1 (g19372), .I2 (g19383));
OR4X1 gate16573(.O (I29985), .I1 (g29385), .I2 (g31376), .I3 (g30735), .I4 (g30825));
OR3X1 gate16574(.O (I22958), .I1 (g21603), .I2 (g21386), .I3 (g21365));
OR2X1 gate16575(.O (g34231), .I1 (g33898), .I2 (g33902));
OR2X1 gate16576(.O (g29504), .I1 (g28143), .I2 (g25875));
OR2X1 gate16577(.O (g25706), .I1 (g25030), .I2 (g18748));
OR2X1 gate16578(.O (g25597), .I1 (g24892), .I2 (g21719));
OR2X1 gate16579(.O (g32037), .I1 (g30566), .I2 (g29329));
OR2X1 gate16580(.O (g33989), .I1 (g33870), .I2 (g18398));
OR2X1 gate16581(.O (g33056), .I1 (g32327), .I2 (g22004));
OR2X1 gate16582(.O (g13570), .I1 (g9223), .I2 (g11130));
OR2X1 gate16583(.O (g25689), .I1 (g24849), .I2 (g21888));
OR2X1 gate16584(.O (g13914), .I1 (g8643), .I2 (g11380));
OR2X1 gate16585(.O (g33611), .I1 (g33243), .I2 (g18632));
OR2X1 gate16586(.O (g31924), .I1 (g31486), .I2 (g22049));
OR2X1 gate16587(.O (g32984), .I1 (g31934), .I2 (g18264));
OR2X1 gate16588(.O (g33988), .I1 (g33861), .I2 (g18397));
OR2X1 gate16589(.O (g25688), .I1 (g24812), .I2 (g21887));
OR2X1 gate16590(.O (g28750), .I1 (g27525), .I2 (g16765));
OR2X1 gate16591(.O (g25624), .I1 (g24408), .I2 (g18224));
OR2X1 gate16592(.O (g26916), .I1 (g25916), .I2 (g18232));
OR2X1 gate16593(.O (g30511), .I1 (g30180), .I2 (g22032));
OR2X1 gate16594(.O (g20241), .I1 (g16233), .I2 (g13541));
OR2X1 gate16595(.O (g32352), .I1 (g29852), .I2 (g31282));
OR4X1 gate16596(.O (I30746), .I1 (g32047), .I2 (g31985), .I3 (g31991), .I4 (g32309));
OR2X1 gate16597(.O (g24241), .I1 (g22920), .I2 (g18252));
OR2X1 gate16598(.O (g33271), .I1 (g32120), .I2 (g29549));
OR2X1 gate16599(.O (g27972), .I1 (g26131), .I2 (g26105));
OR2X1 gate16600(.O (g32155), .I1 (g30935), .I2 (g29475));
OR2X1 gate16601(.O (g15017), .I1 (g10776), .I2 (g8703));
OR2X1 gate16602(.O (g28091), .I1 (g27665), .I2 (g21913));
OR2X1 gate16603(.O (g32266), .I1 (g30604), .I2 (g29354));
OR2X1 gate16604(.O (g29245), .I1 (g28676), .I2 (g18384));
OR2X1 gate16605(.O (g26721), .I1 (g10776), .I2 (g24444));
OR2X1 gate16606(.O (g29299), .I1 (g28587), .I2 (g18794));
OR2X1 gate16607(.O (g33031), .I1 (g32315), .I2 (g21841));
OR2X1 gate16608(.O (g30456), .I1 (g29378), .I2 (g21869));
OR2X1 gate16609(.O (g34456), .I1 (g34395), .I2 (g18669));
OR2X1 gate16610(.O (g29298), .I1 (g28571), .I2 (g18793));
OR2X1 gate16611(.O (g24235), .I1 (g22632), .I2 (g18238));
OR2X1 gate16612(.O (g13941), .I1 (g11019), .I2 (g11023));
OR2X1 gate16613(.O (g31887), .I1 (g31292), .I2 (g21820));
OR2X1 gate16614(.O (g28390), .I1 (g27207), .I2 (g15861));
OR2X1 gate16615(.O (g30480), .I1 (g29321), .I2 (g21972));
OR2X1 gate16616(.O (g30916), .I1 (g13853), .I2 (g29799));
OR2X1 gate16617(.O (g29775), .I1 (g25966), .I2 (g28232));
OR4X1 gate16618(.O (I26523), .I1 (g20720), .I2 (g20857), .I3 (g20998), .I4 (g21143));
OR2X1 gate16619(.O (g25885), .I1 (g25522), .I2 (g23957));
OR2X1 gate16620(.O (g30550), .I1 (g30226), .I2 (g22121));
OR2X1 gate16621(.O (g30314), .I1 (g28268), .I2 (g27266));
OR2X1 gate16622(.O (g23615), .I1 (g20109), .I2 (g20131));
OR2X1 gate16623(.O (g30287), .I1 (g28653), .I2 (g27677));
OR2X1 gate16624(.O (g34314), .I1 (g25831), .I2 (g34061));
OR2X1 gate16625(.O (g30307), .I1 (g28256), .I2 (g27260));
OR2X1 gate16626(.O (g33393), .I1 (g32286), .I2 (g29984));
OR2X1 gate16627(.O (g23720), .I1 (g20165), .I2 (g16801));
OR4X1 gate16628(.O (I12902), .I1 (g4235), .I2 (g4232), .I3 (g4229), .I4 (g4226));
OR2X1 gate16629(.O (g25763), .I1 (g25113), .I2 (g18817));
OR2X1 gate16630(.O (g29232), .I1 (g28183), .I2 (g18231));
OR2X1 gate16631(.O (g31764), .I1 (g30015), .I2 (g30032));
OR2X1 gate16632(.O (g23275), .I1 (g19680), .I2 (g16160));
OR2X1 gate16633(.O (g34721), .I1 (g34696), .I2 (g18135));
OR2X1 gate16634(.O (g31869), .I1 (g30592), .I2 (g18221));
OR4X1 gate16635(.O (I30193), .I1 (g31070), .I2 (g30614), .I3 (g30673), .I4 (g31528));
OR2X1 gate16636(.O (g30431), .I1 (g29875), .I2 (g21815));
OR2X1 gate16637(.O (g33960), .I1 (g33759), .I2 (g21701));
OR2X1 gate16638(.O (g25660), .I1 (g24726), .I2 (g21785));
OR2X1 gate16639(.O (g29261), .I1 (g28247), .I2 (g18605));
OR2X1 gate16640(.O (g31868), .I1 (g30600), .I2 (g18204));
OR2X1 gate16641(.O (g26335), .I1 (g1526), .I2 (g24609));
OR2X1 gate16642(.O (g19572), .I1 (g17133), .I2 (g14193));
OR2X1 gate16643(.O (g22152), .I1 (g21188), .I2 (g17469));
OR2X1 gate16644(.O (g26930), .I1 (g26799), .I2 (g18544));
OR2X1 gate16645(.O (g34269), .I1 (g34083), .I2 (g18732));
OR2X1 gate16646(.O (g30341), .I1 (g29380), .I2 (g18246));
OR2X1 gate16647(.O (g26694), .I1 (g24444), .I2 (g10704));
OR2X1 gate16648(.O (g26965), .I1 (g26336), .I2 (g24317));
OR2X1 gate16649(.O (g33709), .I1 (g32414), .I2 (g33441));
OR2X1 gate16650(.O (g34268), .I1 (g34082), .I2 (g18730));
OR2X1 gate16651(.O (g31259), .I1 (g25992), .I2 (g29554));
OR2X1 gate16652(.O (g32285), .I1 (g31222), .I2 (g29740));
OR2X1 gate16653(.O (g33259), .I1 (g32109), .I2 (g29521));
OR2X1 gate16654(.O (g28536), .I1 (g27293), .I2 (g26205));
OR4X1 gate16655(.O (I30727), .I1 (g31759), .I2 (g32196), .I3 (g31933), .I4 (g31941));
OR2X1 gate16656(.O (g31258), .I1 (g25991), .I2 (g29550));
OR2X1 gate16657(.O (g24206), .I1 (g23386), .I2 (g18110));
OR2X1 gate16658(.O (g13728), .I1 (g6804), .I2 (g12527));
OR2X1 gate16659(.O (g28702), .I1 (g27457), .I2 (g16670));
OR2X1 gate16660(.O (g30734), .I1 (g13808), .I2 (g29774));
OR3X1 gate16661(.O (I22298), .I1 (g20371), .I2 (g20161), .I3 (g20151));
OR2X1 gate16662(.O (g30335), .I1 (g29746), .I2 (g18174));
OR2X1 gate16663(.O (g34734), .I1 (g34681), .I2 (g18652));
OR2X1 gate16664(.O (g25721), .I1 (g25057), .I2 (g18766));
OR2X1 gate16665(.O (g28621), .I1 (g27359), .I2 (g16518));
OR2X1 gate16666(.O (g25596), .I1 (g24865), .I2 (g21718));
OR4X1 gate16667(.O (I31853), .I1 (g33488), .I2 (g33489), .I3 (g33490), .I4 (g33491));
OR2X1 gate16668(.O (g33043), .I1 (g32195), .I2 (g24325));
OR2X1 gate16669(.O (g31244), .I1 (g25963), .I2 (g29515));
OR2X1 gate16670(.O (g20082), .I1 (g16026), .I2 (g13321));
OR2X1 gate16671(.O (g28564), .I1 (g27314), .I2 (g26252));
OR2X1 gate16672(.O (g23193), .I1 (g19556), .I2 (g15937));
OR4X1 gate16673(.O (I23756), .I1 (g23457), .I2 (g23480), .I3 (g23494), .I4 (g23511));
OR2X1 gate16674(.O (g26278), .I1 (g24545), .I2 (g24549));
OR2X1 gate16675(.O (g33069), .I1 (g32009), .I2 (g22113));
OR2X1 gate16676(.O (g33602), .I1 (g33425), .I2 (g18511));
OR2X1 gate16677(.O (g25942), .I1 (g24422), .I2 (g22298));
OR2X1 gate16678(.O (g31774), .I1 (g30046), .I2 (g30057));
OR2X1 gate16679(.O (g7834), .I1 (g2886), .I2 (g2946));
OR2X1 gate16680(.O (g30487), .I1 (g30187), .I2 (g21983));
OR2X1 gate16681(.O (g31375), .I1 (g29628), .I2 (g28339));
OR2X1 gate16682(.O (g33068), .I1 (g31994), .I2 (g22112));
OR3X1 gate16683(.O (g33955), .I1 (g33505), .I2 (I31858), .I3 (I31859));
OR2X1 gate16684(.O (g24345), .I1 (g23606), .I2 (g18788));
OR2X1 gate16685(.O (g25655), .I1 (g24645), .I2 (g18607));
OR2X1 gate16686(.O (g31879), .I1 (g31475), .I2 (g21745));
OR2X1 gate16687(.O (g30502), .I1 (g30232), .I2 (g22023));
OR2X1 gate16688(.O (g28062), .I1 (g27288), .I2 (g21746));
OR2X1 gate16689(.O (g30557), .I1 (g30247), .I2 (g22128));
OR2X1 gate16690(.O (g33970), .I1 (g33868), .I2 (g18322));
OR2X1 gate16691(.O (g34619), .I1 (g34528), .I2 (g18581));
OR3X1 gate16692(.O (I22880), .I1 (g21509), .I2 (g21356), .I3 (g21351));
OR2X1 gate16693(.O (g25670), .I1 (g24967), .I2 (g18626));
OR2X1 gate16694(.O (g29271), .I1 (g28333), .I2 (g18637));
OR2X1 gate16695(.O (g31878), .I1 (g31015), .I2 (g21733));
OR4X1 gate16696(.O (I31864), .I1 (g33510), .I2 (g33511), .I3 (g33512), .I4 (g33513));
OR2X1 gate16697(.O (g30443), .I1 (g29808), .I2 (g21852));
OR2X1 gate16698(.O (g34618), .I1 (g34527), .I2 (g18580));
OR2X1 gate16699(.O (g24398), .I1 (g23801), .I2 (g21296));
OR2X1 gate16700(.O (g30279), .I1 (g28637), .I2 (g27668));
OR2X1 gate16701(.O (g34443), .I1 (g34385), .I2 (g18545));
OR2X1 gate16702(.O (g25734), .I1 (g25058), .I2 (g18782));
OR2X1 gate16703(.O (g28634), .I1 (g27374), .I2 (g16536));
OR2X1 gate16704(.O (g28851), .I1 (g27558), .I2 (g16870));
OR2X1 gate16705(.O (g31886), .I1 (g31481), .I2 (g21791));
OR2X1 gate16706(.O (g29753), .I1 (g28213), .I2 (g22720));
OR4X1 gate16707(.O (g25839), .I1 (g25507), .I2 (g25485), .I3 (g25459), .I4 (g25420));
OR2X1 gate16708(.O (g34278), .I1 (g26829), .I2 (g34212));
OR2X1 gate16709(.O (g30469), .I1 (g30153), .I2 (g21940));
OR2X1 gate16710(.O (g33967), .I1 (g33842), .I2 (g18319));
OR2X1 gate16711(.O (g33994), .I1 (g33841), .I2 (g18424));
OR2X1 gate16712(.O (g27506), .I1 (g26021), .I2 (g24639));
OR2X1 gate16713(.O (g30286), .I1 (g28191), .I2 (g28186));
OR2X1 gate16714(.O (g25694), .I1 (g24638), .I2 (g18738));
OR2X1 gate16715(.O (g25667), .I1 (g24682), .I2 (g18619));
OR2X1 gate16716(.O (g24263), .I1 (g23497), .I2 (g18529));
OR2X1 gate16717(.O (g34286), .I1 (g26842), .I2 (g34216));
OR2X1 gate16718(.O (g30468), .I1 (g30238), .I2 (g21939));
OR2X1 gate16719(.O (g34468), .I1 (g34342), .I2 (g18718));
OR2X1 gate16720(.O (g34039), .I1 (g33743), .I2 (g18736));
OR2X1 gate16721(.O (g34306), .I1 (g25782), .I2 (g34054));
OR4X1 gate16722(.O (g29529), .I1 (g28303), .I2 (g28293), .I3 (g28283), .I4 (g28267));
OR2X1 gate16723(.O (g22640), .I1 (g18951), .I2 (g15613));
OR2X1 gate16724(.O (g34038), .I1 (g33731), .I2 (g18735));
OR2X1 gate16725(.O (g31919), .I1 (g31758), .I2 (g22044));
OR2X1 gate16726(.O (g32454), .I1 (g30322), .I2 (g31795));
OR2X1 gate16727(.O (g25619), .I1 (g24961), .I2 (g18193));
OR2X1 gate16728(.O (g15124), .I1 (g13605), .I2 (g4581));
OR2X1 gate16729(.O (g26884), .I1 (g26511), .I2 (g24190));
OR2X1 gate16730(.O (g28574), .I1 (g27324), .I2 (g26270));
OR2X1 gate16731(.O (g31918), .I1 (g31786), .I2 (g22015));
OR2X1 gate16732(.O (g28047), .I1 (g27676), .I2 (g18160));
OR2X1 gate16733(.O (g33010), .I1 (g32301), .I2 (g18473));
OR2X1 gate16734(.O (g34601), .I1 (g34488), .I2 (g18211));
OR2X1 gate16735(.O (g29764), .I1 (g28219), .I2 (g28226));
OR2X1 gate16736(.O (g25618), .I1 (g25491), .I2 (g18192));
OR2X1 gate16737(.O (g34975), .I1 (g34871), .I2 (g34964));
OR2X1 gate16738(.O (g24500), .I1 (g24011), .I2 (g21605));
OR2X1 gate16739(.O (g33545), .I1 (g33399), .I2 (g18324));
OR2X1 gate16740(.O (g9013), .I1 (g2472), .I2 (g2491));
OR2X1 gate16741(.O (g26363), .I1 (g2965), .I2 (g24965));
OR2X1 gate16742(.O (g33599), .I1 (g33087), .I2 (g18500));
OR2X1 gate16743(.O (g32239), .I1 (g30595), .I2 (g29350));
OR2X1 gate16744(.O (g28051), .I1 (g27699), .I2 (g18166));
OR2X1 gate16745(.O (g27240), .I1 (g25883), .I2 (g24467));
OR2X1 gate16746(.O (g28072), .I1 (g27086), .I2 (g21874));
OR2X1 gate16747(.O (g33598), .I1 (g33364), .I2 (g18496));
OR2X1 gate16748(.O (g32238), .I1 (g30594), .I2 (g29349));
OR4X1 gate16749(.O (I29352), .I1 (g29322), .I2 (g29315), .I3 (g30315), .I4 (g30308));
OR2X1 gate16750(.O (g28592), .I1 (g27333), .I2 (g26288));
OR4X1 gate16751(.O (I31874), .I1 (g33528), .I2 (g33529), .I3 (g33530), .I4 (g33531));
OR2X1 gate16752(.O (g34791), .I1 (g34771), .I2 (g18184));
OR2X1 gate16753(.O (g22662), .I1 (g19069), .I2 (g15679));
OR2X1 gate16754(.O (g34884), .I1 (g34858), .I2 (g21666));
OR2X1 gate16755(.O (g29259), .I1 (g28304), .I2 (g18603));
OR2X1 gate16756(.O (g29225), .I1 (g28451), .I2 (g18158));
OR2X1 gate16757(.O (g30410), .I1 (g29857), .I2 (g21769));
OR2X1 gate16758(.O (g31322), .I1 (g26128), .I2 (g29635));
OR2X1 gate16759(.O (g14062), .I1 (g11047), .I2 (g11116));
OR2X1 gate16760(.O (g34168), .I1 (g33787), .I2 (g19784));
OR2X1 gate16761(.O (g27563), .I1 (g26104), .I2 (g24704));
OR2X1 gate16762(.O (g29258), .I1 (g28238), .I2 (g18601));
OR2X1 gate16763(.O (g31901), .I1 (g31516), .I2 (g21909));
OR2X1 gate16764(.O (g33159), .I1 (g32016), .I2 (g30730));
OR2X1 gate16765(.O (g30479), .I1 (g29320), .I2 (g21950));
OR2X1 gate16766(.O (g33977), .I1 (g33876), .I2 (g18348));
OR2X1 gate16767(.O (g30363), .I1 (g30121), .I2 (g18407));
OR2X1 gate16768(.O (g25601), .I1 (g24660), .I2 (g18112));
OR2X1 gate16769(.O (g12981), .I1 (g12219), .I2 (g9967));
OR2X1 gate16770(.O (g24273), .I1 (g23166), .I2 (g18630));
OR2X1 gate16771(.O (g25677), .I1 (g24684), .I2 (g21834));
OR2X1 gate16772(.O (g31783), .I1 (I29351), .I2 (I29352));
OR2X1 gate16773(.O (g23209), .I1 (g19585), .I2 (g19601));
OR2X1 gate16774(.O (g30478), .I1 (g30248), .I2 (g21949));
OR2X1 gate16775(.O (g34015), .I1 (g33858), .I2 (g18502));
OR2X1 gate16776(.O (g29244), .I1 (g28692), .I2 (g18380));
OR2X1 gate16777(.O (g33561), .I1 (g33408), .I2 (g18376));
OR2X1 gate16778(.O (g30486), .I1 (g30177), .I2 (g21982));
OR2X1 gate16779(.O (g31295), .I1 (g26090), .I2 (g29598));
OR2X1 gate16780(.O (g26922), .I1 (g25902), .I2 (g18288));
OR2X1 gate16781(.O (g28731), .I1 (g27504), .I2 (g16733));
OR2X1 gate16782(.O (g33295), .I1 (g32153), .I2 (g29605));
OR2X1 gate16783(.O (g31144), .I1 (g29477), .I2 (g28193));
OR2X1 gate16784(.O (g25937), .I1 (g24406), .I2 (g22216));
OR2X1 gate16785(.O (g30556), .I1 (g30236), .I2 (g22127));
OR2X1 gate16786(.O (g24234), .I1 (g22622), .I2 (g18237));
OR2X1 gate16787(.O (g13973), .I1 (g11024), .I2 (g11028));
OR2X1 gate16788(.O (g29068), .I1 (g27628), .I2 (g17119));
OR4X1 gate16789(.O (g25791), .I1 (g25411), .I2 (g25371), .I3 (g25328), .I4 (g25290));
OR2X1 gate16790(.O (g28691), .I1 (g27437), .I2 (g16642));
OR2X1 gate16791(.O (g29879), .I1 (g28289), .I2 (g26096));
OR2X1 gate16792(.O (g26953), .I1 (g26486), .I2 (g24291));
OR2X1 gate16793(.O (g28405), .I1 (g27216), .I2 (g15875));
OR2X1 gate16794(.O (g33966), .I1 (g33837), .I2 (g18318));
OR2X1 gate16795(.O (g25666), .I1 (g24788), .I2 (g21793));
OR2X1 gate16796(.O (g33017), .I1 (g32292), .I2 (g18510));
OR2X1 gate16797(.O (g26800), .I1 (g24922), .I2 (g24929));
OR2X1 gate16798(.O (g34321), .I1 (g25866), .I2 (g34065));
OR2X1 gate16799(.O (g30531), .I1 (g30274), .I2 (g22077));
OR2X1 gate16800(.O (g23346), .I1 (g19736), .I2 (g16204));
OR2X1 gate16801(.O (g29792), .I1 (g28235), .I2 (g28244));
OR2X1 gate16802(.O (g12832), .I1 (g10347), .I2 (g10348));
OR2X1 gate16803(.O (g13761), .I1 (g490), .I2 (g12527));
OR2X1 gate16804(.O (g16022), .I1 (g13048), .I2 (g10707));
OR2X1 gate16805(.O (g26334), .I1 (g1171), .I2 (g24591));
OR2X1 gate16806(.O (g28046), .I1 (g27667), .I2 (g18157));
OR2X1 gate16807(.O (g32349), .I1 (g29840), .I2 (g31275));
OR2X1 gate16808(.O (g31289), .I1 (g29580), .I2 (g29591));
OR2X1 gate16809(.O (g30373), .I1 (g30111), .I2 (g18461));
OR2X1 gate16810(.O (g33289), .I1 (g32148), .I2 (g29588));
OR2X1 gate16811(.O (g22331), .I1 (g21405), .I2 (g17809));
OR2X1 gate16812(.O (g26964), .I1 (g26259), .I2 (g24316));
OR2X1 gate16813(.O (g34373), .I1 (g26292), .I2 (g34138));
OR2X1 gate16814(.O (g33023), .I1 (g32313), .I2 (g21751));
OR2X1 gate16815(.O (g31288), .I1 (g2955), .I2 (g29914));
OR2X1 gate16816(.O (g23153), .I1 (g19521), .I2 (g15876));
OR2X1 gate16817(.O (g33288), .I1 (g32147), .I2 (g29587));
OR2X1 gate16818(.O (g31308), .I1 (g26101), .I2 (g29614));
OR2X1 gate16819(.O (g33571), .I1 (g33367), .I2 (g18409));
OR2X1 gate16820(.O (g30417), .I1 (g29874), .I2 (g21801));
OR2X1 gate16821(.O (g34800), .I1 (g34752), .I2 (g18586));
OR2X1 gate16822(.O (g34417), .I1 (g27678), .I2 (g34196));
OR2X1 gate16823(.O (g28357), .I1 (g27148), .I2 (g15836));
OR2X1 gate16824(.O (g30334), .I1 (g29837), .I2 (g18143));
OR2X1 gate16825(.O (g28105), .I1 (g27997), .I2 (g22135));
OR2X1 gate16826(.O (g28743), .I1 (g27517), .I2 (g16758));
OR2X1 gate16827(.O (g29078), .I1 (g27633), .I2 (g26572));
OR2X1 gate16828(.O (g26909), .I1 (g26543), .I2 (g24227));
OR3X1 gate16829(.O (I18385), .I1 (g14413), .I2 (g14391), .I3 (g14360));
OR2X1 gate16830(.O (g34762), .I1 (g34687), .I2 (g34524));
OR2X1 gate16831(.O (g25740), .I1 (g25164), .I2 (g22055));
OR2X1 gate16832(.O (g26908), .I1 (g26358), .I2 (g24225));
OR2X1 gate16833(.O (g28640), .I1 (g27384), .I2 (g16590));
OR2X1 gate16834(.O (g30423), .I1 (g29887), .I2 (g21807));
OR2X1 gate16835(.O (g33976), .I1 (g33869), .I2 (g18347));
OR2X1 gate16836(.O (g33985), .I1 (g33896), .I2 (g18382));
OR3X1 gate16837(.O (g24946), .I1 (g22360), .I2 (g22409), .I3 (g8130));
OR2X1 gate16838(.O (g25676), .I1 (g24668), .I2 (g21833));
OR2X1 gate16839(.O (g25685), .I1 (g24476), .I2 (g21866));
OR4X1 gate16840(.O (I30750), .I1 (g31788), .I2 (g32310), .I3 (g32054), .I4 (g32070));
OR3X1 gate16841(.O (g33954), .I1 (g33496), .I2 (I31853), .I3 (I31854));
OR2X1 gate16842(.O (g21891), .I1 (g19948), .I2 (g15103));
OR2X1 gate16843(.O (g24344), .I1 (g22145), .I2 (g18787));
OR2X1 gate16844(.O (g25654), .I1 (g24634), .I2 (g18606));
OR2X1 gate16845(.O (g25936), .I1 (g24403), .I2 (g22209));
OR2X1 gate16846(.O (g30543), .I1 (g29338), .I2 (g22110));
OR4X1 gate16847(.O (I26522), .I1 (g19890), .I2 (g19935), .I3 (g19984), .I4 (g26365));
OR2X1 gate16848(.O (g31260), .I1 (g25993), .I2 (g29555));
OR2X1 gate16849(.O (g34000), .I1 (g33943), .I2 (g18441));
OR2X1 gate16850(.O (g26751), .I1 (g24903), .I2 (g24912));
OR2X1 gate16851(.O (g33260), .I1 (g32110), .I2 (g29524));
OR2X1 gate16852(.O (g29295), .I1 (g28663), .I2 (g18780));
OR2X1 gate16853(.O (g31668), .I1 (g29924), .I2 (g28558));
OR2X1 gate16854(.O (g14583), .I1 (g10685), .I2 (g542));
OR2X1 gate16855(.O (g25762), .I1 (g25095), .I2 (g18816));
OR2X1 gate16856(.O (g28662), .I1 (g27407), .I2 (g16612));
OR2X1 gate16857(.O (g26293), .I1 (g24550), .I2 (g24555));
OR2X1 gate16858(.O (g33559), .I1 (g33073), .I2 (g18368));
OR4X1 gate16859(.O (I30192), .I1 (g29385), .I2 (g31376), .I3 (g30735), .I4 (g30825));
OR2X1 gate16860(.O (g33016), .I1 (g32284), .I2 (g18509));
OR2X1 gate16861(.O (g25587), .I1 (g21682), .I2 (g24157));
OR2X1 gate16862(.O (g33558), .I1 (g33350), .I2 (g18364));
OR2X1 gate16863(.O (g23750), .I1 (g20174), .I2 (g16840));
OR2X1 gate16864(.O (g31893), .I1 (g31490), .I2 (g21837));
OR2X1 gate16865(.O (g34807), .I1 (g34764), .I2 (g18596));
OR2X1 gate16866(.O (g34974), .I1 (g34870), .I2 (g34963));
OR2X1 gate16867(.O (g31865), .I1 (g31149), .I2 (g21709));
OR2X1 gate16868(.O (g33544), .I1 (g33392), .I2 (g18317));
OR2X1 gate16869(.O (g34639), .I1 (g34486), .I2 (g18722));
OR2X1 gate16870(.O (g12911), .I1 (g10278), .I2 (g12768));
OR2X1 gate16871(.O (g30293), .I1 (g28236), .I2 (g27246));
OR3X1 gate16872(.O (g23796), .I1 (g21462), .I2 (g21433), .I3 (I22958));
OR2X1 gate16873(.O (g28778), .I1 (g27540), .I2 (g16808));
OR2X1 gate16874(.O (g16239), .I1 (g7892), .I2 (g13432));
OR2X1 gate16875(.O (g34293), .I1 (g26854), .I2 (g34224));
OR2X1 gate16876(.O (g34638), .I1 (g34484), .I2 (g18721));
OR2X1 gate16877(.O (g34265), .I1 (g34117), .I2 (g18711));
OR2X1 gate16878(.O (g30416), .I1 (g29858), .I2 (g21800));
OR2X1 gate16879(.O (g27591), .I1 (g26181), .I2 (g24765));
OR2X1 gate16880(.O (g34416), .I1 (g34191), .I2 (g25159));
OR2X1 gate16881(.O (g29289), .I1 (g28642), .I2 (g18763));
OR2X1 gate16882(.O (g25747), .I1 (g25130), .I2 (g18795));
OR2X1 gate16883(.O (g28647), .I1 (g27389), .I2 (g16596));
OR2X1 gate16884(.O (g33610), .I1 (g33242), .I2 (g18616));
OR2X1 gate16885(.O (g29309), .I1 (g28722), .I2 (g18818));
OR2X1 gate16886(.O (g30391), .I1 (g30080), .I2 (g18557));
OR2X1 gate16887(.O (g33042), .I1 (g32193), .I2 (g24324));
OR2X1 gate16888(.O (g27147), .I1 (g25802), .I2 (g24399));
OR2X1 gate16889(.O (g31255), .I1 (g25982), .I2 (g29536));
OR2X1 gate16890(.O (g29288), .I1 (g28630), .I2 (g18762));
OR2X1 gate16891(.O (g33255), .I1 (g32106), .I2 (g29514));
OR2X1 gate16892(.O (g29224), .I1 (g28919), .I2 (g18156));
OR2X1 gate16893(.O (g30510), .I1 (g30263), .I2 (g22031));
OR2X1 gate16894(.O (g29308), .I1 (g28612), .I2 (g18815));
OR2X1 gate16895(.O (g24240), .I1 (g22861), .I2 (g18251));
OR2X1 gate16896(.O (g33270), .I1 (g32119), .I2 (g29547));
OR2X1 gate16897(.O (g28090), .I1 (g27275), .I2 (g18733));
OR2X1 gate16898(.O (g30579), .I1 (g30173), .I2 (g14571));
OR2X1 gate16899(.O (g27858), .I1 (g17405), .I2 (g26737));
OR2X1 gate16900(.O (g25751), .I1 (g25061), .I2 (g22098));
OR2X1 gate16901(.O (g28651), .I1 (g27392), .I2 (g16599));
OR2X1 gate16902(.O (g29495), .I1 (g28563), .I2 (g27614));
OR2X1 gate16903(.O (g33383), .I1 (g32244), .I2 (g29940));
OR2X1 gate16904(.O (g25639), .I1 (g25122), .I2 (g18530));
OR2X1 gate16905(.O (g34014), .I1 (g33647), .I2 (g18493));
OR2X1 gate16906(.O (g33030), .I1 (g32166), .I2 (g21826));
OR2X1 gate16907(.O (g31267), .I1 (g29548), .I2 (g28263));
OR2X1 gate16908(.O (g25638), .I1 (g24977), .I2 (g18316));
OR2X1 gate16909(.O (g34007), .I1 (g33640), .I2 (g18467));
OR2X1 gate16910(.O (g16883), .I1 (g13509), .I2 (g11115));
OR2X1 gate16911(.O (g33267), .I1 (g32115), .I2 (g29535));
OR2X1 gate16912(.O (g33294), .I1 (g32152), .I2 (g29604));
OR2X1 gate16913(.O (g27394), .I1 (g25957), .I2 (g24573));
OR2X1 gate16914(.O (g28331), .I1 (g27129), .I2 (g15814));
OR2X1 gate16915(.O (g30442), .I1 (g29797), .I2 (g21851));
OR2X1 gate16916(.O (g33065), .I1 (g32008), .I2 (g22068));
OR2X1 gate16917(.O (g34442), .I1 (g34380), .I2 (g18542));
OR2X1 gate16918(.O (g28513), .I1 (g27276), .I2 (g26123));
OR2X1 gate16919(.O (g31875), .I1 (g31066), .I2 (g21730));
OR2X1 gate16920(.O (g29643), .I1 (g28192), .I2 (g27145));
OR2X1 gate16921(.O (g34615), .I1 (g34516), .I2 (g18576));
OR3X1 gate16922(.O (g33219), .I1 (g32335), .I2 (I30760), .I3 (I30761));
OR2X1 gate16923(.O (g24262), .I1 (g23387), .I2 (g18315));
OR2X1 gate16924(.O (g28404), .I1 (g27215), .I2 (g15874));
OR2X1 gate16925(.O (g34720), .I1 (g34694), .I2 (g18134));
OR2X1 gate16926(.O (g34041), .I1 (g33829), .I2 (g18739));
OR2X1 gate16927(.O (g28717), .I1 (g27482), .I2 (g16701));
OR2X1 gate16928(.O (g30430), .I1 (g29859), .I2 (g21814));
OR2X1 gate16929(.O (g30493), .I1 (g30198), .I2 (g21989));
OR2X1 gate16930(.O (g28212), .I1 (g27030), .I2 (g27035));
OR2X1 gate16931(.O (g29260), .I1 (g28315), .I2 (g18604));
OR2X1 gate16932(.O (g25835), .I1 (g25367), .I2 (g23855));
OR2X1 gate16933(.O (g30465), .I1 (g30164), .I2 (g21936));
OR2X1 gate16934(.O (g34465), .I1 (g34295), .I2 (g18712));
OR2X1 gate16935(.O (g25586), .I1 (g21678), .I2 (g24156));
OR2X1 gate16936(.O (g34237), .I1 (g32715), .I2 (g33955));
OR2X1 gate16937(.O (g30340), .I1 (g29377), .I2 (g18245));
OR2X1 gate16938(.O (g29489), .I1 (g28550), .I2 (g27601));
OR2X1 gate16939(.O (g34035), .I1 (g33721), .I2 (g18714));
OR2X1 gate16940(.O (g29488), .I1 (g28547), .I2 (g27600));
OR2X1 gate16941(.O (g34806), .I1 (g34763), .I2 (g18595));
OR2X1 gate16942(.O (g23183), .I1 (g19545), .I2 (g15911));
OR2X1 gate16943(.O (g28723), .I1 (g27490), .I2 (g16706));
OR2X1 gate16944(.O (g33617), .I1 (g33263), .I2 (g24326));
OR2X1 gate16945(.O (g31915), .I1 (g31520), .I2 (g22001));
OR2X1 gate16946(.O (g25615), .I1 (g24803), .I2 (g18162));
OR2X1 gate16947(.O (g30517), .I1 (g30244), .I2 (g22038));
OR2X1 gate16948(.O (g28387), .I1 (g27203), .I2 (g15858));
OR2X1 gate16949(.O (g31277), .I1 (g29570), .I2 (g28285));
OR2X1 gate16950(.O (g25720), .I1 (g25042), .I2 (g18765));
OR2X1 gate16951(.O (g24247), .I1 (g22623), .I2 (g18259));
OR2X1 gate16952(.O (g33277), .I1 (g32129), .I2 (g29568));
OR3X1 gate16953(.O (g14182), .I1 (g11741), .I2 (g11721), .I3 (g753));
OR2X1 gate16954(.O (g15935), .I1 (g13029), .I2 (g10665));
OR2X1 gate16955(.O (g28097), .I1 (g27682), .I2 (g22005));
OR2X1 gate16956(.O (g28104), .I1 (g27697), .I2 (g22108));
OR2X1 gate16957(.O (g25746), .I1 (g25217), .I2 (g22063));
OR2X1 gate16958(.O (g28646), .I1 (g27388), .I2 (g16595));
OR2X1 gate16959(.O (g33595), .I1 (g33368), .I2 (g18489));
OR2X1 gate16960(.O (g32235), .I1 (g31151), .I2 (g29662));
OR2X1 gate16961(.O (g27562), .I1 (g26102), .I2 (g24703));
OR2X1 gate16962(.O (g33623), .I1 (g33370), .I2 (g18792));
OR4X1 gate16963(.O (I30756), .I1 (g32088), .I2 (g32163), .I3 (g32098), .I4 (g32105));
OR2X1 gate16964(.O (g33037), .I1 (g32177), .I2 (g24310));
OR2X1 gate16965(.O (g30362), .I1 (g30120), .I2 (g18392));
OR2X1 gate16966(.O (g34193), .I1 (g33809), .I2 (g33814));
OR2X1 gate16967(.O (g24251), .I1 (g22637), .I2 (g18296));
OR2X1 gate16968(.O (g24272), .I1 (g23056), .I2 (g18629));
OR2X1 gate16969(.O (g31782), .I1 (g30060), .I2 (g30070));
OR2X1 gate16970(.O (g27290), .I1 (g25926), .I2 (g25928));
OR2X1 gate16971(.O (g28369), .I1 (g27160), .I2 (g25938));
OR2X1 gate16972(.O (g30523), .I1 (g30245), .I2 (g22069));
OR2X1 gate16973(.O (g33984), .I1 (g33881), .I2 (g18374));
OR2X1 gate16974(.O (g25684), .I1 (g24983), .I2 (g18643));
OR2X1 gate16975(.O (g29255), .I1 (g28714), .I2 (g18516));
OR2X1 gate16976(.O (g28368), .I1 (g27158), .I2 (g27184));
OR2X1 gate16977(.O (g26703), .I1 (g24447), .I2 (g10705));
OR2X1 gate16978(.O (g29270), .I1 (g28258), .I2 (g18635));
OR2X1 gate16979(.O (g32991), .I1 (g32322), .I2 (g18349));
OR2X1 gate16980(.O (g30475), .I1 (g30220), .I2 (g21946));
OR2X1 gate16981(.O (g34006), .I1 (g33897), .I2 (g18462));
OR2X1 gate16982(.O (g28850), .I1 (g27557), .I2 (g16869));
OR2X1 gate16983(.O (g33266), .I1 (g32114), .I2 (g29532));
OR2X1 gate16984(.O (g23574), .I1 (g20093), .I2 (g20108));
OR2X1 gate16985(.O (g13972), .I1 (g11232), .I2 (g11203));
OR2X1 gate16986(.O (g34727), .I1 (g34655), .I2 (g18213));
OR2X1 gate16987(.O (g26781), .I1 (g24913), .I2 (g24921));
OR2X1 gate16988(.O (g30437), .I1 (g29876), .I2 (g21846));
OR2X1 gate16989(.O (g26952), .I1 (g26360), .I2 (g24290));
OR2X1 gate16990(.O (g29294), .I1 (g28645), .I2 (g18779));
OR2X1 gate16991(.O (g29267), .I1 (g28257), .I2 (g18622));
OR2X1 gate16992(.O (g19619), .I1 (g15712), .I2 (g13080));
OR2X1 gate16993(.O (g8863), .I1 (g1644), .I2 (g1664));
OR2X1 gate16994(.O (g19557), .I1 (g17123), .I2 (g14190));
OR3X1 gate16995(.O (I22830), .I1 (g21429), .I2 (g21338), .I3 (g21307));
OR2X1 gate16996(.O (g27403), .I1 (g25962), .I2 (g24581));
OR2X1 gate16997(.O (g33589), .I1 (g33340), .I2 (g18469));
OR2X1 gate16998(.O (g30347), .I1 (g29383), .I2 (g18304));
OR2X1 gate16999(.O (g28716), .I1 (g27481), .I2 (g13887));
OR2X1 gate17000(.O (g34347), .I1 (g25986), .I2 (g34102));
OR2X1 gate17001(.O (g33588), .I1 (g33334), .I2 (g18468));
OR2X1 gate17002(.O (g34253), .I1 (g34171), .I2 (g24300));
OR2X1 gate17003(.O (g27226), .I1 (g25872), .I2 (g24436));
OR2X1 gate17004(.O (g28582), .I1 (g27330), .I2 (g26277));
OR2X1 gate17005(.O (g34600), .I1 (g34538), .I2 (g18182));
OR2X1 gate17006(.O (g24447), .I1 (g10948), .I2 (g22450));
OR2X1 gate17007(.O (g14387), .I1 (g9086), .I2 (g11048));
OR2X1 gate17008(.O (g34781), .I1 (g33431), .I2 (g34715));
OR2X1 gate17009(.O (g27551), .I1 (g26091), .I2 (g24675));
OR2X1 gate17010(.O (g27572), .I1 (g26129), .I2 (g24724));
OR2X1 gate17011(.O (g33119), .I1 (g32420), .I2 (g32428));
OR2X1 gate17012(.O (g28310), .I1 (g27107), .I2 (g15797));
OR2X1 gate17013(.O (g34236), .I1 (g32650), .I2 (g33954));
OR2X1 gate17014(.O (g30351), .I1 (g30084), .I2 (g18339));
OR2X1 gate17015(.O (g30372), .I1 (g30110), .I2 (g18446));
OR2X1 gate17016(.O (g25727), .I1 (g25163), .I2 (g22010));
OR2X1 gate17017(.O (g33118), .I1 (g32413), .I2 (g32418));
OR2X1 gate17018(.O (g34372), .I1 (g26287), .I2 (g34137));
OR2X1 gate17019(.O (g31864), .I1 (g31271), .I2 (g21703));
OR2X1 gate17020(.O (g33022), .I1 (g32306), .I2 (g21750));
OR2X1 gate17021(.O (g26422), .I1 (g24774), .I2 (g23104));
OR2X1 gate17022(.O (g31749), .I1 (g29974), .I2 (g29988));
OR2X1 gate17023(.O (g16052), .I1 (g13060), .I2 (g10724));
OR2X1 gate17024(.O (g7450), .I1 (g1277), .I2 (g1283));
OR2X1 gate17025(.O (g28050), .I1 (g27692), .I2 (g18165));
OR2X1 gate17026(.O (g33616), .I1 (g33237), .I2 (g24314));
OR2X1 gate17027(.O (g33313), .I1 (g29649), .I2 (g32171));
OR2X1 gate17028(.O (g30516), .I1 (g30233), .I2 (g22037));
OR2X1 gate17029(.O (g34264), .I1 (g34081), .I2 (g18701));
OR2X1 gate17030(.O (g28386), .I1 (g27202), .I2 (g13277));
OR2X1 gate17031(.O (g34790), .I1 (g34774), .I2 (g18151));
OR2X1 gate17032(.O (g31276), .I1 (g29567), .I2 (g28282));
OR2X1 gate17033(.O (g25703), .I1 (g25087), .I2 (g21922));
OR2X1 gate17034(.O (g28603), .I1 (g27340), .I2 (g26300));
OR2X1 gate17035(.O (g24246), .I1 (g23372), .I2 (g18257));
OR2X1 gate17036(.O (g33276), .I1 (g32128), .I2 (g29566));
OR2X1 gate17037(.O (g28096), .I1 (g27988), .I2 (g21997));
OR2X1 gate17038(.O (g32399), .I1 (g31527), .I2 (g30062));
OR2X1 gate17039(.O (g33053), .I1 (g31967), .I2 (g21974));
OR2X1 gate17040(.O (g31254), .I1 (g25981), .I2 (g29534));
OR2X1 gate17041(.O (g27980), .I1 (g26105), .I2 (g26131));
OR2X1 gate17042(.O (g33254), .I1 (g32104), .I2 (g29512));
OR2X1 gate17043(.O (g31900), .I1 (g31484), .I2 (g21908));
OR2X1 gate17044(.O (g31466), .I1 (g26160), .I2 (g29650));
OR2X1 gate17045(.O (g32398), .I1 (g31526), .I2 (g30061));
OR3X1 gate17046(.O (I22267), .I1 (g20236), .I2 (g20133), .I3 (g20111));
OR2X1 gate17047(.O (g25600), .I1 (g24650), .I2 (g18111));
OR2X1 gate17048(.O (g26913), .I1 (g25848), .I2 (g18225));
OR2X1 gate17049(.O (g28681), .I1 (g27428), .I2 (g16634));
OR2X1 gate17050(.O (g23405), .I1 (g19791), .I2 (g16245));
OR2X1 gate17051(.O (g29277), .I1 (g28440), .I2 (g18710));
OR2X1 gate17052(.O (g30422), .I1 (g29795), .I2 (g21806));
OR2X1 gate17053(.O (g33036), .I1 (g32168), .I2 (g24309));
OR2X1 gate17054(.O (g28429), .I1 (g27228), .I2 (g15913));
OR2X1 gate17055(.O (g33560), .I1 (g33404), .I2 (g18369));
OR2X1 gate17056(.O (g24355), .I1 (g23799), .I2 (g18824));
OR2X1 gate17057(.O (g28730), .I1 (g27503), .I2 (g13912));
OR2X1 gate17058(.O (g26905), .I1 (g26397), .I2 (g24222));
OR4X1 gate17059(.O (g25821), .I1 (g25482), .I2 (g25456), .I3 (g25417), .I4 (g25377));
OR2X1 gate17060(.O (g28428), .I1 (g27227), .I2 (g15912));
OR2X1 gate17061(.O (g30542), .I1 (g29337), .I2 (g22088));
OR2X1 gate17062(.O (g30453), .I1 (g29902), .I2 (g21862));
OR2X1 gate17063(.O (g33064), .I1 (g31993), .I2 (g22067));
OR2X1 gate17064(.O (g19363), .I1 (g17810), .I2 (g14913));
OR2X1 gate17065(.O (g28690), .I1 (g27436), .I2 (g16641));
OR2X1 gate17066(.O (g34021), .I1 (g33652), .I2 (g18519));
OR2X1 gate17067(.O (g34453), .I1 (g34410), .I2 (g18666));
OR2X1 gate17068(.O (g27426), .I1 (g25967), .I2 (g24588));
OR2X1 gate17069(.O (g28549), .I1 (g27304), .I2 (g26233));
OR2X1 gate17070(.O (g24151), .I1 (g18088), .I2 (g21661));
OR2X1 gate17071(.O (g33733), .I1 (g33105), .I2 (g32012));
OR2X1 gate17072(.O (g32361), .I1 (g29869), .I2 (g31300));
OR2X1 gate17073(.O (g34726), .I1 (g34665), .I2 (g18212));
OR2X1 gate17074(.O (g28548), .I1 (g27303), .I2 (g26232));
OR2X1 gate17075(.O (g31874), .I1 (g31016), .I2 (g21729));
OR2X1 gate17076(.O (g30436), .I1 (g29860), .I2 (g21845));
OR2X1 gate17077(.O (g19486), .I1 (g15589), .I2 (g12979));
OR2X1 gate17078(.O (g34614), .I1 (g34518), .I2 (g18568));
OR2X1 gate17079(.O (g29266), .I1 (g28330), .I2 (g18621));
OR2X1 gate17080(.O (g34607), .I1 (g34567), .I2 (g15081));
OR2X1 gate17081(.O (g30530), .I1 (g30224), .I2 (g22076));
OR2X1 gate17082(.O (g28317), .I1 (g27114), .I2 (g15805));
OR2X1 gate17083(.O (g33009), .I1 (g32273), .I2 (g18458));
OR2X1 gate17084(.O (g34274), .I1 (g27822), .I2 (g34205));
OR2X1 gate17085(.O (g30346), .I1 (g29381), .I2 (g18303));
OR2X1 gate17086(.O (g25834), .I1 (g25366), .I2 (g23854));
OR2X1 gate17087(.O (g27024), .I1 (g26826), .I2 (g17692));
OR4X1 gate17088(.O (I31849), .I1 (g33483), .I2 (g33484), .I3 (g33485), .I4 (g33486));
OR2X1 gate17089(.O (g33008), .I1 (g32261), .I2 (g18457));
OR2X1 gate17090(.O (g30464), .I1 (g30152), .I2 (g21935));
OR2X1 gate17091(.O (g32221), .I1 (g31140), .I2 (g29634));
OR2X1 gate17092(.O (g34464), .I1 (g34340), .I2 (g18687));
OR2X1 gate17093(.O (g31892), .I1 (g31019), .I2 (g21825));
OR4X1 gate17094(.O (I31848), .I1 (g33479), .I2 (g33480), .I3 (g33481), .I4 (g33482));
OR2X1 gate17095(.O (g28057), .I1 (g27033), .I2 (g18218));
OR2X1 gate17096(.O (g34034), .I1 (g33719), .I2 (g18713));
OR2X1 gate17097(.O (g33555), .I1 (g33355), .I2 (g18357));
OR2X1 gate17098(.O (g34641), .I1 (g34479), .I2 (g18724));
OR2X1 gate17099(.O (g34797), .I1 (g34747), .I2 (g18574));
OR2X1 gate17100(.O (g25726), .I1 (g25148), .I2 (g22009));
OR2X1 gate17101(.O (g33570), .I1 (g33420), .I2 (g18405));
OR2X1 gate17102(.O (g31914), .I1 (g31499), .I2 (g22000));
OR2X1 gate17103(.O (g34292), .I1 (g26853), .I2 (g34223));
OR2X1 gate17104(.O (g28323), .I1 (g27118), .I2 (g15810));
OR2X1 gate17105(.O (g33914), .I1 (g33305), .I2 (g33311));
OR2X1 gate17106(.O (g34153), .I1 (g33899), .I2 (g33451));
OR2X1 gate17107(.O (g27126), .I1 (g24378), .I2 (g25787));
OR2X1 gate17108(.O (g25614), .I1 (g24797), .I2 (g18161));
OR2X1 gate17109(.O (g28533), .I1 (g27291), .I2 (g26203));
OR2X1 gate17110(.O (g31907), .I1 (g31492), .I2 (g21954));
OR2X1 gate17111(.O (g30409), .I1 (g29842), .I2 (g21768));
OR2X1 gate17112(.O (g27250), .I1 (g25901), .I2 (g15738));
OR2X1 gate17113(.O (g26891), .I1 (g26652), .I2 (g24197));
OR2X1 gate17114(.O (g24203), .I1 (g22982), .I2 (g18107));
OR2X1 gate17115(.O (g25607), .I1 (g24773), .I2 (g18118));
OR2X1 gate17116(.O (g10802), .I1 (g7533), .I2 (g1296));
OR4X1 gate17117(.O (g15732), .I1 (g13411), .I2 (g13384), .I3 (g13349), .I4 (g11016));
OR2X1 gate17118(.O (g28775), .I1 (g27537), .I2 (g16806));
OR2X1 gate17119(.O (g30408), .I1 (g29806), .I2 (g21767));
OR2X1 gate17120(.O (g29864), .I1 (g28272), .I2 (g26086));
OR2X1 gate17121(.O (g34635), .I1 (g34485), .I2 (g18692));
OR2X1 gate17122(.O (g25593), .I1 (g24716), .I2 (g21707));
OR2X1 gate17123(.O (g33567), .I1 (g33081), .I2 (g18394));
OR2X1 gate17124(.O (g33594), .I1 (g33421), .I2 (g18485));
OR2X1 gate17125(.O (g32371), .I1 (g29883), .I2 (g31313));
OR2X1 gate17126(.O (g29313), .I1 (g28284), .I2 (g27270));
OR2X1 gate17127(.O (g24281), .I1 (g23397), .I2 (g18656));
OR2X1 gate17128(.O (g33238), .I1 (g32048), .I2 (g32051));
OR2X1 gate17129(.O (g26327), .I1 (g8462), .I2 (g24591));
OR2X1 gate17130(.O (g22225), .I1 (g21332), .I2 (g17654));
OR2X1 gate17131(.O (g29748), .I1 (g28210), .I2 (g28214));
OR2X1 gate17132(.O (g22708), .I1 (g19266), .I2 (g15711));
OR2X1 gate17133(.O (g29276), .I1 (g28616), .I2 (g18709));
OR2X1 gate17134(.O (g29285), .I1 (g28639), .I2 (g18750));
OR2X1 gate17135(.O (g29305), .I1 (g28602), .I2 (g18811));
OR2X1 gate17136(.O (g29254), .I1 (g28725), .I2 (g18512));
OR3X1 gate17137(.O (g33176), .I1 (g32198), .I2 (I30734), .I3 (I30735));
OR2X1 gate17138(.O (g16882), .I1 (g13508), .I2 (g11114));
OR2X1 gate17139(.O (g30474), .I1 (g30208), .I2 (g21945));
OR2X1 gate17140(.O (g25635), .I1 (g24504), .I2 (g18293));
OR2X1 gate17141(.O (g31883), .I1 (g31132), .I2 (g21777));
OR2X1 gate17142(.O (g30537), .I1 (g30246), .I2 (g22083));
OR2X1 gate17143(.O (g19587), .I1 (g15700), .I2 (g13046));
OR4X1 gate17144(.O (I30331), .I1 (g31672), .I2 (g31710), .I3 (g31021), .I4 (g30937));
OR2X1 gate17145(.O (g34537), .I1 (g34324), .I2 (g34084));
OR2X1 gate17146(.O (g13794), .I1 (g7396), .I2 (g10684));
OR2X1 gate17147(.O (g34283), .I1 (g26839), .I2 (g34215));
OR2X1 gate17148(.O (g30492), .I1 (g30188), .I2 (g21988));
OR2X1 gate17149(.O (g34606), .I1 (g34564), .I2 (g15080));
OR2X1 gate17150(.O (g34303), .I1 (g25768), .I2 (g34045));
OR2X1 gate17151(.O (g28316), .I1 (g27113), .I2 (g15804));
OR2X1 gate17152(.O (g27581), .I1 (g26161), .I2 (g24750));
OR2X1 gate17153(.O (g27450), .I1 (g2917), .I2 (g26483));
OR4X1 gate17154(.O (I30717), .I1 (g31787), .I2 (g32200), .I3 (g31940), .I4 (g31949));
OR2X1 gate17155(.O (g33577), .I1 (g33405), .I2 (g18430));
OR2X1 gate17156(.O (g30381), .I1 (g30126), .I2 (g18497));
OR2X1 gate17157(.O (g25575), .I1 (g24139), .I2 (g24140));
OR2X1 gate17158(.O (g28056), .I1 (g27230), .I2 (g18210));
OR2X1 gate17159(.O (g32359), .I1 (g29867), .I2 (g31298));
OR2X1 gate17160(.O (g27257), .I1 (g25904), .I2 (g24498));
OR2X1 gate17161(.O (g29166), .I1 (g27653), .I2 (g17153));
OR2X1 gate17162(.O (g25711), .I1 (g25105), .I2 (g21962));
OR2X1 gate17163(.O (g28611), .I1 (g27348), .I2 (g16485));
OR2X1 gate17164(.O (g24715), .I1 (g22189), .I2 (g22207));
OR2X1 gate17165(.O (g32358), .I1 (g29866), .I2 (g31297));
OR2X1 gate17166(.O (g34796), .I1 (g34745), .I2 (g18573));
OR2X1 gate17167(.O (g29892), .I1 (g28300), .I2 (g26120));
OR2X1 gate17168(.O (g27590), .I1 (g26179), .I2 (g24764));
OR2X1 gate17169(.O (g29476), .I1 (g28108), .I2 (g28112));
OR2X1 gate17170(.O (g29485), .I1 (g28535), .I2 (g27594));
OR2X1 gate17171(.O (g31906), .I1 (g31477), .I2 (g21953));
OR2X1 gate17172(.O (g30390), .I1 (g29985), .I2 (g18555));
OR2X1 gate17173(.O (g32344), .I1 (g29804), .I2 (g31266));
OR2X1 gate17174(.O (g31284), .I1 (g29575), .I2 (g28290));
OR2X1 gate17175(.O (g25606), .I1 (g24761), .I2 (g18117));
OR2X1 gate17176(.O (g28342), .I1 (g27134), .I2 (g15819));
OR2X1 gate17177(.O (g31304), .I1 (g29594), .I2 (g29608));
OR3X1 gate17178(.O (g29914), .I1 (g22531), .I2 (g22585), .I3 (I28147));
OR2X1 gate17179(.O (g21897), .I1 (g20095), .I2 (g15111));
OR2X1 gate17180(.O (g33622), .I1 (g33366), .I2 (g18791));
OR2X1 gate17181(.O (g33566), .I1 (g33356), .I2 (g18390));
OR2X1 gate17182(.O (g25750), .I1 (g25543), .I2 (g18802));
OR2X1 gate17183(.O (g26949), .I1 (g26356), .I2 (g24287));
OR2X1 gate17184(.O (g28650), .I1 (g27391), .I2 (g16598));
OR2X1 gate17185(.O (g30522), .I1 (g29332), .I2 (g22064));
OR2X1 gate17186(.O (g27150), .I1 (g25804), .I2 (g24400));
OR2X1 gate17187(.O (g34663), .I1 (g32028), .I2 (g34500));
OR2X1 gate17188(.O (g29239), .I1 (g28427), .I2 (g18297));
OR2X1 gate17189(.O (g26948), .I1 (g26399), .I2 (g24286));
OR2X1 gate17190(.O (g24354), .I1 (g23775), .I2 (g18823));
OR2X1 gate17191(.O (g27019), .I1 (g26822), .I2 (g14610));
OR2X1 gate17192(.O (g26904), .I1 (g26393), .I2 (g24221));
OR2X1 gate17193(.O (g29238), .I1 (g28178), .I2 (g18292));
OR2X1 gate17194(.O (g30483), .I1 (g30241), .I2 (g21979));
OR2X1 gate17195(.O (g30553), .I1 (g30205), .I2 (g22124));
OR2X1 gate17196(.O (g22901), .I1 (g19384), .I2 (g15745));
OR2X1 gate17197(.O (g28132), .I1 (g27932), .I2 (g27957));
OR2X1 gate17198(.O (g13997), .I1 (g11029), .I2 (g11036));
OR2X1 gate17199(.O (g29176), .I1 (g27661), .I2 (g17177));
OR2X1 gate17200(.O (g30536), .I1 (g30234), .I2 (g22082));
OR2X1 gate17201(.O (g26673), .I1 (g24433), .I2 (g10674));
OR2X1 gate17202(.O (g34040), .I1 (g33818), .I2 (g18737));
OR2X1 gate17203(.O (g33963), .I1 (g33830), .I2 (g18124));
OR2X1 gate17204(.O (g25663), .I1 (g24666), .I2 (g21788));
OR2X1 gate17205(.O (g34252), .I1 (g34146), .I2 (g18180));
OR2X1 gate17206(.O (g34621), .I1 (g34517), .I2 (g18583));
OR2X1 gate17207(.O (g28708), .I1 (g27462), .I2 (g16674));
OR2X1 gate17208(.O (g26933), .I1 (g26808), .I2 (g18551));
OR2X1 gate17209(.O (g28087), .I1 (g27255), .I2 (g18720));
OR2X1 gate17210(.O (g33576), .I1 (g33401), .I2 (g18423));
OR2X1 gate17211(.O (g33585), .I1 (g33411), .I2 (g18456));
OR2X1 gate17212(.O (g24211), .I1 (g23572), .I2 (g18138));
OR2X1 gate17213(.O (g28043), .I1 (g27323), .I2 (g21714));
OR2X1 gate17214(.O (g33554), .I1 (g33407), .I2 (g18353));
OR2X1 gate17215(.O (g32240), .I1 (g24757), .I2 (g31182));
OR2X1 gate17216(.O (g30397), .I1 (g29747), .I2 (g21756));
OR4X1 gate17217(.O (I26742), .I1 (g23430), .I2 (g23445), .I3 (g23458), .I4 (g23481));
OR2X1 gate17218(.O (g33609), .I1 (g33239), .I2 (g18615));
OR2X1 gate17219(.O (g29501), .I1 (g28583), .I2 (g27634));
OR2X1 gate17220(.O (g33312), .I1 (g29646), .I2 (g32170));
OR2X1 gate17221(.O (g30509), .I1 (g30210), .I2 (g22030));
OR2X1 gate17222(.O (g33608), .I1 (g33322), .I2 (g18537));
OR2X1 gate17223(.O (g28069), .I1 (g27564), .I2 (g21865));
OR2X1 gate17224(.O (g33115), .I1 (g32397), .I2 (g32401));
OR2X1 gate17225(.O (g25702), .I1 (g25068), .I2 (g21921));
OR2X1 gate17226(.O (g25757), .I1 (g25132), .I2 (g22104));
OR2X1 gate17227(.O (g28774), .I1 (g27536), .I2 (g16804));
OR2X1 gate17228(.O (g30508), .I1 (g30199), .I2 (g22029));
OR2X1 gate17229(.O (g31921), .I1 (g31508), .I2 (g22046));
OR2X1 gate17230(.O (g28068), .I1 (g27310), .I2 (g21838));
OR2X1 gate17231(.O (g32981), .I1 (g32425), .I2 (g18206));
OR2X1 gate17232(.O (g28375), .I1 (g27183), .I2 (g15851));
OR2X1 gate17233(.O (g33052), .I1 (g31961), .I2 (g21973));
OR2X1 gate17234(.O (g34634), .I1 (g34483), .I2 (g18691));
OR2X1 gate17235(.O (g25621), .I1 (g24523), .I2 (g18205));
OR2X1 gate17236(.O (g31745), .I1 (g29959), .I2 (g29973));
OR2X1 gate17237(.O (g21896), .I1 (g20084), .I2 (g15110));
OR2X1 gate17238(.O (g24250), .I1 (g22633), .I2 (g18295));
OR2X1 gate17239(.O (g26912), .I1 (g25946), .I2 (g18209));
OR2X1 gate17240(.O (g27231), .I1 (g25873), .I2 (g15699));
OR2X1 gate17241(.O (g29284), .I1 (g28554), .I2 (g18747));
OR2X1 gate17242(.O (g32395), .I1 (g31523), .I2 (g30049));
OR2X1 gate17243(.O (g24339), .I1 (g23690), .I2 (g18756));
OR2X1 gate17244(.O (g33973), .I1 (g33840), .I2 (g18344));
OR2X1 gate17245(.O (g29304), .I1 (g28588), .I2 (g18810));
OR2X1 gate17246(.O (g32262), .I1 (g31186), .I2 (g29710));
OR2X1 gate17247(.O (g23716), .I1 (g9194), .I2 (g20905));
OR2X1 gate17248(.O (g25673), .I1 (g24727), .I2 (g21830));
OR2X1 gate17249(.O (g32990), .I1 (g32281), .I2 (g18341));
OR3X1 gate17250(.O (I18417), .I1 (g14444), .I2 (g14414), .I3 (g14392));
OR2X1 gate17251(.O (g24338), .I1 (g23658), .I2 (g18755));
OR2X1 gate17252(.O (g11370), .I1 (g8807), .I2 (g550));
OR2X1 gate17253(.O (g30452), .I1 (g29891), .I2 (g21861));
OR2X1 gate17254(.O (g34452), .I1 (g34401), .I2 (g18665));
OR2X1 gate17255(.O (g13858), .I1 (g209), .I2 (g10685));
OR2X1 gate17256(.O (g33732), .I1 (g33104), .I2 (g32011));
OR2X1 gate17257(.O (g30311), .I1 (g28265), .I2 (g27265));
OR3X1 gate17258(.O (g24968), .I1 (g22360), .I2 (g22409), .I3 (g23389));
OR2X1 gate17259(.O (g25634), .I1 (g24559), .I2 (g18284));
OR2X1 gate17260(.O (g31761), .I1 (g30009), .I2 (g30028));
OR2X1 gate17261(.O (g33692), .I1 (g32400), .I2 (g33428));
OR2X1 gate17262(.O (g19475), .I1 (g16930), .I2 (g14126));
OR2X1 gate17263(.O (g27456), .I1 (g25978), .I2 (g24607));
OR2X1 gate17264(.O (g26396), .I1 (g24762), .I2 (g23062));
OR2X1 gate17265(.O (g28545), .I1 (g27301), .I2 (g26230));
OR2X1 gate17266(.O (g28078), .I1 (g27140), .I2 (g21880));
OR2X1 gate17267(.O (g33013), .I1 (g32283), .I2 (g18484));
OR2X1 gate17268(.O (g22669), .I1 (g7763), .I2 (g19525));
OR2X1 gate17269(.O (g32247), .I1 (g31168), .I2 (g29686));
OR3X1 gate17270(.O (I18543), .I1 (g14568), .I2 (g14540), .I3 (g14516));
OR2X1 gate17271(.O (g28086), .I1 (g27268), .I2 (g18702));
OR2X1 gate17272(.O (g32389), .I1 (g31496), .I2 (g29966));
OR2X1 gate17273(.O (g30350), .I1 (g30118), .I2 (g18334));
OR2X1 gate17274(.O (g34350), .I1 (g26048), .I2 (g34106));
OR2X1 gate17275(.O (g33539), .I1 (g33245), .I2 (g18178));
OR2X1 gate17276(.O (g32388), .I1 (g31495), .I2 (g29962));
OR2X1 gate17277(.O (g33005), .I1 (g32260), .I2 (g18432));
OR2X1 gate17278(.O (g27596), .I1 (g26207), .I2 (g24775));
OR2X1 gate17279(.O (g11025), .I1 (g2980), .I2 (g7831));
OR2X1 gate17280(.O (g28817), .I1 (g27548), .I2 (g16845));
OR2X1 gate17281(.O (g33538), .I1 (g33252), .I2 (g18144));
OR2X1 gate17282(.O (g28322), .I1 (g27117), .I2 (g15809));
OR2X1 gate17283(.O (g27243), .I1 (g25884), .I2 (g24475));
OR2X1 gate17284(.O (g30396), .I1 (g29856), .I2 (g21755));
OR2X1 gate17285(.O (g32251), .I1 (g30599), .I2 (g29352));
OR2X1 gate17286(.O (g13540), .I1 (g10822), .I2 (g10827));
OR2X1 gate17287(.O (g27431), .I1 (g24582), .I2 (g25977));
OR2X1 gate17288(.O (g20202), .I1 (g16211), .I2 (g13507));
OR2X1 gate17289(.O (g34731), .I1 (g34662), .I2 (g18272));
OR2X1 gate17290(.O (g29484), .I1 (g28124), .I2 (g22191));
OR2X1 gate17291(.O (g24202), .I1 (g22899), .I2 (g18106));
OR2X1 gate17292(.O (g26929), .I1 (g26635), .I2 (g18543));
OR2X1 gate17293(.O (g24257), .I1 (g22938), .I2 (g18310));
OR2X1 gate17294(.O (g30413), .I1 (g30001), .I2 (g21772));
OR2X1 gate17295(.O (g24496), .I1 (g24008), .I2 (g21557));
OR2X1 gate17296(.O (g31241), .I1 (g25959), .I2 (g29510));
OR2X1 gate17297(.O (g26928), .I1 (g26713), .I2 (g18541));
OR4X1 gate17298(.O (g17488), .I1 (g14361), .I2 (g14335), .I3 (g11954), .I4 (I18417));
OR2X1 gate17299(.O (g25592), .I1 (g24672), .I2 (g21706));
OR2X1 gate17300(.O (g25756), .I1 (g25112), .I2 (g22103));
OR2X1 gate17301(.O (g28561), .I1 (g27312), .I2 (g26250));
OR2X1 gate17302(.O (g28295), .I1 (g27094), .I2 (g15783));
OR2X1 gate17303(.O (g28680), .I1 (g27427), .I2 (g16633));
OR2X1 gate17304(.O (g32997), .I1 (g32269), .I2 (g18378));
OR2X1 gate17305(.O (g30405), .I1 (g29767), .I2 (g21764));
OR2X1 gate17306(.O (g16173), .I1 (g8796), .I2 (g13464));
OR2X1 gate17307(.O (g34405), .I1 (g34183), .I2 (g25103));
OR2X1 gate17308(.O (g33235), .I1 (g32040), .I2 (g30982));
OR2X1 gate17309(.O (g23317), .I1 (g19715), .I2 (g16191));
OR3X1 gate17310(.O (I22852), .I1 (g21459), .I2 (g21350), .I3 (g21339));
OR2X1 gate17311(.O (g29813), .I1 (g26020), .I2 (g28261));
OR2X1 gate17312(.O (g22679), .I1 (g19145), .I2 (g15701));
OR2X1 gate17313(.O (g23129), .I1 (g19500), .I2 (g15863));
OR2X1 gate17314(.O (g13699), .I1 (g10921), .I2 (g10947));
OR2X1 gate17315(.O (g34020), .I1 (g33904), .I2 (g18514));
OR2X1 gate17316(.O (g25731), .I1 (g25128), .I2 (g22014));
OR2X1 gate17317(.O (g28631), .I1 (g27372), .I2 (g16534));
OR4X1 gate17318(.O (I28567), .I1 (g29204), .I2 (g29205), .I3 (g29206), .I4 (g29207));
OR3X1 gate17319(.O (I24117), .I1 (g23088), .I2 (g23154), .I3 (g23172));
OR2X1 gate17320(.O (g32360), .I1 (g29868), .I2 (g31299));
OR2X1 gate17321(.O (g16506), .I1 (g13294), .I2 (g10966));
OR2X1 gate17322(.O (g15789), .I1 (g10819), .I2 (g13211));
OR4X1 gate17323(.O (I30261), .I1 (g29385), .I2 (g31376), .I3 (g30735), .I4 (g30825));
OR2X1 gate17324(.O (g34046), .I1 (g33906), .I2 (g33908));
OR2X1 gate17325(.O (g31882), .I1 (g31115), .I2 (g21776));
OR2X1 gate17326(.O (g33991), .I1 (g33885), .I2 (g18400));
OR2X1 gate17327(.O (g14078), .I1 (g10776), .I2 (g8703));
OR2X1 gate17328(.O (g20196), .I1 (g16207), .I2 (g13497));
OR2X1 gate17329(.O (g25691), .I1 (g24536), .I2 (g21890));
OR2X1 gate17330(.O (g27487), .I1 (g25990), .I2 (g24629));
OR2X1 gate17331(.O (g34282), .I1 (g26838), .I2 (g34214));
OR2X1 gate17332(.O (g23298), .I1 (g19693), .I2 (g16179));
OR2X1 gate17333(.O (g30357), .I1 (g30107), .I2 (g18366));
OR2X1 gate17334(.O (g28309), .I1 (g27106), .I2 (g15796));
OR2X1 gate17335(.O (g32220), .I1 (g31139), .I2 (g29633));
OR2X1 gate17336(.O (g26881), .I1 (g26629), .I2 (g24187));
OR2X1 gate17337(.O (g16927), .I1 (g13524), .I2 (g11126));
OR2X1 gate17338(.O (g25929), .I1 (g24395), .I2 (g22193));
OR2X1 gate17339(.O (g28308), .I1 (g27105), .I2 (g15795));
OR2X1 gate17340(.O (g27278), .I1 (g15786), .I2 (g25921));
OR2X1 gate17341(.O (g29692), .I1 (g28197), .I2 (g10873));
OR2X1 gate17342(.O (g24457), .I1 (g10902), .I2 (g22400));
OR2X1 gate17343(.O (g14977), .I1 (g10776), .I2 (g8703));
OR2X1 gate17344(.O (g25583), .I1 (g21666), .I2 (g24153));
OR2X1 gate17345(.O (g33584), .I1 (g33406), .I2 (g18449));
OR2X1 gate17346(.O (g34640), .I1 (g34487), .I2 (g18723));
OR2X1 gate17347(.O (g19274), .I1 (g17753), .I2 (g14791));
OR2X1 gate17348(.O (g19593), .I1 (g17145), .I2 (g14210));
OR2X1 gate17349(.O (g34803), .I1 (g34758), .I2 (g18590));
OR2X1 gate17350(.O (g28816), .I1 (g27547), .I2 (g16843));
OR2X1 gate17351(.O (g20077), .I1 (g16025), .I2 (g13320));
OR2X1 gate17352(.O (g23261), .I1 (g19660), .I2 (g16125));
OR2X1 gate17353(.O (g26890), .I1 (g26630), .I2 (g24196));
OR2X1 gate17354(.O (g28687), .I1 (g27434), .I2 (g16638));
OR2X1 gate17355(.O (g29539), .I1 (g2864), .I2 (g28220));
OR2X1 gate17356(.O (g32355), .I1 (g29855), .I2 (g31286));
OR2X1 gate17357(.O (g34881), .I1 (g34866), .I2 (g18187));
OR2X1 gate17358(.O (g24256), .I1 (g22873), .I2 (g18309));
OR2X1 gate17359(.O (g32370), .I1 (g29882), .I2 (g31312));
OR2X1 gate17360(.O (g28374), .I1 (g27181), .I2 (g15850));
OR2X1 gate17361(.O (g24280), .I1 (g23292), .I2 (g15109));
OR2X1 gate17362(.O (g25743), .I1 (g25110), .I2 (g22058));
OR2X1 gate17363(.O (g28643), .I1 (g27386), .I2 (g16592));
OR2X1 gate17364(.O (g27937), .I1 (g14506), .I2 (g26793));
OR2X1 gate17365(.O (g32996), .I1 (g32256), .I2 (g18377));
OR2X1 gate17366(.O (g34027), .I1 (g33718), .I2 (g18683));
OR2X1 gate17367(.O (g29241), .I1 (g28638), .I2 (g18332));
OR2X1 gate17368(.O (g13385), .I1 (g11967), .I2 (g9479));
ND2X1 gate17369(.O (g11980), .I1 (I14817), .I2 (I14818));
ND2X1 gate17370(.O (g13889), .I1 (g11566), .I2 (g11435));
ND2X1 gate17371(.O (g13980), .I1 (g10295), .I2 (g11435));
ND2X1 gate17372(.O (g12169), .I1 (g9804), .I2 (g5448));
ND2X1 gate17373(.O (I22761), .I1 (g11939), .I2 (I22760));
ND2X1 gate17374(.O (I13443), .I1 (g262), .I2 (I13442));
ND2X1 gate17375(.O (I14185), .I1 (g8442), .I2 (g3470));
ND4X1 gate17376(.O (g16719), .I1 (g3243), .I2 (g13700), .I3 (g3310), .I4 (g11350));
ND2X1 gate17377(.O (I14518), .I1 (g661), .I2 (I14516));
ND4X1 gate17378(.O (g10224), .I1 (g6661), .I2 (g6704), .I3 (g6675), .I4 (g6697));
ND2X1 gate17379(.O (g17595), .I1 (g8616), .I2 (g14367));
ND2X1 gate17380(.O (g22984), .I1 (g20114), .I2 (g2868));
ND2X1 gate17381(.O (I12346), .I1 (g3111), .I2 (I12344));
ND2X1 gate17382(.O (g12478), .I1 (I15299), .I2 (I15300));
ND4X1 gate17383(.O (g21432), .I1 (g17790), .I2 (g14820), .I3 (g17761), .I4 (g14780));
ND3X1 gate17384(.O (g28830), .I1 (g27886), .I2 (g7451), .I3 (g7369));
ND2X1 gate17385(.O (I14883), .I1 (g9500), .I2 (g5489));
ND2X1 gate17386(.O (g19474), .I1 (g11609), .I2 (g17794));
ND2X1 gate17387(.O (g11426), .I1 (g8742), .I2 (g4878));
ND2X1 gate17388(.O (g11190), .I1 (g8539), .I2 (g3447));
ND2X1 gate17389(.O (g9852), .I1 (g3684), .I2 (g4871));
ND2X1 gate17390(.O (g23342), .I1 (g6928), .I2 (g21163));
ND2X1 gate17391(.O (g27223), .I1 (I25908), .I2 (I25909));
ND2X1 gate17392(.O (I15089), .I1 (g2393), .I2 (I15087));
ND2X1 gate17393(.O (g22853), .I1 (g20219), .I2 (g2922));
ND2X1 gate17394(.O (g25003), .I1 (g21353), .I2 (g23462));
ND2X1 gate17395(.O (I15088), .I1 (g9832), .I2 (I15087));
ND2X1 gate17396(.O (g24916), .I1 (g19450), .I2 (g23154));
ND2X1 gate17397(.O (g25779), .I1 (g19694), .I2 (g24362));
ND2X1 gate17398(.O (g12084), .I1 (g2342), .I2 (g8211));
ND3X1 gate17399(.O (g28270), .I1 (g10504), .I2 (g26105), .I3 (g26987));
ND2X1 gate17400(.O (g22836), .I1 (g18918), .I2 (g2852));
ND2X1 gate17401(.O (g21330), .I1 (g11401), .I2 (g17157));
ND2X1 gate17402(.O (g20076), .I1 (g13795), .I2 (g16521));
ND4X1 gate17403(.O (g21365), .I1 (g15744), .I2 (g13119), .I3 (g15730), .I4 (g13100));
ND2X1 gate17404(.O (g23132), .I1 (g8155), .I2 (g19932));
ND2X1 gate17405(.O (I22683), .I1 (g11893), .I2 (g21434));
ND2X1 gate17406(.O (g28938), .I1 (g27796), .I2 (g8205));
ND2X1 gate17407(.O (g9825), .I1 (I13391), .I2 (I13392));
ND2X1 gate17408(.O (g7201), .I1 (I11865), .I2 (I11866));
ND4X1 gate17409(.O (g15719), .I1 (g5256), .I2 (g14490), .I3 (g5335), .I4 (g9780));
ND3X1 gate17410(.O (g27654), .I1 (g164), .I2 (g26598), .I3 (g23042));
ND2X1 gate17411(.O (g22864), .I1 (g7780), .I2 (g21156));
ND2X1 gate17412(.O (I20165), .I1 (g16246), .I2 (g990));
ND2X1 gate17413(.O (g14489), .I1 (g12126), .I2 (g5084));
ND2X1 gate17414(.O (g29082), .I1 (g27837), .I2 (g9694));
ND2X1 gate17415(.O (g25233), .I1 (g20838), .I2 (g23623));
ND2X1 gate17416(.O (g24942), .I1 (g20039), .I2 (g23172));
ND2X1 gate17417(.O (I26459), .I1 (g26576), .I2 (g14306));
ND3X1 gate17418(.O (g15832), .I1 (g7903), .I2 (g7479), .I3 (g13256));
ND4X1 gate17419(.O (g14830), .I1 (g6605), .I2 (g12211), .I3 (g6723), .I4 (g12721));
ND2X1 gate17420(.O (I32431), .I1 (g34056), .I2 (g34051));
ND2X1 gate17421(.O (g9972), .I1 (I13510), .I2 (I13511));
ND2X1 gate17422(.O (I20222), .I1 (g16272), .I2 (I20221));
ND3X1 gate17423(.O (g17748), .I1 (g562), .I2 (g14708), .I3 (g12323));
ND2X1 gate17424(.O (g11969), .I1 (g7252), .I2 (g1636));
ND2X1 gate17425(.O (g20734), .I1 (g14408), .I2 (g17312));
ND3X1 gate17426(.O (g28837), .I1 (g27800), .I2 (g7374), .I3 (g2197));
ND2X1 gate17427(.O (I25244), .I1 (g24744), .I2 (I25242));
ND3X1 gate17428(.O (g11968), .I1 (g837), .I2 (g9334), .I3 (g9086));
ND4X1 gate17429(.O (g13968), .I1 (g3913), .I2 (g11255), .I3 (g4031), .I4 (g11631));
ND2X1 gate17430(.O (g15045), .I1 (g12716), .I2 (g7142));
ND2X1 gate17431(.O (g12423), .I1 (I15242), .I2 (I15243));
ND4X1 gate17432(.O (g27587), .I1 (g24917), .I2 (g25018), .I3 (g24918), .I4 (g26857));
ND2X1 gate17433(.O (g20838), .I1 (g5041), .I2 (g17284));
ND2X1 gate17434(.O (g13855), .I1 (g4944), .I2 (g11804));
ND3X1 gate17435(.O (g19483), .I1 (g15969), .I2 (g10841), .I3 (g10922));
ND2X1 gate17436(.O (g10610), .I1 (g7462), .I2 (g7490));
ND2X1 gate17437(.O (g11411), .I1 (g9713), .I2 (g3625));
ND2X1 gate17438(.O (I13110), .I1 (g5808), .I2 (I13109));
ND2X1 gate17439(.O (g22642), .I1 (g7870), .I2 (g19560));
ND2X1 gate17440(.O (g12587), .I1 (g7497), .I2 (g6315));
ND2X1 gate17441(.O (g13870), .I1 (g11773), .I2 (g4732));
ND4X1 gate17442(.O (g13527), .I1 (g182), .I2 (g168), .I3 (g203), .I4 (g12812));
ND2X1 gate17443(.O (g23810), .I1 (I22973), .I2 (I22974));
ND2X1 gate17444(.O (g20619), .I1 (g14317), .I2 (g17217));
ND4X1 gate17445(.O (g16628), .I1 (g3602), .I2 (g11207), .I3 (g3618), .I4 (g13902));
ND2X1 gate17446(.O (I23119), .I1 (g20076), .I2 (I23118));
ND4X1 gate17447(.O (g10124), .I1 (g5276), .I2 (g5320), .I3 (g5290), .I4 (g5313));
ND2X1 gate17448(.O (g12000), .I1 (g8418), .I2 (g2610));
ND2X1 gate17449(.O (I23118), .I1 (g20076), .I2 (g417));
ND2X1 gate17450(.O (g22874), .I1 (g18918), .I2 (g2844));
ND2X1 gate17451(.O (g10939), .I1 (g7352), .I2 (g1459));
ND2X1 gate17452(.O (g13867), .I1 (g11312), .I2 (g8449));
ND4X1 gate17453(.O (g14686), .I1 (g5268), .I2 (g12059), .I3 (g5276), .I4 (g12239));
ND2X1 gate17454(.O (I12840), .I1 (g4222), .I2 (g4235));
ND2X1 gate17455(.O (g29049), .I1 (g9640), .I2 (g27779));
ND4X1 gate17456(.O (g16776), .I1 (g3945), .I2 (g13772), .I3 (g4012), .I4 (g11419));
ND2X1 gate17457(.O (g13315), .I1 (g1459), .I2 (g10715));
ND2X1 gate17458(.O (g11707), .I1 (g8718), .I2 (g4864));
ND2X1 gate17459(.O (I18530), .I1 (g1811), .I2 (I18529));
ND2X1 gate17460(.O (g20039), .I1 (g11250), .I2 (g17794));
ND2X1 gate17461(.O (I14609), .I1 (g8993), .I2 (g8678));
ND2X1 gate17462(.O (I13334), .I1 (g1687), .I2 (g1691));
ND2X1 gate17463(.O (g13257), .I1 (g1389), .I2 (g10544));
ND2X1 gate17464(.O (g29004), .I1 (g27933), .I2 (g8330));
ND4X1 gate17465(.O (g21459), .I1 (g17814), .I2 (g14854), .I3 (g17605), .I4 (g17581));
ND2X1 gate17466(.O (g11979), .I1 (g9861), .I2 (g5452));
ND3X1 gate17467(.O (g13496), .I1 (g1351), .I2 (g11336), .I3 (g11815));
ND3X1 gate17468(.O (g11590), .I1 (g6928), .I2 (g3990), .I3 (g4049));
ND3X1 gate17469(.O (g12639), .I1 (g10194), .I2 (g6682), .I3 (g6732));
ND2X1 gate17470(.O (g22712), .I1 (g18957), .I2 (g2864));
ND2X1 gate17471(.O (g23010), .I1 (g20516), .I2 (g2984));
ND2X1 gate17472(.O (g7897), .I1 (I12288), .I2 (I12289));
ND2X1 gate17473(.O (g24601), .I1 (g22957), .I2 (g2965));
ND2X1 gate17474(.O (g13986), .I1 (g10323), .I2 (g11747));
ND2X1 gate17475(.O (g12293), .I1 (g7436), .I2 (g5283));
ND2X1 gate17476(.O (g24677), .I1 (g22957), .I2 (g2975));
ND2X1 gate17477(.O (g12638), .I1 (g7514), .I2 (g6661));
ND2X1 gate17478(.O (g24975), .I1 (g21388), .I2 (g23363));
ND4X1 gate17479(.O (g10160), .I1 (g5623), .I2 (g5666), .I3 (g5637), .I4 (g5659));
ND4X1 gate17480(.O (g17712), .I1 (g5599), .I2 (g14425), .I3 (g5666), .I4 (g12301));
ND3X1 gate17481(.O (g12416), .I1 (g10133), .I2 (g7064), .I3 (g10166));
ND2X1 gate17482(.O (g14160), .I1 (g11626), .I2 (g8958));
ND3X1 gate17483(.O (g28853), .I1 (g27742), .I2 (g1636), .I3 (g7252));
ND4X1 gate17484(.O (g13067), .I1 (g5240), .I2 (g12059), .I3 (g5331), .I4 (g9780));
ND2X1 gate17485(.O (g28167), .I1 (g925), .I2 (g27046));
ND2X1 gate17486(.O (I18635), .I1 (g14713), .I2 (I18633));
ND2X1 gate17487(.O (g10617), .I1 (g10151), .I2 (g9909));
ND3X1 gate17488(.O (g16319), .I1 (g8224), .I2 (g8170), .I3 (g13736));
ND2X1 gate17489(.O (I32187), .I1 (g33661), .I2 (I32185));
ND2X1 gate17490(.O (I12252), .I1 (g1124), .I2 (I12251));
ND2X1 gate17491(.O (g14915), .I1 (g12553), .I2 (g10266));
ND2X1 gate17492(.O (g22941), .I1 (g20219), .I2 (g2970));
ND2X1 gate17493(.O (I17406), .I1 (g1472), .I2 (I17404));
ND2X1 gate17494(.O (g12578), .I1 (g7791), .I2 (g10341));
ND4X1 gate17495(.O (g27586), .I1 (g24924), .I2 (g24916), .I3 (g24905), .I4 (g26863));
ND2X1 gate17496(.O (g12014), .I1 (g7197), .I2 (g703));
ND2X1 gate17497(.O (g14075), .I1 (g11658), .I2 (g11527));
ND3X1 gate17498(.O (g15591), .I1 (g4332), .I2 (g4322), .I3 (g13202));
ND3X1 gate17499(.O (g28864), .I1 (g27886), .I2 (g7411), .I3 (g1996));
ND2X1 gate17500(.O (g10623), .I1 (g10181), .I2 (g9976));
ND4X1 gate17501(.O (g17675), .I1 (g5252), .I2 (g14399), .I3 (g5320), .I4 (g12239));
ND2X1 gate17502(.O (g23656), .I1 (I22800), .I2 (I22801));
ND2X1 gate17503(.O (g21353), .I1 (g11467), .I2 (g17157));
ND2X1 gate17504(.O (I13751), .I1 (g4584), .I2 (I13749));
ND2X1 gate17505(.O (g14782), .I1 (g12755), .I2 (g10491));
ND2X1 gate17506(.O (I14400), .I1 (g3654), .I2 (I14398));
ND2X1 gate17507(.O (g12116), .I1 (g2051), .I2 (g8255));
ND2X1 gate17508(.O (g14984), .I1 (g7812), .I2 (g12680));
ND4X1 gate17509(.O (g13866), .I1 (g3239), .I2 (g11194), .I3 (g3321), .I4 (g11519));
ND2X1 gate17510(.O (I18537), .I1 (g2236), .I2 (I18536));
ND3X1 gate17511(.O (g16281), .I1 (g4754), .I2 (g13937), .I3 (g12054));
ND3X1 gate17512(.O (g28900), .I1 (g27886), .I2 (g7451), .I3 (g2040));
ND2X1 gate17513(.O (g14822), .I1 (g12755), .I2 (g12632));
ND2X1 gate17514(.O (g14170), .I1 (g11715), .I2 (g11537));
ND3X1 gate17515(.O (g15844), .I1 (g14714), .I2 (g9340), .I3 (g12378));
ND2X1 gate17516(.O (I22972), .I1 (g9657), .I2 (g19638));
ND4X1 gate17517(.O (g21364), .I1 (g15787), .I2 (g15781), .I3 (g15753), .I4 (g13131));
ND2X1 gate17518(.O (I13391), .I1 (g1821), .I2 (I13390));
ND3X1 gate17519(.O (g13256), .I1 (g11846), .I2 (g11294), .I3 (g11812));
ND2X1 gate17520(.O (I13510), .I1 (g2089), .I2 (I13509));
ND2X1 gate17521(.O (g11923), .I1 (I14734), .I2 (I14735));
ND2X1 gate17522(.O (g12340), .I1 (g4888), .I2 (g8984));
ND2X1 gate17523(.O (g12035), .I1 (g10000), .I2 (g6144));
ND2X1 gate17524(.O (g13923), .I1 (g11692), .I2 (g11527));
ND2X1 gate17525(.O (I15300), .I1 (g1982), .I2 (I15298));
ND2X1 gate17526(.O (g9830), .I1 (I13402), .I2 (I13403));
ND2X1 gate17527(.O (g20186), .I1 (g16926), .I2 (g8177));
ND2X1 gate17528(.O (g20676), .I1 (g14379), .I2 (g17287));
ND2X1 gate17529(.O (g21289), .I1 (g14616), .I2 (g17493));
ND2X1 gate17530(.O (I12205), .I1 (g1135), .I2 (I12203));
ND2X1 gate17531(.O (g13102), .I1 (g7523), .I2 (g10759));
ND3X1 gate17532(.O (g25429), .I1 (g22417), .I2 (g1917), .I3 (g8302));
ND2X1 gate17533(.O (g23309), .I1 (g6905), .I2 (g21024));
ND3X1 gate17534(.O (g28874), .I1 (g27907), .I2 (g7424), .I3 (g2421));
ND2X1 gate17535(.O (g29121), .I1 (g9755), .I2 (g27886));
ND2X1 gate17536(.O (g21288), .I1 (g14616), .I2 (g17492));
ND2X1 gate17537(.O (g7582), .I1 (g1361), .I2 (g1373));
ND2X1 gate17538(.O (I13442), .I1 (g262), .I2 (g239));
ND3X1 gate17539(.O (g13066), .I1 (g4430), .I2 (g7178), .I3 (g10590));
ND4X1 gate17540(.O (g24936), .I1 (g20186), .I2 (g20173), .I3 (g23379), .I4 (g14029));
ND3X1 gate17541(.O (g31262), .I1 (g767), .I2 (g29916), .I3 (g11679));
ND2X1 gate17542(.O (g10022), .I1 (g6474), .I2 (g6466));
ND2X1 gate17543(.O (g14864), .I1 (g7791), .I2 (g10421));
ND2X1 gate17544(.O (g8769), .I1 (g691), .I2 (g714));
ND2X1 gate17545(.O (g7227), .I1 (g4584), .I2 (g4593));
ND2X1 gate17546(.O (I32186), .I1 (g33665), .I2 (I32185));
ND2X1 gate17547(.O (g12523), .I1 (g7563), .I2 (g6346));
ND3X1 gate17548(.O (g28892), .I1 (g27779), .I2 (g1772), .I3 (g7275));
ND2X1 gate17549(.O (g13854), .I1 (g4765), .I2 (g11797));
ND2X1 gate17550(.O (g11511), .I1 (I14481), .I2 (I14482));
ND2X1 gate17551(.O (I14991), .I1 (g9685), .I2 (g6527));
ND2X1 gate17552(.O (g8967), .I1 (g4264), .I2 (g4258));
ND4X1 gate17553(.O (g13511), .I1 (g182), .I2 (g174), .I3 (g203), .I4 (g12812));
ND2X1 gate17554(.O (g20216), .I1 (I20487), .I2 (I20488));
ND3X1 gate17555(.O (g14254), .I1 (g11968), .I2 (g11933), .I3 (g11951));
ND3X1 gate17556(.O (g28914), .I1 (g27937), .I2 (g7462), .I3 (g2555));
ND2X1 gate17557(.O (g29134), .I1 (g9762), .I2 (g27907));
ND3X1 gate17558(.O (g28907), .I1 (g27858), .I2 (g2361), .I3 (g2287));
ND2X1 gate17559(.O (g12222), .I1 (g8310), .I2 (g2028));
ND2X1 gate17560(.O (g29028), .I1 (g27933), .I2 (g8381));
ND2X1 gate17561(.O (g22852), .I1 (g18957), .I2 (g2856));
ND2X1 gate17562(.O (g14101), .I1 (g11653), .I2 (g11729));
ND2X1 gate17563(.O (g25002), .I1 (g19474), .I2 (g23154));
ND2X1 gate17564(.O (I29297), .I1 (g12117), .I2 (I29295));
ND3X1 gate17565(.O (g14177), .I1 (g11741), .I2 (g11721), .I3 (g753));
ND2X1 gate17566(.O (g11480), .I1 (g10323), .I2 (g8906));
ND2X1 gate17567(.O (I26460), .I1 (g26576), .I2 (I26459));
ND2X1 gate17568(.O (I22946), .I1 (g19620), .I2 (I22944));
ND2X1 gate17569(.O (I18536), .I1 (g2236), .I2 (g14642));
ND2X1 gate17570(.O (I15287), .I1 (g10061), .I2 (g6697));
ND2X1 gate17571(.O (I14206), .I1 (g3821), .I2 (I14204));
ND4X1 gate17572(.O (g16956), .I1 (g3925), .I2 (g13824), .I3 (g4019), .I4 (g11631));
ND2X1 gate17573(.O (I26093), .I1 (g26055), .I2 (g13539));
ND2X1 gate17574(.O (I15307), .I1 (g10116), .I2 (I15306));
ND2X1 gate17575(.O (g23195), .I1 (g20136), .I2 (g37));
ND2X1 gate17576(.O (g13307), .I1 (g1116), .I2 (g10695));
ND2X1 gate17577(.O (I15243), .I1 (g6351), .I2 (I15241));
ND4X1 gate17578(.O (g16181), .I1 (g13475), .I2 (g13495), .I3 (g13057), .I4 (g13459));
ND2X1 gate17579(.O (g12351), .I1 (I15194), .I2 (I15195));
ND2X1 gate17580(.O (g24814), .I1 (g20011), .I2 (g23167));
ND2X1 gate17581(.O (g22312), .I1 (g907), .I2 (g19063));
ND3X1 gate17582(.O (g28935), .I1 (g27800), .I2 (g2227), .I3 (g7328));
ND2X1 gate17583(.O (g24807), .I1 (I23979), .I2 (I23980));
ND2X1 gate17584(.O (I15341), .I1 (g10154), .I2 (I15340));
ND2X1 gate17585(.O (g14665), .I1 (g12604), .I2 (g12798));
ND2X1 gate17586(.O (g24974), .I1 (g21301), .I2 (g23363));
ND2X1 gate17587(.O (g31997), .I1 (g22306), .I2 (g30580));
ND2X1 gate17588(.O (g14008), .I1 (g11610), .I2 (g11435));
ND2X1 gate17589(.O (I14399), .I1 (g8542), .I2 (I14398));
ND2X1 gate17590(.O (I22760), .I1 (g11939), .I2 (g21434));
ND2X1 gate17591(.O (g9258), .I1 (I13044), .I2 (I13045));
ND2X1 gate17592(.O (g22921), .I1 (g20219), .I2 (g2950));
ND3X1 gate17593(.O (g15715), .I1 (g336), .I2 (g305), .I3 (g13385));
ND2X1 gate17594(.O (g17312), .I1 (g7297), .I2 (g14248));
ND2X1 gate17595(.O (g25995), .I1 (g24621), .I2 (g22853));
ND2X1 gate17596(.O (g14892), .I1 (g12700), .I2 (g12515));
ND4X1 gate17597(.O (g17608), .I1 (g5953), .I2 (g12067), .I3 (g5969), .I4 (g14701));
ND2X1 gate17598(.O (I14398), .I1 (g8542), .I2 (g3654));
ND2X1 gate17599(.O (g15572), .I1 (g12969), .I2 (g7219));
ND2X1 gate17600(.O (I18634), .I1 (g2504), .I2 (I18633));
ND2X1 gate17601(.O (I15335), .I1 (g2116), .I2 (I15333));
ND2X1 gate17602(.O (g34056), .I1 (I31984), .I2 (I31985));
ND4X1 gate17603(.O (g14570), .I1 (g3933), .I2 (g11255), .I3 (g4023), .I4 (g8595));
ND2X1 gate17604(.O (g11993), .I1 (g1894), .I2 (g8302));
ND4X1 gate17605(.O (g13993), .I1 (g3961), .I2 (g11255), .I3 (g3969), .I4 (g11419));
ND2X1 gate17606(.O (I23963), .I1 (g13631), .I2 (I23961));
ND2X1 gate17607(.O (g9975), .I1 (I13519), .I2 (I13520));
ND2X1 gate17608(.O (g21124), .I1 (g5731), .I2 (g17393));
ND2X1 gate17609(.O (I14332), .I1 (g9966), .I2 (I14330));
ND2X1 gate17610(.O (g13667), .I1 (g3723), .I2 (g11119));
ND4X1 gate17611(.O (g13131), .I1 (g6243), .I2 (g12101), .I3 (g6377), .I4 (g10003));
ND2X1 gate17612(.O (g10567), .I1 (g1862), .I2 (g7405));
ND2X1 gate17613(.O (g20007), .I1 (g11512), .I2 (g17794));
ND2X1 gate17614(.O (I23585), .I1 (g22409), .I2 (g4332));
ND4X1 gate17615(.O (g28349), .I1 (g27074), .I2 (g24770), .I3 (g27187), .I4 (g19644));
ND2X1 gate17616(.O (g29719), .I1 (g28406), .I2 (g13739));
ND2X1 gate17617(.O (g21294), .I1 (g11324), .I2 (g17157));
ND3X1 gate17618(.O (g25498), .I1 (g22498), .I2 (g2610), .I3 (g8418));
ND2X1 gate17619(.O (g28906), .I1 (g27796), .I2 (g8150));
ND2X1 gate17620(.O (g13210), .I1 (g7479), .I2 (g10521));
ND2X1 gate17621(.O (g34650), .I1 (I32757), .I2 (I32758));
ND4X1 gate17622(.O (g16625), .I1 (g3203), .I2 (g13700), .I3 (g3274), .I4 (g11519));
ND4X1 gate17623(.O (g17732), .I1 (g3937), .I2 (g13824), .I3 (g4012), .I4 (g13933));
ND4X1 gate17624(.O (g10185), .I1 (g5969), .I2 (g6012), .I3 (g5983), .I4 (g6005));
ND2X1 gate17625(.O (g11443), .I1 (g9916), .I2 (g3649));
ND2X1 gate17626(.O (g12436), .I1 (I15263), .I2 (I15264));
ND2X1 gate17627(.O (g11279), .I1 (g8504), .I2 (g3443));
ND4X1 gate17628(.O (g14519), .I1 (g3889), .I2 (g11225), .I3 (g4000), .I4 (g8595));
ND2X1 gate17629(.O (I29296), .I1 (g29495), .I2 (I29295));
ND2X1 gate17630(.O (g14675), .I1 (g12317), .I2 (g9898));
ND2X1 gate17631(.O (I25219), .I1 (g482), .I2 (g24718));
ND4X1 gate17632(.O (g27593), .I1 (g24972), .I2 (g24950), .I3 (g24906), .I4 (g26861));
ND2X1 gate17633(.O (I26419), .I1 (g14247), .I2 (I26417));
ND2X1 gate17634(.O (I22755), .I1 (g21434), .I2 (I22753));
ND2X1 gate17635(.O (g12073), .I1 (g10058), .I2 (g6490));
ND2X1 gate17636(.O (g14154), .I1 (g11669), .I2 (g8958));
ND4X1 gate17637(.O (g17761), .I1 (g6291), .I2 (g14529), .I3 (g6358), .I4 (g12423));
ND2X1 gate17638(.O (I26418), .I1 (g26519), .I2 (I26417));
ND2X1 gate17639(.O (g13469), .I1 (g4983), .I2 (g10862));
ND2X1 gate17640(.O (g25432), .I1 (g12374), .I2 (g22384));
ND2X1 gate17641(.O (g10935), .I1 (g1459), .I2 (g7352));
ND2X1 gate17642(.O (g14637), .I1 (g12255), .I2 (g9815));
ND2X1 gate17643(.O (I15306), .I1 (g10116), .I2 (g2407));
ND2X1 gate17644(.O (g16296), .I1 (g9360), .I2 (g13501));
ND2X1 gate17645(.O (g25271), .I1 (I24462), .I2 (I24463));
ND2X1 gate17646(.O (g7133), .I1 (I11825), .I2 (I11826));
ND3X1 gate17647(.O (g12464), .I1 (g10169), .I2 (g7087), .I3 (g10191));
ND2X1 gate17648(.O (g7846), .I1 (g4843), .I2 (g4878));
ND4X1 gate17649(.O (g12797), .I1 (g10275), .I2 (g7655), .I3 (g7643), .I4 (g7627));
ND2X1 gate17650(.O (I22794), .I1 (g21434), .I2 (I22792));
ND2X1 gate17651(.O (I22845), .I1 (g12113), .I2 (I22844));
ND2X1 gate17652(.O (g7803), .I1 (I12204), .I2 (I12205));
ND2X1 gate17653(.O (g31950), .I1 (g7285), .I2 (g30573));
ND2X1 gate17654(.O (g12292), .I1 (g4698), .I2 (g8933));
ND2X1 gate17655(.O (g9461), .I1 (I13140), .I2 (I13141));
ND2X1 gate17656(.O (g12153), .I1 (g2610), .I2 (g8330));
ND2X1 gate17657(.O (g25199), .I1 (I24364), .I2 (I24365));
ND2X1 gate17658(.O (I22899), .I1 (g12193), .I2 (g21228));
ND2X1 gate17659(.O (g8829), .I1 (g5011), .I2 (g4836));
ND2X1 gate17660(.O (g11975), .I1 (g8267), .I2 (g8316));
ND2X1 gate17661(.O (I12204), .I1 (g1094), .I2 (I12203));
ND3X1 gate17662(.O (g19513), .I1 (g15969), .I2 (g10841), .I3 (g10922));
ND2X1 gate17663(.O (g23617), .I1 (I22761), .I2 (I22762));
ND2X1 gate17664(.O (g15024), .I1 (g12780), .I2 (g10421));
ND2X1 gate17665(.O (I20205), .I1 (g11147), .I2 (I20203));
ND2X1 gate17666(.O (g12136), .I1 (I14992), .I2 (I14993));
ND2X1 gate17667(.O (I22719), .I1 (g21434), .I2 (I22717));
ND2X1 gate17668(.O (g9904), .I1 (I13443), .I2 (I13444));
ND4X1 gate17669(.O (g13143), .I1 (g10695), .I2 (g7661), .I3 (g979), .I4 (g1061));
ND2X1 gate17670(.O (I13453), .I1 (g1955), .I2 (I13452));
ND2X1 gate17671(.O (I22718), .I1 (g11916), .I2 (I22717));
ND3X1 gate17672(.O (g33394), .I1 (g10159), .I2 (g4474), .I3 (g32426));
ND2X1 gate17673(.O (g11169), .I1 (I14229), .I2 (I14230));
ND2X1 gate17674(.O (I29315), .I1 (g12154), .I2 (I29313));
ND2X1 gate17675(.O (I15168), .I1 (g9823), .I2 (I15166));
ND2X1 gate17676(.O (g13884), .I1 (g11797), .I2 (g4727));
ND3X1 gate17677(.O (g11410), .I1 (g6875), .I2 (g6895), .I3 (g8696));
ND2X1 gate17678(.O (g23623), .I1 (g9364), .I2 (g20717));
ND2X1 gate17679(.O (g9391), .I1 (I13110), .I2 (I13111));
ND2X1 gate17680(.O (I15363), .I1 (g10182), .I2 (g2675));
ND2X1 gate17681(.O (g8124), .I1 (I12402), .I2 (I12403));
ND2X1 gate17682(.O (g24362), .I1 (g21370), .I2 (g22136));
ND3X1 gate17683(.O (g11479), .I1 (g6875), .I2 (g3288), .I3 (g3347));
ND2X1 gate17684(.O (g23782), .I1 (g2741), .I2 (g21062));
ND2X1 gate17685(.O (g13666), .I1 (g11190), .I2 (g8441));
ND4X1 gate17686(.O (g13479), .I1 (g12686), .I2 (g12639), .I3 (g12590), .I4 (g12526));
ND2X1 gate17687(.O (g8069), .I1 (I12373), .I2 (I12374));
ND2X1 gate17688(.O (I32517), .I1 (g34424), .I2 (I32516));
ND2X1 gate17689(.O (g13217), .I1 (g4082), .I2 (g10808));
ND2X1 gate17690(.O (g10622), .I1 (g10178), .I2 (g9973));
ND2X1 gate17691(.O (g10566), .I1 (g7315), .I2 (g7356));
ND4X1 gate17692(.O (g13478), .I1 (g12511), .I2 (g12460), .I3 (g12414), .I4 (g12344));
ND2X1 gate17693(.O (I13565), .I1 (g2648), .I2 (I13564));
ND2X1 gate17694(.O (I13464), .I1 (g2384), .I2 (I13462));
ND3X1 gate17695(.O (g13486), .I1 (g10862), .I2 (g4983), .I3 (g4966));
ND2X1 gate17696(.O (g25258), .I1 (I24439), .I2 (I24440));
ND2X1 gate17697(.O (g23266), .I1 (g18918), .I2 (g2894));
ND4X1 gate17698(.O (g13580), .I1 (g11849), .I2 (g7503), .I3 (g7922), .I4 (g10544));
ND2X1 gate17699(.O (g10653), .I1 (g10204), .I2 (g10042));
ND2X1 gate17700(.O (g14139), .I1 (g11626), .I2 (g11584));
ND4X1 gate17701(.O (g16741), .I1 (g3207), .I2 (g13765), .I3 (g3303), .I4 (g11519));
ND2X1 gate17702(.O (I14789), .I1 (g9891), .I2 (I14788));
ND2X1 gate17703(.O (g23167), .I1 (g8219), .I2 (g19981));
ND4X1 gate17704(.O (g13084), .I1 (g5587), .I2 (g12093), .I3 (g5677), .I4 (g9864));
ND3X1 gate17705(.O (g28973), .I1 (g27907), .I2 (g2465), .I3 (g7387));
ND4X1 gate17706(.O (g14636), .I1 (g5595), .I2 (g12029), .I3 (g5677), .I4 (g12563));
ND2X1 gate17707(.O (I14788), .I1 (g9891), .I2 (g6167));
ND4X1 gate17708(.O (g14333), .I1 (g12042), .I2 (g12014), .I3 (g11990), .I4 (g11892));
ND2X1 gate17709(.O (I17462), .I1 (g1300), .I2 (I17460));
ND4X1 gate17710(.O (g21401), .I1 (g17755), .I2 (g14730), .I3 (g17712), .I4 (g14695));
ND4X1 gate17711(.O (g27796), .I1 (g21228), .I2 (g25263), .I3 (g26424), .I4 (g26171));
ND4X1 gate17712(.O (g20236), .I1 (g16875), .I2 (g14014), .I3 (g16625), .I4 (g16604));
ND2X1 gate17713(.O (g12796), .I1 (g4467), .I2 (g6961));
ND2X1 gate17714(.O (g9654), .I1 (g2485), .I2 (g2453));
ND3X1 gate17715(.O (g15867), .I1 (g14714), .I2 (g9417), .I3 (g9340));
ND3X1 gate17716(.O (g25337), .I1 (g22342), .I2 (g1648), .I3 (g8187));
ND2X1 gate17717(.O (g28934), .I1 (g27882), .I2 (g14641));
ND4X1 gate17718(.O (g14664), .I1 (g5220), .I2 (g12059), .I3 (g5339), .I4 (g12497));
ND4X1 gate17719(.O (g16196), .I1 (g13496), .I2 (g13513), .I3 (g13079), .I4 (g13476));
ND4X1 gate17720(.O (g11676), .I1 (g358), .I2 (g8944), .I3 (g376), .I4 (g385));
ND3X1 gate17721(.O (g34545), .I1 (g11679), .I2 (g794), .I3 (g34354));
ND2X1 gate17722(.O (I22871), .I1 (g12150), .I2 (g21228));
ND2X1 gate17723(.O (g11953), .I1 (g8195), .I2 (g8241));
ND2X1 gate17724(.O (g13676), .I1 (g11834), .I2 (g11283));
ND2X1 gate17725(.O (g23616), .I1 (I22754), .I2 (I22755));
ND2X1 gate17726(.O (g29355), .I1 (g24383), .I2 (g28109));
ND2X1 gate17727(.O (g15581), .I1 (g7232), .I2 (g12999));
ND2X1 gate17728(.O (g10585), .I1 (g1996), .I2 (g7451));
ND2X1 gate17729(.O (g9595), .I1 (g2351), .I2 (g2319));
ND2X1 gate17730(.O (g23748), .I1 (I22872), .I2 (I22873));
ND2X1 gate17731(.O (I14291), .I1 (g3835), .I2 (I14289));
ND2X1 gate17732(.O (g11936), .I1 (g8241), .I2 (g1783));
ND2X1 gate17733(.O (I15334), .I1 (g10152), .I2 (I15333));
ND2X1 gate17734(.O (g12192), .I1 (g8267), .I2 (g2319));
ND2X1 gate17735(.O (g10609), .I1 (g10111), .I2 (g9826));
ND2X1 gate17736(.O (I13109), .I1 (g5808), .I2 (g5813));
ND2X1 gate17737(.O (g22940), .I1 (g18918), .I2 (g2860));
ND2X1 gate17738(.O (I12097), .I1 (g1339), .I2 (I12096));
ND2X1 gate17739(.O (g25425), .I1 (g20081), .I2 (g23172));
ND3X1 gate17740(.O (g12522), .I1 (g10133), .I2 (g5990), .I3 (g6040));
ND2X1 gate17741(.O (g23809), .I1 (I22966), .I2 (I22967));
ND4X1 gate17742(.O (g17744), .I1 (g6303), .I2 (g14529), .I3 (g6373), .I4 (g12672));
ND2X1 gate17743(.O (I17447), .I1 (g13336), .I2 (I17446));
ND3X1 gate17744(.O (g28207), .I1 (g12546), .I2 (g26131), .I3 (g27977));
ND3X1 gate17745(.O (g17399), .I1 (g9626), .I2 (g9574), .I3 (g14535));
ND2X1 gate17746(.O (g14921), .I1 (g12492), .I2 (g10266));
ND4X1 gate17747(.O (g15741), .I1 (g5244), .I2 (g14490), .I3 (g5320), .I4 (g14631));
ND2X1 gate17748(.O (I32516), .I1 (g34424), .I2 (g34422));
ND2X1 gate17749(.O (g9629), .I1 (g6462), .I2 (g6466));
ND2X1 gate17750(.O (I13750), .I1 (g4608), .I2 (I13749));
ND2X1 gate17751(.O (g14813), .I1 (g7766), .I2 (g12824));
ND2X1 gate17752(.O (g11543), .I1 (g9714), .I2 (g3969));
ND2X1 gate17753(.O (I12850), .I1 (g4277), .I2 (I12848));
ND4X1 gate17754(.O (g13909), .I1 (g11396), .I2 (g8847), .I3 (g11674), .I4 (g8803));
ND2X1 gate17755(.O (g23733), .I1 (g20751), .I2 (g11178));
ND4X1 gate17756(.O (g15735), .I1 (g5547), .I2 (g14425), .I3 (g5659), .I4 (g9864));
ND3X1 gate17757(.O (g15877), .I1 (g14833), .I2 (g9340), .I3 (g12543));
ND2X1 gate17758(.O (g9800), .I1 (g5436), .I2 (g5428));
ND4X1 gate17759(.O (g14674), .I1 (g5941), .I2 (g12067), .I3 (g6023), .I4 (g12614));
ND3X1 gate17760(.O (g11117), .I1 (g8087), .I2 (g8186), .I3 (g8239));
ND3X1 gate17761(.O (g29025), .I1 (g27937), .I2 (g2629), .I3 (g7462));
ND2X1 gate17762(.O (g13000), .I1 (g7228), .I2 (g10598));
ND2X1 gate17763(.O (I22754), .I1 (g11937), .I2 (I22753));
ND2X1 gate17764(.O (g29540), .I1 (g28336), .I2 (g13464));
ND2X1 gate17765(.O (g23630), .I1 (g20739), .I2 (g11123));
ND3X1 gate17766(.O (g22833), .I1 (g1193), .I2 (g19560), .I3 (g10666));
ND2X1 gate17767(.O (g15695), .I1 (g1266), .I2 (g13125));
ND2X1 gate17768(.O (g25532), .I1 (g21360), .I2 (g23363));
ND2X1 gate17769(.O (g15018), .I1 (g12739), .I2 (g12515));
ND2X1 gate17770(.O (I13390), .I1 (g1821), .I2 (g1825));
ND2X1 gate17771(.O (g14732), .I1 (g12662), .I2 (g12515));
ND2X1 gate17772(.O (g24905), .I1 (g534), .I2 (g23088));
ND2X1 gate17773(.O (I15242), .I1 (g10003), .I2 (I15241));
ND2X1 gate17774(.O (g19857), .I1 (g13628), .I2 (g16296));
ND2X1 gate17775(.O (g17500), .I1 (g14573), .I2 (g14548));
ND2X1 gate17776(.O (I15123), .I1 (g2102), .I2 (I15121));
ND2X1 gate17777(.O (g14761), .I1 (g12651), .I2 (g10281));
ND2X1 gate17778(.O (I22844), .I1 (g12113), .I2 (g21228));
ND4X1 gate17779(.O (g21555), .I1 (g17846), .I2 (g14946), .I3 (g17686), .I4 (g17650));
ND4X1 gate17780(.O (g16854), .I1 (g3965), .I2 (g13824), .I3 (g3976), .I4 (g8595));
ND2X1 gate17781(.O (g11974), .I1 (g2185), .I2 (g8259));
ND2X1 gate17782(.O (g31671), .I1 (I29262), .I2 (I29263));
ND4X1 gate17783(.O (g27933), .I1 (g21228), .I2 (g25356), .I3 (g26424), .I4 (g26236));
ND3X1 gate17784(.O (g19549), .I1 (g15969), .I2 (g10841), .I3 (g10899));
ND4X1 gate17785(.O (g8806), .I1 (g358), .I2 (g370), .I3 (g376), .I4 (g385));
ND2X1 gate17786(.O (g11639), .I1 (g8933), .I2 (g4722));
ND2X1 gate17787(.O (g9823), .I1 (I13383), .I2 (I13384));
ND2X1 gate17788(.O (g12933), .I1 (g7150), .I2 (g10515));
ND2X1 gate17789(.O (I25907), .I1 (g26256), .I2 (g24782));
ND4X1 gate17790(.O (g10207), .I1 (g6315), .I2 (g6358), .I3 (g6329), .I4 (g6351));
ND2X1 gate17791(.O (I20204), .I1 (g16246), .I2 (I20203));
ND2X1 gate17792(.O (g26752), .I1 (g9397), .I2 (g25189));
ND2X1 gate17793(.O (g14005), .I1 (g11514), .I2 (g11729));
ND4X1 gate17794(.O (g16660), .I1 (g3953), .I2 (g11225), .I3 (g3969), .I4 (g13933));
ND2X1 gate17795(.O (I26439), .I1 (g26549), .I2 (I26438));
ND4X1 gate17796(.O (g17605), .I1 (g5559), .I2 (g14425), .I3 (g5630), .I4 (g12563));
ND2X1 gate17797(.O (g11992), .I1 (g7275), .I2 (g1772));
ND2X1 gate17798(.O (I29314), .I1 (g29501), .I2 (I29313));
ND2X1 gate17799(.O (I26438), .I1 (g26549), .I2 (g14271));
ND2X1 gate17800(.O (I12096), .I1 (g1339), .I2 (g1322));
ND2X1 gate17801(.O (I23962), .I1 (g23184), .I2 (I23961));
ND2X1 gate17802(.O (I17446), .I1 (g13336), .I2 (g956));
ND3X1 gate17803(.O (g28206), .I1 (g12546), .I2 (g26105), .I3 (g27985));
ND2X1 gate17804(.O (g25309), .I1 (g22384), .I2 (g12021));
ND2X1 gate17805(.O (I13564), .I1 (g2648), .I2 (g2652));
ND2X1 gate17806(.O (I12730), .I1 (g4287), .I2 (I12728));
ND2X1 gate17807(.O (g7857), .I1 (I12241), .I2 (I12242));
ND3X1 gate17808(.O (g28758), .I1 (g27779), .I2 (g7356), .I3 (g7275));
ND2X1 gate17809(.O (I29269), .I1 (g29486), .I2 (g12050));
ND4X1 gate17810(.O (g14771), .I1 (g5961), .I2 (g12129), .I3 (g5969), .I4 (g12351));
ND2X1 gate17811(.O (g8913), .I1 (I12877), .I2 (I12878));
ND3X1 gate17812(.O (g11442), .I1 (g8644), .I2 (g3288), .I3 (g3343));
ND2X1 gate17813(.O (I13183), .I1 (g6500), .I2 (I13182));
ND2X1 gate17814(.O (g14683), .I1 (g12553), .I2 (g12443));
ND4X1 gate17815(.O (g17514), .I1 (g3917), .I2 (g13772), .I3 (g4019), .I4 (g8595));
ND2X1 gate17816(.O (g25495), .I1 (g12483), .I2 (g22472));
ND2X1 gate17817(.O (g12592), .I1 (I15364), .I2 (I15365));
ND2X1 gate17818(.O (I13509), .I1 (g2089), .I2 (g2093));
ND2X1 gate17819(.O (I14247), .I1 (g1322), .I2 (g8091));
ND2X1 gate17820(.O (I15041), .I1 (g9752), .I2 (g1834));
ND2X1 gate17821(.O (g10515), .I1 (g10337), .I2 (g5022));
ND2X1 gate17822(.O (I13851), .I1 (g862), .I2 (I13850));
ND2X1 gate17823(.O (g25985), .I1 (g24631), .I2 (g23956));
ND2X1 gate17824(.O (g14882), .I1 (g12558), .I2 (g12453));
ND2X1 gate17825(.O (g34424), .I1 (I32440), .I2 (I32441));
ND2X1 gate17826(.O (g14407), .I1 (g12008), .I2 (g9807));
ND3X1 gate17827(.O (g19856), .I1 (g13626), .I2 (g16278), .I3 (g8105));
ND2X1 gate17828(.O (I23951), .I1 (g13603), .I2 (I23949));
ND2X1 gate17829(.O (I15340), .I1 (g10154), .I2 (g2541));
ND2X1 gate17830(.O (g26255), .I1 (g8075), .I2 (g24779));
ND2X1 gate17831(.O (g12152), .I1 (g2485), .I2 (g8324));
ND2X1 gate17832(.O (g22325), .I1 (g1252), .I2 (g19140));
ND2X1 gate17833(.O (g13983), .I1 (g11658), .I2 (g8906));
ND4X1 gate17834(.O (g16694), .I1 (g3905), .I2 (g13772), .I3 (g3976), .I4 (g11631));
ND4X1 gate17835(.O (g17788), .I1 (g5232), .I2 (g14490), .I3 (g5327), .I4 (g12497));
ND2X1 gate17836(.O (g12413), .I1 (g7521), .I2 (g5654));
ND2X1 gate17837(.O (g10584), .I1 (g7362), .I2 (g7405));
ND2X1 gate17838(.O (g28406), .I1 (g27064), .I2 (g13675));
ND2X1 gate17839(.O (I13452), .I1 (g1955), .I2 (g1959));
ND3X1 gate17840(.O (g28962), .I1 (g27886), .I2 (g2040), .I3 (g7369));
ND2X1 gate17841(.O (I29279), .I1 (g12081), .I2 (I29277));
ND3X1 gate17842(.O (g28500), .I1 (g590), .I2 (g27629), .I3 (g12323));
ND2X1 gate17843(.O (g10759), .I1 (g7537), .I2 (g324));
ND3X1 gate17844(.O (g15721), .I1 (g7564), .I2 (g311), .I3 (g13385));
ND2X1 gate17845(.O (I29278), .I1 (g29488), .I2 (I29277));
ND2X1 gate17846(.O (I14766), .I1 (g5821), .I2 (I14764));
ND2X1 gate17847(.O (I15130), .I1 (g2527), .I2 (I15128));
ND2X1 gate17848(.O (I15193), .I1 (g9935), .I2 (g6005));
ND2X1 gate17849(.O (I29286), .I1 (g12085), .I2 (I29284));
ND2X1 gate17850(.O (g14758), .I1 (g7704), .I2 (g12405));
ND2X1 gate17851(.O (g11130), .I1 (g1221), .I2 (g7918));
ND2X1 gate17852(.O (g14082), .I1 (g11697), .I2 (g11537));
ND2X1 gate17853(.O (g11193), .I1 (I14258), .I2 (I14259));
ND3X1 gate17854(.O (g13130), .I1 (g1351), .I2 (g11815), .I3 (g11336));
ND2X1 gate17855(.O (g14107), .I1 (g11571), .I2 (g11527));
ND3X1 gate17856(.O (g16278), .I1 (g8102), .I2 (g8057), .I3 (g13664));
ND2X1 gate17857(.O (g12020), .I1 (g2028), .I2 (g8365));
ND3X1 gate17858(.O (g19611), .I1 (g1070), .I2 (g1199), .I3 (g15995));
ND2X1 gate17859(.O (g23139), .I1 (g21163), .I2 (g10756));
ND3X1 gate17860(.O (g16306), .I1 (g4944), .I2 (g13971), .I3 (g12088));
ND2X1 gate17861(.O (I12261), .I1 (g1454), .I2 (g1448));
ND2X1 gate17862(.O (g14940), .I1 (g12744), .I2 (g12581));
ND2X1 gate17863(.O (I18627), .I1 (g14712), .I2 (I18625));
ND3X1 gate17864(.O (g13475), .I1 (g1008), .I2 (g11294), .I3 (g11786));
ND2X1 gate17865(.O (g14848), .I1 (g12651), .I2 (g12453));
ND4X1 gate17866(.O (g27282), .I1 (g11192), .I2 (g26269), .I3 (g26248), .I4 (g479));
ND4X1 gate17867(.O (g21415), .I1 (g17773), .I2 (g14771), .I3 (g17740), .I4 (g14739));
ND4X1 gate17868(.O (g16815), .I1 (g3909), .I2 (g13824), .I3 (g4005), .I4 (g11631));
ND4X1 gate17869(.O (g13727), .I1 (g174), .I2 (g203), .I3 (g168), .I4 (g12812));
ND4X1 gate17870(.O (g15734), .I1 (g5228), .I2 (g12059), .I3 (g5290), .I4 (g14631));
ND2X1 gate17871(.O (g14804), .I1 (g12651), .I2 (g12798));
ND2X1 gate17872(.O (g25255), .I1 (g20979), .I2 (g23659));
ND2X1 gate17873(.O (I13731), .I1 (g4537), .I2 (I13729));
ND2X1 gate17874(.O (g12357), .I1 (g7439), .I2 (g6329));
ND2X1 gate17875(.O (g31978), .I1 (g30580), .I2 (g15591));
ND2X1 gate17876(.O (I22824), .I1 (g21434), .I2 (I22822));
ND2X1 gate17877(.O (I15253), .I1 (g10078), .I2 (g1848));
ND2X1 gate17878(.O (g24621), .I1 (g22957), .I2 (g2927));
ND2X1 gate17879(.O (I18681), .I1 (g2638), .I2 (I18680));
ND2X1 gate17880(.O (g14962), .I1 (g12558), .I2 (g10281));
ND2X1 gate17881(.O (g13600), .I1 (g3021), .I2 (g11039));
ND2X1 gate17882(.O (I22931), .I1 (g21228), .I2 (I22929));
ND2X1 gate17883(.O (g9645), .I1 (g2060), .I2 (g2028));
ND2X1 gate17884(.O (g23576), .I1 (I22718), .I2 (I22719));
ND2X1 gate17885(.O (g19764), .I1 (I20166), .I2 (I20167));
ND2X1 gate17886(.O (g11952), .I1 (g1624), .I2 (g8187));
ND2X1 gate17887(.O (I15175), .I1 (g9977), .I2 (I15174));
ND2X1 gate17888(.O (I32757), .I1 (g34469), .I2 (I32756));
ND2X1 gate17889(.O (I14370), .I1 (g3303), .I2 (I14368));
ND2X1 gate17890(.O (g26782), .I1 (g9467), .I2 (g25203));
ND2X1 gate17891(.O (g13821), .I1 (g11251), .I2 (g8340));
ND2X1 gate17892(.O (g14048), .I1 (g11658), .I2 (g11483));
ND2X1 gate17893(.O (I15264), .I1 (g2273), .I2 (I15262));
ND2X1 gate17894(.O (g22755), .I1 (g20136), .I2 (g18984));
ND2X1 gate17895(.O (g28421), .I1 (g27074), .I2 (g13715));
ND3X1 gate17896(.O (g26352), .I1 (g744), .I2 (g24875), .I3 (g11679));
ND2X1 gate17897(.O (I12271), .I1 (g956), .I2 (I12269));
ND3X1 gate17898(.O (g13264), .I1 (g11869), .I2 (g11336), .I3 (g11849));
ND2X1 gate17899(.O (g24933), .I1 (g19466), .I2 (g23154));
ND4X1 gate17900(.O (g13137), .I1 (g10699), .I2 (g7675), .I3 (g1322), .I4 (g1404));
ND4X1 gate17901(.O (g13516), .I1 (g11533), .I2 (g11490), .I3 (g11444), .I4 (g11412));
ND2X1 gate17902(.O (g15039), .I1 (g12755), .I2 (g7142));
ND2X1 gate17903(.O (g29060), .I1 (g9649), .I2 (g27800));
ND4X1 gate17904(.O (g17755), .I1 (g5619), .I2 (g14522), .I3 (g5630), .I4 (g9864));
ND2X1 gate17905(.O (g13873), .I1 (g11566), .I2 (g11729));
ND2X1 gate17906(.O (I31974), .I1 (g33631), .I2 (I31972));
ND2X1 gate17907(.O (g14947), .I1 (g12785), .I2 (g10491));
ND2X1 gate17908(.O (g10605), .I1 (g2555), .I2 (g7490));
ND2X1 gate17909(.O (g12482), .I1 (I15307), .I2 (I15308));
ND3X1 gate17910(.O (g25470), .I1 (g22457), .I2 (g2051), .I3 (g8365));
ND2X1 gate17911(.O (g13834), .I1 (g4754), .I2 (g11773));
ND3X1 gate17912(.O (g16321), .I1 (g4955), .I2 (g13996), .I3 (g12088));
ND2X1 gate17913(.O (g10951), .I1 (g7845), .I2 (g7868));
ND3X1 gate17914(.O (g28920), .I1 (g27779), .I2 (g1802), .I3 (g7315));
ND2X1 gate17915(.O (g24574), .I1 (g22709), .I2 (g22687));
ND2X1 gate17916(.O (g14234), .I1 (g9177), .I2 (g11881));
ND2X1 gate17917(.O (g31706), .I1 (I29270), .I2 (I29271));
ND2X1 gate17918(.O (I18626), .I1 (g2079), .I2 (I18625));
ND3X1 gate17919(.O (g28946), .I1 (g27907), .I2 (g2495), .I3 (g2421));
ND2X1 gate17920(.O (g25467), .I1 (g12432), .I2 (g22417));
ND2X1 gate17921(.O (g23761), .I1 (I22893), .I2 (I22894));
ND2X1 gate17922(.O (g23692), .I1 (g9501), .I2 (g20995));
ND2X1 gate17923(.O (g27380), .I1 (I26071), .I2 (I26072));
ND2X1 gate17924(.O (g12356), .I1 (g7438), .I2 (g6012));
ND2X1 gate17925(.O (g9591), .I1 (g1926), .I2 (g1894));
ND3X1 gate17926(.O (g12999), .I1 (g4392), .I2 (g10476), .I3 (g4401));
ND3X1 gate17927(.O (g11320), .I1 (g4633), .I2 (g4621), .I3 (g7202));
ND2X1 gate17928(.O (g25984), .I1 (g24567), .I2 (g22668));
ND2X1 gate17929(.O (g19886), .I1 (g11403), .I2 (g17794));
ND2X1 gate17930(.O (I15122), .I1 (g9910), .I2 (I15121));
ND2X1 gate17931(.O (g13346), .I1 (g4854), .I2 (g11012));
ND2X1 gate17932(.O (g19792), .I1 (I20204), .I2 (I20205));
ND2X1 gate17933(.O (I14957), .I1 (g6181), .I2 (I14955));
ND3X1 gate17934(.O (g26053), .I1 (g22875), .I2 (g24677), .I3 (g22941));
ND3X1 gate17935(.O (g13464), .I1 (g10831), .I2 (g4793), .I3 (g4776));
ND2X1 gate17936(.O (g13797), .I1 (g8102), .I2 (g11273));
ND2X1 gate17937(.O (g11292), .I1 (I14331), .I2 (I14332));
ND2X1 gate17938(.O (I32756), .I1 (g34469), .I2 (g25779));
ND2X1 gate17939(.O (g11153), .I1 (I14205), .I2 (I14206));
ND2X1 gate17940(.O (g29094), .I1 (g27858), .I2 (g9700));
ND3X1 gate17941(.O (g12449), .I1 (g7004), .I2 (g5297), .I3 (g5352));
ND2X1 gate17942(.O (I14290), .I1 (g8282), .I2 (I14289));
ND2X1 gate17943(.O (g11409), .I1 (g9842), .I2 (g3298));
ND2X1 gate17944(.O (I22894), .I1 (g21228), .I2 (I22892));
ND2X1 gate17945(.O (I14427), .I1 (g8595), .I2 (g4005));
ND4X1 gate17946(.O (g14829), .I1 (g6621), .I2 (g12137), .I3 (g6675), .I4 (g12471));
ND2X1 gate17947(.O (I31983), .I1 (g33653), .I2 (g33648));
ND2X1 gate17948(.O (g14434), .I1 (g6415), .I2 (g11945));
ND2X1 gate17949(.O (g29018), .I1 (g9586), .I2 (g27742));
ND2X1 gate17950(.O (I12878), .I1 (g4180), .I2 (I12876));
ND2X1 gate17951(.O (g10946), .I1 (g1489), .I2 (g7876));
ND3X1 gate17952(.O (g28927), .I1 (g27837), .I2 (g1906), .I3 (g7322));
ND4X1 gate17953(.O (g14946), .I1 (g6247), .I2 (g12173), .I3 (g6346), .I4 (g12672));
ND2X1 gate17954(.O (g9750), .I1 (I13335), .I2 (I13336));
ND2X1 gate17955(.O (I11826), .I1 (g4601), .I2 (I11824));
ND2X1 gate17956(.O (g14344), .I1 (g5377), .I2 (g11885));
ND2X1 gate17957(.O (g24583), .I1 (g22753), .I2 (g22711));
ND2X1 gate17958(.O (I13182), .I1 (g6500), .I2 (g6505));
ND2X1 gate17959(.O (I17496), .I1 (g1448), .I2 (I17494));
ND3X1 gate17960(.O (g28903), .I1 (g27800), .I2 (g2197), .I3 (g7280));
ND2X1 gate17961(.O (g14682), .I1 (g4933), .I2 (g11780));
ND2X1 gate17962(.O (g12149), .I1 (g8205), .I2 (g2185));
ND2X1 gate17963(.O (I14481), .I1 (g10074), .I2 (I14480));
ND3X1 gate17964(.O (g28755), .I1 (g27742), .I2 (g7268), .I3 (g1592));
ND2X1 gate17965(.O (g12148), .I1 (g2060), .I2 (g8310));
ND4X1 gate17966(.O (g13109), .I1 (g6279), .I2 (g12173), .I3 (g6369), .I4 (g10003));
ND4X1 gate17967(.O (g16772), .I1 (g3558), .I2 (g13799), .I3 (g3654), .I4 (g11576));
ND2X1 gate17968(.O (g24787), .I1 (g3391), .I2 (g23079));
ND3X1 gate17969(.O (g29001), .I1 (g27937), .I2 (g2599), .I3 (g7431));
ND4X1 gate17970(.O (g13108), .I1 (g5551), .I2 (g12029), .I3 (g5685), .I4 (g9864));
ND2X1 gate17971(.O (g12343), .I1 (g7470), .I2 (g5630));
ND3X1 gate17972(.O (g13283), .I1 (g12440), .I2 (g12399), .I3 (g9843));
ND2X1 gate17973(.O (I22801), .I1 (g21434), .I2 (I22799));
ND3X1 gate17974(.O (g11492), .I1 (g6928), .I2 (g6941), .I3 (g8756));
ND3X1 gate17975(.O (g12971), .I1 (g9024), .I2 (g8977), .I3 (g10664));
ND2X1 gate17976(.O (I12545), .I1 (g191), .I2 (I12544));
ND2X1 gate17977(.O (g9528), .I1 (I13183), .I2 (I13184));
ND2X1 gate17978(.O (g12369), .I1 (g9049), .I2 (g637));
ND2X1 gate17979(.O (g28395), .I1 (g27074), .I2 (g13655));
ND2X1 gate17980(.O (I14956), .I1 (g9620), .I2 (I14955));
ND2X1 gate17981(.O (g11381), .I1 (g9660), .I2 (g3274));
ND2X1 gate17982(.O (g28899), .I1 (g27833), .I2 (g14612));
ND2X1 gate17983(.O (I18529), .I1 (g1811), .I2 (g14640));
ND2X1 gate17984(.O (g28990), .I1 (g27882), .I2 (g8310));
ND3X1 gate17985(.O (g17220), .I1 (g9369), .I2 (g9298), .I3 (g14376));
ND2X1 gate17986(.O (I15174), .I1 (g9977), .I2 (g2661));
ND2X1 gate17987(.O (g29157), .I1 (g9835), .I2 (g27937));
ND3X1 gate17988(.O (g17246), .I1 (g9439), .I2 (g9379), .I3 (g14405));
ND3X1 gate17989(.O (g12412), .I1 (g10044), .I2 (g5297), .I3 (g5348));
ND2X1 gate17990(.O (I26049), .I1 (g25997), .I2 (g13500));
ND3X1 gate17991(.O (g26382), .I1 (g577), .I2 (g24953), .I3 (g12323));
ND3X1 gate17992(.O (g33930), .I1 (g33394), .I2 (g12767), .I3 (g9848));
ND2X1 gate17993(.O (g22754), .I1 (g20114), .I2 (g19376));
ND2X1 gate17994(.O (g33838), .I1 (g33083), .I2 (g4369));
ND2X1 gate17995(.O (g14927), .I1 (g12695), .I2 (g10281));
ND2X1 gate17996(.O (g16586), .I1 (g13851), .I2 (g13823));
ND2X1 gate17997(.O (I22866), .I1 (g21228), .I2 (I22864));
ND2X1 gate17998(.O (g21345), .I1 (g11429), .I2 (g17157));
ND3X1 gate17999(.O (g27582), .I1 (g10857), .I2 (g26131), .I3 (g26105));
ND2X1 gate18000(.O (g9372), .I1 (g5080), .I2 (g5084));
ND3X1 gate18001(.O (g28861), .I1 (g27837), .I2 (g7405), .I3 (g1906));
ND2X1 gate18002(.O (I20461), .I1 (g17515), .I2 (I20460));
ND3X1 gate18003(.O (g25476), .I1 (g22472), .I2 (g2476), .I3 (g8373));
ND2X1 gate18004(.O (g8359), .I1 (I12545), .I2 (I12546));
ND2X1 gate18005(.O (g24662), .I1 (g22957), .I2 (g2955));
ND2X1 gate18006(.O (I24461), .I1 (g23796), .I2 (g14437));
ND2X1 gate18007(.O (g10604), .I1 (g7424), .I2 (g7456));
ND4X1 gate18008(.O (g15751), .I1 (g5591), .I2 (g14522), .I3 (g5666), .I4 (g14669));
ND4X1 gate18009(.O (g10755), .I1 (g7352), .I2 (g7675), .I3 (g1322), .I4 (g1404));
ND2X1 gate18010(.O (g24890), .I1 (g13852), .I2 (g22929));
ND2X1 gate18011(.O (g14755), .I1 (g12593), .I2 (g12772));
ND3X1 gate18012(.O (g19495), .I1 (g15969), .I2 (g10841), .I3 (g7781));
ND2X1 gate18013(.O (g27925), .I1 (I26439), .I2 (I26440));
ND2X1 gate18014(.O (I22923), .I1 (g21284), .I2 (I22921));
ND2X1 gate18015(.O (g29660), .I1 (g28448), .I2 (g9582));
ND3X1 gate18016(.O (g20248), .I1 (g17056), .I2 (g14146), .I3 (g14123));
ND2X1 gate18017(.O (g16275), .I1 (g9291), .I2 (g13480));
ND2X1 gate18018(.O (g14981), .I1 (g12785), .I2 (g12632));
ND2X1 gate18019(.O (I14211), .I1 (g9252), .I2 (g9295));
ND2X1 gate18020(.O (g9334), .I1 (g827), .I2 (g832));
ND2X1 gate18021(.O (g12112), .I1 (g8139), .I2 (g1624));
ND2X1 gate18022(.O (I17923), .I1 (g13378), .I2 (g1478));
ND3X1 gate18023(.O (g33306), .I1 (g776), .I2 (g32212), .I3 (g11679));
ND4X1 gate18024(.O (g11326), .I1 (g8993), .I2 (g376), .I3 (g365), .I4 (g370));
ND2X1 gate18025(.O (g20081), .I1 (g11325), .I2 (g17794));
ND2X1 gate18026(.O (g14794), .I1 (g12492), .I2 (g12772));
ND2X1 gate18027(.O (g14845), .I1 (g12558), .I2 (g12798));
ND2X1 gate18028(.O (I14497), .I1 (g9020), .I2 (g8737));
ND2X1 gate18029(.O (I24365), .I1 (g14320), .I2 (I24363));
ND2X1 gate18030(.O (I13850), .I1 (g862), .I2 (g7397));
ND4X1 gate18031(.O (g13040), .I1 (g5196), .I2 (g12002), .I3 (g5308), .I4 (g9780));
ND2X1 gate18032(.O (g13948), .I1 (g11610), .I2 (g8864));
ND2X1 gate18033(.O (g14899), .I1 (g12744), .I2 (g10421));
ND2X1 gate18034(.O (g29085), .I1 (g9694), .I2 (g27837));
ND2X1 gate18035(.O (g28997), .I1 (g27903), .I2 (g8324));
ND2X1 gate18036(.O (g25382), .I1 (g12333), .I2 (g22342));
ND2X1 gate18037(.O (I12289), .I1 (g1300), .I2 (I12287));
ND4X1 gate18038(.O (g14898), .I1 (g5901), .I2 (g12129), .I3 (g6000), .I4 (g12614));
ND2X1 gate18039(.O (I32204), .I1 (g33670), .I2 (I32202));
ND2X1 gate18040(.O (I23950), .I1 (g23162), .I2 (I23949));
ND2X1 gate18041(.O (g15014), .I1 (g12785), .I2 (g12680));
ND2X1 gate18042(.O (I12288), .I1 (g1484), .I2 (I12287));
ND2X1 gate18043(.O (g24380), .I1 (I23601), .I2 (I23602));
ND2X1 gate18044(.O (g12429), .I1 (g7473), .I2 (g6675));
ND2X1 gate18045(.O (g14521), .I1 (g12170), .I2 (g5428));
ND2X1 gate18046(.O (I25221), .I1 (g24718), .I2 (I25219));
ND2X1 gate18047(.O (g12428), .I1 (g7472), .I2 (g6358));
ND3X1 gate18048(.O (g28871), .I1 (g27858), .I2 (g7418), .I3 (g2331));
ND2X1 gate18049(.O (I17885), .I1 (g1135), .I2 (I17883));
ND2X1 gate18050(.O (g9908), .I1 (I13453), .I2 (I13454));
ND2X1 gate18051(.O (g22902), .I1 (g18957), .I2 (g2848));
ND2X1 gate18052(.O (I16780), .I1 (g12332), .I2 (I16778));
ND2X1 gate18053(.O (g10573), .I1 (g7992), .I2 (g8179));
ND2X1 gate18054(.O (g9567), .I1 (g6116), .I2 (g6120));
ND2X1 gate18055(.O (g14861), .I1 (g12744), .I2 (g10341));
ND2X1 gate18056(.O (g14573), .I1 (g9506), .I2 (g12249));
ND2X1 gate18057(.O (g24932), .I1 (g19886), .I2 (g23172));
ND4X1 gate18058(.O (g15720), .I1 (g5917), .I2 (g14497), .I3 (g6019), .I4 (g9935));
ND3X1 gate18059(.O (g11933), .I1 (g837), .I2 (g9334), .I3 (g7197));
ND2X1 gate18060(.O (I14855), .I1 (g5142), .I2 (I14853));
ND2X1 gate18061(.O (g14045), .I1 (g11571), .I2 (g11747));
ND2X1 gate18062(.O (g29335), .I1 (g25540), .I2 (g28131));
ND2X1 gate18063(.O (g13634), .I1 (g11797), .I2 (g11261));
ND2X1 gate18064(.O (g13851), .I1 (g8224), .I2 (g11360));
ND2X1 gate18065(.O (g27317), .I1 (g24793), .I2 (g26255));
ND2X1 gate18066(.O (I12374), .I1 (g3462), .I2 (I12372));
ND2X1 gate18067(.O (g25215), .I1 (I24384), .I2 (I24385));
ND2X1 gate18068(.O (g7850), .I1 (g554), .I2 (g807));
ND2X1 gate18069(.O (g12317), .I1 (g10026), .I2 (g6486));
ND2X1 gate18070(.O (g29694), .I1 (g28391), .I2 (g13709));
ND2X1 gate18071(.O (g14098), .I1 (g11566), .I2 (g8864));
ND2X1 gate18072(.O (g17699), .I1 (I18681), .I2 (I18682));
ND2X1 gate18073(.O (g25439), .I1 (g22498), .I2 (g12122));
ND3X1 gate18074(.O (g28911), .I1 (g27907), .I2 (g7456), .I3 (g2465));
ND2X1 gate18075(.O (g23972), .I1 (g7097), .I2 (g20751));
ND3X1 gate18076(.O (g17290), .I1 (g9506), .I2 (g9449), .I3 (g14431));
ND2X1 gate18077(.O (I29253), .I1 (g29482), .I2 (g12017));
ND2X1 gate18078(.O (g29131), .I1 (g27907), .I2 (g9762));
ND2X1 gate18079(.O (I15213), .I1 (g10035), .I2 (I15212));
ND2X1 gate18080(.O (I12842), .I1 (g4235), .I2 (I12840));
ND2X1 gate18081(.O (g25349), .I1 (g22432), .I2 (g12051));
ND2X1 gate18082(.O (g12245), .I1 (g7344), .I2 (g5637));
ND2X1 gate18083(.O (g12323), .I1 (g9480), .I2 (g640));
ND2X1 gate18084(.O (I14714), .I1 (g5128), .I2 (I14712));
ND2X1 gate18085(.O (g22661), .I1 (g20136), .I2 (g94));
ND2X1 gate18086(.O (I13730), .I1 (g4534), .I2 (I13729));
ND4X1 gate18087(.O (g27775), .I1 (g21228), .I2 (g25262), .I3 (g26424), .I4 (g26166));
ND3X1 gate18088(.O (g16236), .I1 (g13573), .I2 (g13554), .I3 (g13058));
ND2X1 gate18089(.O (I14257), .I1 (g8154), .I2 (g3133));
ND3X1 gate18090(.O (g28950), .I1 (g27937), .I2 (g7490), .I3 (g2599));
ND2X1 gate18091(.O (I15051), .I1 (g9759), .I2 (g2259));
ND2X1 gate18092(.O (I14818), .I1 (g6513), .I2 (I14816));
ND2X1 gate18093(.O (g9724), .I1 (g5092), .I2 (g5084));
ND2X1 gate18094(.O (g22715), .I1 (g20114), .I2 (g2999));
ND2X1 gate18095(.O (I23120), .I1 (g417), .I2 (I23118));
ND2X1 gate18096(.O (g24620), .I1 (g22902), .I2 (g22874));
ND4X1 gate18097(.O (g14871), .I1 (g6653), .I2 (g12211), .I3 (g6661), .I4 (g12471));
ND2X1 gate18098(.O (I12544), .I1 (g191), .I2 (g194));
ND2X1 gate18099(.O (g13756), .I1 (g203), .I2 (g12812));
ND2X1 gate18100(.O (I18680), .I1 (g2638), .I2 (g14752));
ND2X1 gate18101(.O (g12232), .I1 (g8804), .I2 (g4878));
ND3X1 gate18102(.O (g16264), .I1 (g518), .I2 (g9158), .I3 (g13223));
ND2X1 gate18103(.O (g19875), .I1 (g13667), .I2 (g16316));
ND2X1 gate18104(.O (I22930), .I1 (g12223), .I2 (I22929));
ND3X1 gate18105(.O (g26052), .I1 (g22714), .I2 (g24662), .I3 (g22921));
ND2X1 gate18106(.O (g26745), .I1 (g6856), .I2 (g25317));
ND4X1 gate18107(.O (g17572), .I1 (g3598), .I2 (g13799), .I3 (g3676), .I4 (g8542));
ND2X1 gate18108(.O (g11350), .I1 (I14369), .I2 (I14370));
ND2X1 gate18109(.O (I22965), .I1 (g12288), .I2 (g21228));
ND2X1 gate18110(.O (I32433), .I1 (g34051), .I2 (I32431));
ND2X1 gate18111(.O (g24369), .I1 (I23586), .I2 (I23587));
ND2X1 gate18112(.O (g12512), .I1 (g7766), .I2 (g10312));
ND2X1 gate18113(.O (g21359), .I1 (g11509), .I2 (g17157));
ND2X1 gate18114(.O (g13846), .I1 (g1116), .I2 (g10649));
ND2X1 gate18115(.O (g10472), .I1 (I13851), .I2 (I13852));
ND2X1 gate18116(.O (g11396), .I1 (g8713), .I2 (g4688));
ND2X1 gate18117(.O (I12270), .I1 (g1141), .I2 (I12269));
ND2X1 gate18118(.O (I14735), .I1 (g5475), .I2 (I14733));
ND3X1 gate18119(.O (g19455), .I1 (g15969), .I2 (g10841), .I3 (g7781));
ND4X1 gate18120(.O (g20133), .I1 (g17668), .I2 (g17634), .I3 (g17597), .I4 (g14569));
ND2X1 gate18121(.O (g17297), .I1 (g2729), .I2 (g14291));
ND2X1 gate18122(.O (g21344), .I1 (g11428), .I2 (g17157));
ND4X1 gate18123(.O (g11405), .I1 (g2741), .I2 (g2735), .I3 (g6856), .I4 (g2748));
ND4X1 gate18124(.O (g15781), .I1 (g6267), .I2 (g12173), .I3 (g6329), .I4 (g14745));
ND2X1 gate18125(.O (g20011), .I1 (g3731), .I2 (g16476));
ND2X1 gate18126(.O (g14776), .I1 (g12780), .I2 (g12622));
ND3X1 gate18127(.O (g28203), .I1 (g12546), .I2 (g27985), .I3 (g27977));
ND3X1 gate18128(.O (g10754), .I1 (g7936), .I2 (g7913), .I3 (g8411));
ND2X1 gate18129(.O (g29015), .I1 (g27742), .I2 (g9586));
ND2X1 gate18130(.O (g13929), .I1 (g11669), .I2 (g11763));
ND2X1 gate18131(.O (I12219), .I1 (g1478), .I2 (I12217));
ND2X1 gate18132(.O (g25200), .I1 (g5742), .I2 (g23642));
ND2X1 gate18133(.O (g14825), .I1 (g12806), .I2 (g12680));
ND2X1 gate18134(.O (g14950), .I1 (g7812), .I2 (g12632));
ND2X1 gate18135(.O (g11020), .I1 (g9187), .I2 (g9040));
ND2X1 gate18136(.O (g12080), .I1 (g1917), .I2 (g8201));
ND4X1 gate18137(.O (g13928), .I1 (g3562), .I2 (g11238), .I3 (g3680), .I4 (g11576));
ND2X1 gate18138(.O (I12218), .I1 (g1437), .I2 (I12217));
ND2X1 gate18139(.O (g14858), .I1 (g7766), .I2 (g12515));
ND2X1 gate18140(.O (g19782), .I1 (I20188), .I2 (I20189));
ND2X1 gate18141(.O (g29556), .I1 (g28349), .I2 (g13486));
ND2X1 gate18142(.O (g31747), .I1 (I29296), .I2 (I29297));
ND2X1 gate18143(.O (g14151), .I1 (g11692), .I2 (g11483));
ND2X1 gate18144(.O (g14996), .I1 (g12662), .I2 (g10312));
ND2X1 gate18145(.O (g24925), .I1 (g20092), .I2 (g23154));
ND2X1 gate18146(.O (g24958), .I1 (g21330), .I2 (g23462));
ND4X1 gate18147(.O (g17520), .I1 (g5260), .I2 (g12002), .I3 (g5276), .I4 (g14631));
ND2X1 gate18148(.O (g12461), .I1 (g7536), .I2 (g6000));
ND2X1 gate18149(.O (I24364), .I1 (g23687), .I2 (I24363));
ND3X1 gate18150(.O (g12342), .I1 (g7004), .I2 (g7018), .I3 (g10129));
ND2X1 gate18151(.O (I22937), .I1 (g12226), .I2 (I22936));
ND2X1 gate18152(.O (I26395), .I1 (g14227), .I2 (I26393));
ND2X1 gate18153(.O (I14923), .I1 (g9558), .I2 (g5835));
ND2X1 gate18154(.O (g12145), .I1 (g8195), .I2 (g1760));
ND2X1 gate18155(.O (g11302), .I1 (g9496), .I2 (g3281));
ND2X1 gate18156(.O (I15105), .I1 (g9780), .I2 (g5313));
ND2X1 gate18157(.O (I23980), .I1 (g13670), .I2 (I23978));
ND2X1 gate18158(.O (g24944), .I1 (g21354), .I2 (g23363));
ND4X1 gate18159(.O (g13105), .I1 (g10671), .I2 (g7675), .I3 (g1322), .I4 (g1404));
ND2X1 gate18160(.O (I16779), .I1 (g11292), .I2 (I16778));
ND2X1 gate18161(.O (I12470), .I1 (g392), .I2 (I12468));
ND2X1 gate18162(.O (g9092), .I1 (g3004), .I2 (g3050));
ND2X1 gate18163(.O (I16778), .I1 (g11292), .I2 (g12332));
ND3X1 gate18164(.O (g19589), .I1 (g15969), .I2 (g10841), .I3 (g10884));
ND2X1 gate18165(.O (I12277), .I1 (g1467), .I2 (g1472));
ND2X1 gate18166(.O (I13499), .I1 (g232), .I2 (I13497));
ND2X1 gate18167(.O (I17884), .I1 (g13336), .I2 (I17883));
ND2X1 gate18168(.O (g15021), .I1 (g12711), .I2 (g10341));
ND2X1 gate18169(.O (I12075), .I1 (g996), .I2 (I12074));
ND2X1 gate18170(.O (g27365), .I1 (I26050), .I2 (I26051));
ND2X1 gate18171(.O (g24802), .I1 (I23970), .I2 (I23971));
ND2X1 gate18172(.O (g29186), .I1 (g27051), .I2 (g4507));
ND2X1 gate18173(.O (g29676), .I1 (g28381), .I2 (g13676));
ND3X1 gate18174(.O (g7690), .I1 (g4669), .I2 (g4659), .I3 (g4653));
ND4X1 gate18175(.O (g15726), .I1 (g6263), .I2 (g14529), .I3 (g6365), .I4 (g10003));
ND2X1 gate18176(.O (I13498), .I1 (g255), .I2 (I13497));
ND2X1 gate18177(.O (g24793), .I1 (g3742), .I2 (g23124));
ND2X1 gate18178(.O (g26235), .I1 (g8016), .I2 (g24766));
ND2X1 gate18179(.O (g14058), .I1 (g7121), .I2 (g11537));
ND2X1 gate18180(.O (I26440), .I1 (g14271), .I2 (I26438));
ND2X1 gate18181(.O (g28895), .I1 (g27775), .I2 (g8146));
ND2X1 gate18182(.O (I14885), .I1 (g5489), .I2 (I14883));
ND2X1 gate18183(.O (g11881), .I1 (g9060), .I2 (g3361));
ND2X1 gate18184(.O (I14854), .I1 (g9433), .I2 (I14853));
ND2X1 gate18185(.O (g25400), .I1 (g22472), .I2 (g12086));
ND2X1 gate18186(.O (g12225), .I1 (g8324), .I2 (g2453));
ND2X1 gate18187(.O (g14902), .I1 (g7791), .I2 (g12581));
ND2X1 gate18188(.O (g12471), .I1 (I15288), .I2 (I15289));
ND2X1 gate18189(.O (I29303), .I1 (g29496), .I2 (I29302));
ND2X1 gate18190(.O (g12087), .I1 (g7431), .I2 (g2599));
ND2X1 gate18191(.O (g14120), .I1 (g11780), .I2 (g4907));
ND4X1 gate18192(.O (g14739), .I1 (g5929), .I2 (g12067), .I3 (g5983), .I4 (g12351));
ND2X1 gate18193(.O (g10738), .I1 (g6961), .I2 (g10308));
ND2X1 gate18194(.O (I22922), .I1 (g14677), .I2 (I22921));
ND2X1 gate18195(.O (I25845), .I1 (g26212), .I2 (g24799));
ND2X1 gate18196(.O (g14146), .I1 (g11020), .I2 (g691));
ND2X1 gate18197(.O (g32072), .I1 (g31009), .I2 (g13301));
ND2X1 gate18198(.O (g19466), .I1 (g11562), .I2 (g17794));
ND2X1 gate18199(.O (I15003), .I1 (g9691), .I2 (I15002));
ND2X1 gate18200(.O (g12244), .I1 (g7343), .I2 (g5320));
ND3X1 gate18201(.O (g13248), .I1 (g9985), .I2 (g12399), .I3 (g9843));
ND2X1 gate18202(.O (I14480), .I1 (g10074), .I2 (g655));
ND2X1 gate18203(.O (g28376), .I1 (g27064), .I2 (g13620));
ND2X1 gate18204(.O (g13779), .I1 (g11804), .I2 (g11283));
ND2X1 gate18205(.O (I22685), .I1 (g21434), .I2 (I22683));
ND2X1 gate18206(.O (g27955), .I1 (I26460), .I2 (I26461));
ND2X1 gate18207(.O (g28980), .I1 (g27933), .I2 (g14680));
ND2X1 gate18208(.O (I23987), .I1 (g482), .I2 (I23985));
ND2X1 gate18209(.O (g23719), .I1 (I22845), .I2 (I22846));
ND2X1 gate18210(.O (I12401), .I1 (g3808), .I2 (g3813));
ND2X1 gate18211(.O (g28888), .I1 (g27738), .I2 (g8139));
ND3X1 gate18212(.O (g28824), .I1 (g27779), .I2 (g7356), .I3 (g1772));
ND2X1 gate18213(.O (I20488), .I1 (g16757), .I2 (I20486));
ND2X1 gate18214(.O (I22800), .I1 (g11960), .I2 (I22799));
ND2X1 gate18215(.O (I22936), .I1 (g12226), .I2 (g21228));
ND2X1 gate18216(.O (g11356), .I1 (g9552), .I2 (g3632));
ND4X1 gate18217(.O (g8691), .I1 (g3267), .I2 (g3310), .I3 (g3281), .I4 (g3303));
ND2X1 gate18218(.O (g13945), .I1 (g691), .I2 (g11740));
ND3X1 gate18219(.O (g19874), .I1 (g13665), .I2 (g16299), .I3 (g8163));
ND4X1 gate18220(.O (g17581), .I1 (g5607), .I2 (g12029), .I3 (g5623), .I4 (g14669));
ND3X1 gate18221(.O (g17315), .I1 (g9564), .I2 (g9516), .I3 (g14503));
ND3X1 gate18222(.O (g28931), .I1 (g27886), .I2 (g2070), .I3 (g1996));
ND2X1 gate18223(.O (I23969), .I1 (g22202), .I2 (g490));
ND2X1 gate18224(.O (g14547), .I1 (g9439), .I2 (g12201));
ND2X1 gate18225(.O (g14895), .I1 (g7766), .I2 (g12571));
ND2X1 gate18226(.O (g11998), .I1 (g8324), .I2 (g8373));
ND2X1 gate18227(.O (I22762), .I1 (g21434), .I2 (I22760));
ND2X1 gate18228(.O (g13672), .I1 (g8933), .I2 (g11261));
ND2X1 gate18229(.O (g12459), .I1 (g7437), .I2 (g5623));
ND4X1 gate18230(.O (g16663), .I1 (g13854), .I2 (g13834), .I3 (g14655), .I4 (g12292));
ND2X1 gate18231(.O (g10551), .I1 (g1728), .I2 (g7356));
ND2X1 gate18232(.O (g21388), .I1 (g11608), .I2 (g17157));
ND3X1 gate18233(.O (g24880), .I1 (g23281), .I2 (g23266), .I3 (g22839));
ND2X1 gate18234(.O (g23324), .I1 (g703), .I2 (g20181));
ND2X1 gate18235(.O (g14572), .I1 (g12169), .I2 (g9678));
ND2X1 gate18236(.O (I14734), .I1 (g9732), .I2 (I14733));
ND2X1 gate18237(.O (I20189), .I1 (g1333), .I2 (I20187));
ND2X1 gate18238(.O (g21272), .I1 (g11268), .I2 (g17157));
ND2X1 gate18239(.O (I13043), .I1 (g5115), .I2 (g5120));
ND2X1 gate18240(.O (I14993), .I1 (g6527), .I2 (I14991));
ND2X1 gate18241(.O (I20188), .I1 (g16272), .I2 (I20187));
ND3X1 gate18242(.O (g13513), .I1 (g1351), .I2 (g11815), .I3 (g8002));
ND2X1 gate18243(.O (g14127), .I1 (g11653), .I2 (g11435));
ND4X1 gate18244(.O (g21462), .I1 (g17816), .I2 (g14871), .I3 (g17779), .I4 (g14829));
ND2X1 gate18245(.O (g11961), .I1 (g9777), .I2 (g5105));
ND2X1 gate18246(.O (g12079), .I1 (g1792), .I2 (g8195));
ND2X1 gate18247(.O (g28860), .I1 (g27775), .I2 (g14586));
ND4X1 gate18248(.O (g13897), .I1 (g3211), .I2 (g11217), .I3 (g3329), .I4 (g11519));
ND2X1 gate18249(.O (I20460), .I1 (g17515), .I2 (g14187));
ND2X1 gate18250(.O (I24383), .I1 (g23721), .I2 (g14347));
ND2X1 gate18251(.O (g12078), .I1 (g8187), .I2 (g8093));
ND2X1 gate18252(.O (I26071), .I1 (g26026), .I2 (I26070));
ND2X1 gate18253(.O (I15212), .I1 (g10035), .I2 (g1714));
ND2X1 gate18254(.O (g14956), .I1 (g12604), .I2 (g10281));
ND2X1 gate18255(.O (I11879), .I1 (g4430), .I2 (I11877));
ND2X1 gate18256(.O (g14889), .I1 (g12609), .I2 (g12824));
ND4X1 gate18257(.O (g16757), .I1 (g13911), .I2 (g13886), .I3 (g14120), .I4 (g11675));
ND2X1 gate18258(.O (I11878), .I1 (g4388), .I2 (I11877));
ND3X1 gate18259(.O (g28987), .I1 (g27886), .I2 (g2070), .I3 (g7411));
ND3X1 gate18260(.O (g25435), .I1 (g22432), .I2 (g2342), .I3 (g8316));
ND2X1 gate18261(.O (I23979), .I1 (g23198), .I2 (I23978));
ND2X1 gate18262(.O (g24989), .I1 (g21345), .I2 (g23363));
ND2X1 gate18263(.O (g12159), .I1 (g8765), .I2 (g4864));
ND2X1 gate18264(.O (g12125), .I1 (g9728), .I2 (g5101));
ND2X1 gate18265(.O (I21978), .I1 (g19620), .I2 (I21976));
ND2X1 gate18266(.O (I22974), .I1 (g19638), .I2 (I22972));
ND2X1 gate18267(.O (I23978), .I1 (g23198), .I2 (g13670));
ND2X1 gate18268(.O (g24988), .I1 (g546), .I2 (g23088));
ND2X1 gate18269(.O (g24924), .I1 (g20007), .I2 (g23172));
ND2X1 gate18270(.O (I15149), .I1 (g5659), .I2 (I15147));
ND2X1 gate18271(.O (g21360), .I1 (g11510), .I2 (g17157));
ND2X1 gate18272(.O (I23986), .I1 (g22182), .I2 (I23985));
ND2X1 gate18273(.O (g27295), .I1 (g24776), .I2 (g26208));
ND4X1 gate18274(.O (g20271), .I1 (g16925), .I2 (g14054), .I3 (g16657), .I4 (g16628));
ND2X1 gate18275(.O (g11149), .I1 (g1564), .I2 (g7948));
ND2X1 gate18276(.O (I15148), .I1 (g9864), .I2 (I15147));
ND2X1 gate18277(.O (g28969), .I1 (g27854), .I2 (g8267));
ND2X1 gate18278(.O (I26367), .I1 (g26400), .I2 (I26366));
ND2X1 gate18279(.O (I26394), .I1 (g26488), .I2 (I26393));
ND2X1 gate18280(.O (g12144), .I1 (I15003), .I2 (I15004));
ND2X1 gate18281(.O (g9543), .I1 (g2217), .I2 (g2185));
ND4X1 gate18282(.O (g13097), .I1 (g5204), .I2 (g12002), .I3 (g5339), .I4 (g9780));
ND2X1 gate18283(.O (g10520), .I1 (g7195), .I2 (g7115));
ND2X1 gate18284(.O (g13104), .I1 (g1404), .I2 (g10794));
ND2X1 gate18285(.O (g12336), .I1 (I15175), .I2 (I15176));
ND2X1 gate18286(.O (g14520), .I1 (g9369), .I2 (g12163));
ND2X1 gate18287(.O (I14187), .I1 (g3470), .I2 (I14185));
ND2X1 gate18288(.O (g7150), .I1 (g5016), .I2 (g5062));
ND2X1 gate18289(.O (I25220), .I1 (g482), .I2 (I25219));
ND4X1 gate18290(.O (g20199), .I1 (g16815), .I2 (g13968), .I3 (g16749), .I4 (g13907));
ND2X1 gate18291(.O (g11971), .I1 (g8249), .I2 (g8302));
ND2X1 gate18292(.O (g28870), .I1 (g27796), .I2 (g14588));
ND3X1 gate18293(.O (g34048), .I1 (g33669), .I2 (g10583), .I3 (g7442));
ND2X1 gate18294(.O (I13079), .I1 (g5467), .I2 (I13077));
ND2X1 gate18295(.O (I13444), .I1 (g239), .I2 (I13442));
ND2X1 gate18296(.O (I32432), .I1 (g34056), .I2 (I32431));
ND2X1 gate18297(.O (g14546), .I1 (g12125), .I2 (g9613));
ND2X1 gate18298(.O (g14089), .I1 (g11755), .I2 (g4717));
ND2X1 gate18299(.O (g22688), .I1 (g20219), .I2 (g2936));
ND4X1 gate18300(.O (g20198), .I1 (g16813), .I2 (g13958), .I3 (g16745), .I4 (g13927));
ND4X1 gate18301(.O (g17706), .I1 (g3921), .I2 (g11255), .I3 (g3983), .I4 (g13933));
ND4X1 gate18302(.O (g17597), .I1 (g3191), .I2 (g13700), .I3 (g3303), .I4 (g8481));
ND2X1 gate18303(.O (I12074), .I1 (g996), .I2 (g979));
ND2X1 gate18304(.O (I13078), .I1 (g5462), .I2 (I13077));
ND4X1 gate18305(.O (g14088), .I1 (g3901), .I2 (g11255), .I3 (g4000), .I4 (g11631));
ND2X1 gate18306(.O (g14024), .I1 (g7121), .I2 (g11763));
ND4X1 gate18307(.O (g17689), .I1 (g6645), .I2 (g12137), .I3 (g6661), .I4 (g14786));
ND2X1 gate18308(.O (I18589), .I1 (g14679), .I2 (I18587));
ND2X1 gate18309(.O (g24528), .I1 (g4098), .I2 (g22654));
ND2X1 gate18310(.O (g17624), .I1 (I18588), .I2 (I18589));
ND3X1 gate18311(.O (g28867), .I1 (g27800), .I2 (g2227), .I3 (g2153));
ND2X1 gate18312(.O (I18588), .I1 (g2370), .I2 (I18587));
ND2X1 gate18313(.O (g7836), .I1 (g4653), .I2 (g4688));
ND2X1 gate18314(.O (I20467), .I1 (g16663), .I2 (g16728));
ND2X1 gate18315(.O (I14169), .I1 (g8389), .I2 (g3119));
ND2X1 gate18316(.O (I14884), .I1 (g9500), .I2 (I14883));
ND3X1 gate18317(.O (g11412), .I1 (g8666), .I2 (g6918), .I3 (g8697));
ND2X1 gate18318(.O (g15702), .I1 (g13066), .I2 (g7293));
ND2X1 gate18319(.O (g13850), .I1 (g11279), .I2 (g8396));
ND2X1 gate18320(.O (g15904), .I1 (I17380), .I2 (I17381));
ND2X1 gate18321(.O (g25049), .I1 (g21344), .I2 (g23462));
ND3X1 gate18322(.O (g12289), .I1 (g9978), .I2 (g9766), .I3 (g9708));
ND2X1 gate18323(.O (g14659), .I1 (g12646), .I2 (g12443));
ND4X1 gate18324(.O (g14625), .I1 (g3897), .I2 (g11225), .I3 (g4031), .I4 (g8595));
ND4X1 gate18325(.O (g14987), .I1 (g6593), .I2 (g12211), .I3 (g6692), .I4 (g12721));
ND4X1 gate18326(.O (g20161), .I1 (g17732), .I2 (g17706), .I3 (g17670), .I4 (g14625));
ND2X1 gate18327(.O (g22885), .I1 (g9104), .I2 (g20154));
ND2X1 gate18328(.O (g12023), .I1 (g2453), .I2 (g8373));
ND2X1 gate18329(.O (g28910), .I1 (g27854), .I2 (g14614));
ND4X1 gate18330(.O (g13896), .I1 (g3227), .I2 (g11194), .I3 (g3281), .I4 (g11350));
ND2X1 gate18331(.O (I23917), .I1 (g23975), .I2 (g9333));
ND2X1 gate18332(.O (g25048), .I1 (g542), .I2 (g23088));
ND2X1 gate18333(.O (g12224), .I1 (I15088), .I2 (I15089));
ND2X1 gate18334(.O (g14943), .I1 (g7791), .I2 (g12622));
ND2X1 gate18335(.O (I13336), .I1 (g1691), .I2 (I13334));
ND2X1 gate18336(.O (g27687), .I1 (g25200), .I2 (g26714));
ND2X1 gate18337(.O (g14968), .I1 (g12739), .I2 (g10312));
ND2X1 gate18338(.O (g11959), .I1 (g8316), .I2 (g2342));
ND2X1 gate18339(.O (g13627), .I1 (g11172), .I2 (g8388));
ND2X1 gate18340(.O (I22684), .I1 (g11893), .I2 (I22683));
ND2X1 gate18341(.O (I20167), .I1 (g990), .I2 (I20165));
ND2X1 gate18342(.O (g14855), .I1 (g12700), .I2 (g12824));
ND2X1 gate18343(.O (I12729), .I1 (g4291), .I2 (I12728));
ND4X1 gate18344(.O (g13050), .I1 (g5543), .I2 (g12029), .I3 (g5654), .I4 (g9864));
ND4X1 gate18345(.O (g13958), .I1 (g3610), .I2 (g11238), .I3 (g3618), .I4 (g11389));
ND2X1 gate18346(.O (I12728), .I1 (g4291), .I2 (g4287));
ND3X1 gate18347(.O (g28877), .I1 (g27937), .I2 (g7490), .I3 (g7431));
ND2X1 gate18348(.O (g20068), .I1 (g11293), .I2 (g17794));
ND2X1 gate18349(.O (I26366), .I1 (g26400), .I2 (g14211));
ND2X1 gate18350(.O (I14531), .I1 (g8840), .I2 (I14530));
ND2X1 gate18351(.O (g13742), .I1 (g11780), .I2 (g11283));
ND2X1 gate18352(.O (g11944), .I1 (I14765), .I2 (I14766));
ND2X1 gate18353(.O (g7620), .I1 (I12097), .I2 (I12098));
ND2X1 gate18354(.O (g8010), .I1 (I12345), .I2 (I12346));
ND2X1 gate18355(.O (I14186), .I1 (g8442), .I2 (I14185));
ND2X1 gate18356(.O (g17287), .I1 (g7262), .I2 (g14228));
ND2X1 gate18357(.O (g12195), .I1 (g2619), .I2 (g8381));
ND2X1 gate18358(.O (g17596), .I1 (g8686), .I2 (g14367));
ND2X1 gate18359(.O (g25514), .I1 (g12540), .I2 (g22498));
ND2X1 gate18360(.O (g24792), .I1 (I23950), .I2 (I23951));
ND2X1 gate18361(.O (g17243), .I1 (g7247), .I2 (g14212));
ND2X1 gate18362(.O (g12525), .I1 (g7522), .I2 (g6668));
ND2X1 gate18363(.O (g12016), .I1 (g1648), .I2 (g8093));
ND2X1 gate18364(.O (g23281), .I1 (g18957), .I2 (g2898));
ND2X1 gate18365(.O (g21301), .I1 (g11371), .I2 (g17157));
ND2X1 gate18366(.O (g21377), .I1 (g11560), .I2 (g17157));
ND2X1 gate18367(.O (g14055), .I1 (g11697), .I2 (g11763));
ND4X1 gate18368(.O (g17773), .I1 (g5965), .I2 (g14549), .I3 (g5976), .I4 (g9935));
ND2X1 gate18369(.O (I18485), .I1 (g1677), .I2 (g14611));
ND2X1 gate18370(.O (g14978), .I1 (g12716), .I2 (g10491));
ND4X1 gate18371(.O (g15780), .I1 (g5937), .I2 (g14549), .I3 (g6012), .I4 (g14701));
ND2X1 gate18372(.O (I17475), .I1 (g13336), .I2 (I17474));
ND4X1 gate18373(.O (g14590), .I1 (g3546), .I2 (g11207), .I3 (g3680), .I4 (g8542));
ND2X1 gate18374(.O (g24918), .I1 (g136), .I2 (g23088));
ND4X1 gate18375(.O (g17670), .I1 (g3893), .I2 (g13772), .I3 (g4005), .I4 (g8595));
ND2X1 gate18376(.O (g22839), .I1 (g20114), .I2 (g2988));
ND2X1 gate18377(.O (g23699), .I1 (g21012), .I2 (g11160));
ND2X1 gate18378(.O (I29302), .I1 (g29496), .I2 (g12121));
ND2X1 gate18379(.O (g25473), .I1 (g12437), .I2 (g22432));
ND2X1 gate18380(.O (g14741), .I1 (g12711), .I2 (g10421));
ND2X1 gate18381(.O (g27705), .I1 (g25237), .I2 (g26782));
ND2X1 gate18382(.O (g22838), .I1 (g20219), .I2 (g2960));
ND4X1 gate18383(.O (g17734), .I1 (g5272), .I2 (g14490), .I3 (g5283), .I4 (g9780));
ND2X1 gate18384(.O (g28923), .I1 (g27775), .I2 (g8195));
ND3X1 gate18385(.O (g16282), .I1 (g4933), .I2 (g13939), .I3 (g12088));
ND2X1 gate18386(.O (g9442), .I1 (g5424), .I2 (g5428));
ND2X1 gate18387(.O (g27679), .I1 (g25186), .I2 (g26685));
ND2X1 gate18388(.O (I15129), .I1 (g9914), .I2 (I15128));
ND2X1 gate18389(.O (g12042), .I1 (g9086), .I2 (g703));
ND2X1 gate18390(.O (I15002), .I1 (g9691), .I2 (g1700));
ND2X1 gate18391(.O (I26095), .I1 (g13539), .I2 (I26093));
ND2X1 gate18392(.O (g12255), .I1 (g9958), .I2 (g6140));
ND2X1 gate18393(.O (g11002), .I1 (g7475), .I2 (g862));
ND2X1 gate18394(.O (I15128), .I1 (g9914), .I2 (g2527));
ND2X1 gate18395(.O (g13057), .I1 (g969), .I2 (g11294));
ND2X1 gate18396(.O (g14735), .I1 (g12739), .I2 (g12571));
ND2X1 gate18397(.O (g12188), .I1 (g8249), .I2 (g1894));
ND2X1 gate18398(.O (g12124), .I1 (g8741), .I2 (g4674));
ND2X1 gate18399(.O (I13392), .I1 (g1825), .I2 (I13390));
ND3X1 gate18400(.O (g11245), .I1 (g7636), .I2 (g7733), .I3 (g7697));
ND2X1 gate18401(.O (I15299), .I1 (g10112), .I2 (I15298));
ND3X1 gate18402(.O (g12460), .I1 (g10093), .I2 (g5644), .I3 (g5694));
ND3X1 gate18403(.O (g12686), .I1 (g7097), .I2 (g6682), .I3 (g6736));
ND2X1 gate18404(.O (I20166), .I1 (g16246), .I2 (I20165));
ND2X1 gate18405(.O (g11323), .I1 (I14351), .I2 (I14352));
ND4X1 gate18406(.O (g14695), .I1 (g5583), .I2 (g12029), .I3 (g5637), .I4 (g12301));
ND2X1 gate18407(.O (g14018), .I1 (g10323), .I2 (g11483));
ND2X1 gate18408(.O (I15298), .I1 (g10112), .I2 (g1982));
ND3X1 gate18409(.O (g11533), .I1 (g6905), .I2 (g3639), .I3 (g3698));
ND2X1 gate18410(.O (g21403), .I1 (g11652), .I2 (g17157));
ND2X1 gate18411(.O (g20783), .I1 (g14616), .I2 (g17225));
ND3X1 gate18412(.O (g12294), .I1 (g10044), .I2 (g7018), .I3 (g10090));
ND2X1 gate18413(.O (g17618), .I1 (I18580), .I2 (I18581));
ND3X1 gate18414(.O (g28885), .I1 (g27742), .I2 (g1668), .I3 (g7268));
ND4X1 gate18415(.O (g22306), .I1 (g4584), .I2 (g4616), .I3 (g13202), .I4 (g19071));
ND2X1 gate18416(.O (I22873), .I1 (g21228), .I2 (I22871));
ND2X1 gate18417(.O (I11865), .I1 (g4434), .I2 (I11864));
ND2X1 gate18418(.O (I14230), .I1 (g8055), .I2 (I14228));
ND4X1 gate18419(.O (g17468), .I1 (g3215), .I2 (g13700), .I3 (g3317), .I4 (g8481));
ND2X1 gate18420(.O (I21993), .I1 (g7670), .I2 (I21992));
ND4X1 gate18421(.O (g15787), .I1 (g6283), .I2 (g14575), .I3 (g6358), .I4 (g14745));
ND4X1 gate18422(.O (g14706), .I1 (g6287), .I2 (g12101), .I3 (g6369), .I4 (g12672));
ND2X1 gate18423(.O (I14992), .I1 (g9685), .I2 (I14991));
ND4X1 gate18424(.O (g21385), .I1 (g17736), .I2 (g14696), .I3 (g17679), .I4 (g14636));
ND2X1 gate18425(.O (I14510), .I1 (g8721), .I2 (I14508));
ND4X1 gate18426(.O (g15743), .I1 (g5893), .I2 (g14497), .I3 (g6005), .I4 (g9935));
ND2X1 gate18427(.O (g21354), .I1 (g11468), .I2 (g17157));
ND2X1 gate18428(.O (g14688), .I1 (g12604), .I2 (g12453));
ND3X1 gate18429(.O (g28287), .I1 (g10504), .I2 (g26131), .I3 (g26973));
ND2X1 gate18430(.O (g12915), .I1 (g12806), .I2 (g12632));
ND2X1 gate18431(.O (I13383), .I1 (g269), .I2 (I13382));
ND2X1 gate18432(.O (g11445), .I1 (g9771), .I2 (g3976));
ND2X1 gate18433(.O (g14157), .I1 (g11715), .I2 (g11763));
ND2X1 gate18434(.O (g22666), .I1 (g18957), .I2 (g2878));
ND4X1 gate18435(.O (g13499), .I1 (g11479), .I2 (g11442), .I3 (g11410), .I4 (g11382));
ND2X1 gate18436(.O (I13065), .I1 (g4308), .I2 (g4304));
ND2X1 gate18437(.O (g14066), .I1 (g11514), .I2 (g11473));
ND4X1 gate18438(.O (g13498), .I1 (g12577), .I2 (g12522), .I3 (g12462), .I4 (g12416));
ND2X1 gate18439(.O (I15080), .I1 (g1968), .I2 (I15078));
ND2X1 gate18440(.O (g17363), .I1 (g8635), .I2 (g14367));
ND3X1 gate18441(.O (g28942), .I1 (g27858), .I2 (g2331), .I3 (g7335));
ND2X1 gate18442(.O (g17217), .I1 (g7239), .I2 (g14194));
ND2X1 gate18443(.O (g21190), .I1 (g6077), .I2 (g17420));
ND2X1 gate18444(.O (g14876), .I1 (g12492), .I2 (g12443));
ND2X1 gate18445(.O (g14885), .I1 (g12651), .I2 (g12505));
ND4X1 gate18446(.O (g14854), .I1 (g5555), .I2 (g12093), .I3 (g5654), .I4 (g12563));
ND3X1 gate18447(.O (g10511), .I1 (g4628), .I2 (g7202), .I3 (g4621));
ND2X1 gate18448(.O (g11432), .I1 (g10295), .I2 (g8864));
ND2X1 gate18449(.O (I23601), .I1 (g22360), .I2 (I23600));
ND2X1 gate18450(.O (g13432), .I1 (g4793), .I2 (g10831));
ND2X1 gate18451(.O (I14275), .I1 (g8218), .I2 (g3484));
ND2X1 gate18452(.O (g12155), .I1 (g7753), .I2 (g7717));
ND4X1 gate18453(.O (g12822), .I1 (g6978), .I2 (g7236), .I3 (g7224), .I4 (g7163));
ND2X1 gate18454(.O (g15027), .I1 (g12667), .I2 (g10341));
ND2X1 gate18455(.O (I15342), .I1 (g2541), .I2 (I15340));
ND2X1 gate18456(.O (g28930), .I1 (g27833), .I2 (g8201));
ND2X1 gate18457(.O (I24439), .I1 (g23771), .I2 (I24438));
ND2X1 gate18458(.O (g28965), .I1 (g27882), .I2 (g8255));
ND2X1 gate18459(.O (g30573), .I1 (g29355), .I2 (g19666));
ND2X1 gate18460(.O (I24438), .I1 (g23771), .I2 (g14411));
ND2X1 gate18461(.O (g15710), .I1 (g319), .I2 (g13385));
ND2X1 gate18462(.O (g9715), .I1 (g5011), .I2 (g4836));
ND2X1 gate18463(.O (g28131), .I1 (g27051), .I2 (g25838));
ND3X1 gate18464(.O (g31509), .I1 (g599), .I2 (g29933), .I3 (g12323));
ND2X1 gate18465(.O (g10916), .I1 (g1146), .I2 (g7854));
ND2X1 gate18466(.O (I12241), .I1 (g1111), .I2 (I12240));
ND4X1 gate18467(.O (g33933), .I1 (g33394), .I2 (g12491), .I3 (g12819), .I4 (g12796));
ND2X1 gate18468(.O (g12589), .I1 (g7591), .I2 (g6692));
ND2X1 gate18469(.O (g12194), .I1 (g8373), .I2 (g8273));
ND2X1 gate18470(.O (g10550), .I1 (g7268), .I2 (g7308));
ND4X1 gate18471(.O (g13529), .I1 (g11590), .I2 (g11544), .I3 (g11492), .I4 (g11446));
ND2X1 gate18472(.O (I14517), .I1 (g10147), .I2 (I14516));
ND3X1 gate18473(.O (g12588), .I1 (g10169), .I2 (g6336), .I3 (g6386));
ND2X1 gate18474(.O (g27401), .I1 (I26094), .I2 (I26095));
ND3X1 gate18475(.O (g12524), .I1 (g7074), .I2 (g7087), .I3 (g10212));
ND2X1 gate18476(.O (g23659), .I1 (g9434), .I2 (g20854));
ND2X1 gate18477(.O (g11330), .I1 (g9483), .I2 (g1193));
ND3X1 gate18478(.O (g13528), .I1 (g11294), .I2 (g7549), .I3 (g1008));
ND2X1 gate18479(.O (g13330), .I1 (g4664), .I2 (g11006));
ND2X1 gate18480(.O (g10307), .I1 (I13730), .I2 (I13731));
ND2X1 gate18481(.O (I15365), .I1 (g2675), .I2 (I15363));
ND2X1 gate18482(.O (g14085), .I1 (g7121), .I2 (g11584));
ND4X1 gate18483(.O (g17740), .I1 (g5945), .I2 (g14497), .I3 (g6012), .I4 (g12351));
ND2X1 gate18484(.O (g13764), .I1 (g11252), .I2 (g3072));
ND2X1 gate18485(.O (g8238), .I1 (I12469), .I2 (I12470));
ND4X1 gate18486(.O (g14596), .I1 (g12196), .I2 (g9775), .I3 (g12124), .I4 (g9663));
ND2X1 gate18487(.O (g12119), .I1 (g2351), .I2 (g8267));
ND4X1 gate18488(.O (g14054), .I1 (g3550), .I2 (g11238), .I3 (g3649), .I4 (g11576));
ND2X1 gate18489(.O (I22711), .I1 (g11915), .I2 (I22710));
ND3X1 gate18490(.O (g7701), .I1 (g4859), .I2 (g4849), .I3 (g4843));
ND4X1 gate18491(.O (g21339), .I1 (g15725), .I2 (g13084), .I3 (g15713), .I4 (g13050));
ND2X1 gate18492(.O (g13960), .I1 (g11669), .I2 (g11537));
ND2X1 gate18493(.O (g32057), .I1 (g31003), .I2 (g13297));
ND2X1 gate18494(.O (g12118), .I1 (g8259), .I2 (g8150));
ND2X1 gate18495(.O (g12022), .I1 (g7335), .I2 (g2331));
ND4X1 gate18496(.O (g21338), .I1 (g15741), .I2 (g15734), .I3 (g15728), .I4 (g13097));
ND2X1 gate18497(.O (I26070), .I1 (g26026), .I2 (g13517));
ND2X1 gate18498(.O (I17474), .I1 (g13336), .I2 (g1105));
ND4X1 gate18499(.O (g16723), .I1 (g3606), .I2 (g13730), .I3 (g3676), .I4 (g11576));
ND2X1 gate18500(.O (g14773), .I1 (g12711), .I2 (g12581));
ND3X1 gate18501(.O (g24544), .I1 (g22666), .I2 (g22661), .I3 (g22651));
ND2X1 gate18502(.O (g13709), .I1 (g11755), .I2 (g11261));
ND2X1 gate18503(.O (g25389), .I1 (g22457), .I2 (g12082));
ND2X1 gate18504(.O (g12285), .I1 (I15122), .I2 (I15123));
ND2X1 gate18505(.O (I15087), .I1 (g9832), .I2 (g2393));
ND2X1 gate18506(.O (g14655), .I1 (g4743), .I2 (g11755));
ND2X1 gate18507(.O (g11708), .I1 (g10147), .I2 (g10110));
ND2X1 gate18508(.O (g13708), .I1 (g11200), .I2 (g8507));
ND2X1 gate18509(.O (g12053), .I1 (g2587), .I2 (g8418));
ND2X1 gate18510(.O (g16097), .I1 (g13319), .I2 (g10998));
ND2X1 gate18511(.O (I26094), .I1 (g26055), .I2 (I26093));
ND2X1 gate18512(.O (I24415), .I1 (g23751), .I2 (I24414));
ND2X1 gate18513(.O (I15043), .I1 (g1834), .I2 (I15041));
ND2X1 gate18514(.O (g13043), .I1 (g10521), .I2 (g969));
ND2X1 gate18515(.O (g14930), .I1 (g12609), .I2 (g12515));
ND2X1 gate18516(.O (g14993), .I1 (g12695), .I2 (g12453));
ND2X1 gate18517(.O (I17381), .I1 (g1129), .I2 (I17379));
ND2X1 gate18518(.O (g24678), .I1 (g22994), .I2 (g23010));
ND2X1 gate18519(.O (g14838), .I1 (g12492), .I2 (g12405));
ND2X1 gate18520(.O (g14965), .I1 (g12609), .I2 (g12571));
ND2X1 gate18521(.O (g22908), .I1 (g9104), .I2 (g20175));
ND4X1 gate18522(.O (g13069), .I1 (g5889), .I2 (g12067), .I3 (g6000), .I4 (g9935));
ND2X1 gate18523(.O (g29702), .I1 (g28395), .I2 (g13712));
ND3X1 gate18524(.O (g34162), .I1 (g785), .I2 (g33823), .I3 (g11679));
ND2X1 gate18525(.O (g15717), .I1 (g10754), .I2 (g13092));
ND2X1 gate18526(.O (I13401), .I1 (g2246), .I2 (g2250));
ND2X1 gate18527(.O (g11955), .I1 (g8302), .I2 (g1917));
ND2X1 gate18528(.O (g13955), .I1 (g11621), .I2 (g11527));
ND2X1 gate18529(.O (g11970), .I1 (g1760), .I2 (g8241));
ND2X1 gate18530(.O (g28410), .I1 (g27074), .I2 (g13679));
ND2X1 gate18531(.O (g19962), .I1 (g11470), .I2 (g17794));
ND2X1 gate18532(.O (g10618), .I1 (g10153), .I2 (g9913));
ND2X1 gate18533(.O (I14351), .I1 (g8890), .I2 (I14350));
ND2X1 gate18534(.O (g27693), .I1 (g25216), .I2 (g26752));
ND2X1 gate18535(.O (I11864), .I1 (g4434), .I2 (g4401));
ND2X1 gate18536(.O (g34220), .I1 (I32186), .I2 (I32187));
ND2X1 gate18537(.O (g28363), .I1 (g27064), .I2 (g13593));
ND2X1 gate18538(.O (g17568), .I1 (I18486), .I2 (I18487));
ND2X1 gate18539(.O (g14279), .I1 (g12111), .I2 (g9246));
ND2X1 gate18540(.O (g7887), .I1 (I12278), .I2 (I12279));
ND2X1 gate18541(.O (I13749), .I1 (g4608), .I2 (g4584));
ND2X1 gate18542(.O (g13886), .I1 (g11804), .I2 (g4922));
ND2X1 gate18543(.O (g7228), .I1 (g6398), .I2 (g6444));
ND2X1 gate18544(.O (g11994), .I1 (g8310), .I2 (g8365));
ND2X1 gate18545(.O (g15723), .I1 (g10775), .I2 (g13104));
ND3X1 gate18546(.O (g23978), .I1 (g572), .I2 (g21389), .I3 (g12323));
ND4X1 gate18547(.O (g13967), .I1 (g3929), .I2 (g11225), .I3 (g3983), .I4 (g11419));
ND2X1 gate18548(.O (I12345), .I1 (g3106), .I2 (I12344));
ND2X1 gate18549(.O (I14790), .I1 (g6167), .I2 (I14788));
ND2X1 gate18550(.O (I14516), .I1 (g10147), .I2 (g661));
ND2X1 gate18551(.O (g23590), .I1 (g20682), .I2 (g11111));
ND2X1 gate18552(.O (I12849), .I1 (g4281), .I2 (I12848));
ND2X1 gate18553(.O (g12008), .I1 (g9932), .I2 (g5798));
ND4X1 gate18554(.O (g17814), .I1 (g5579), .I2 (g14522), .I3 (g5673), .I4 (g12563));
ND2X1 gate18555(.O (g22638), .I1 (g18957), .I2 (g2886));
ND2X1 gate18556(.O (I12848), .I1 (g4281), .I2 (g4277));
ND2X1 gate18557(.O (g12476), .I1 (g7498), .I2 (g6704));
ND3X1 gate18558(.O (g13459), .I1 (g7479), .I2 (g11294), .I3 (g11846));
ND4X1 gate18559(.O (g21384), .I1 (g17734), .I2 (g14686), .I3 (g17675), .I4 (g14663));
ND2X1 gate18560(.O (I23587), .I1 (g4332), .I2 (I23585));
ND2X1 gate18561(.O (g8889), .I1 (g3684), .I2 (g4871));
ND2X1 gate18562(.O (g14038), .I1 (g11514), .I2 (g11435));
ND2X1 gate18563(.O (g23067), .I1 (g20887), .I2 (g10721));
ND2X1 gate18564(.O (g10601), .I1 (g896), .I2 (g7397));
ND4X1 gate18565(.O (g13918), .I1 (g3259), .I2 (g11217), .I3 (g3267), .I4 (g11350));
ND4X1 gate18566(.O (g16925), .I1 (g3574), .I2 (g13799), .I3 (g3668), .I4 (g11576));
ND2X1 gate18567(.O (g14601), .I1 (g12318), .I2 (g6466));
ND2X1 gate18568(.O (I18538), .I1 (g14642), .I2 (I18536));
ND2X1 gate18569(.O (g8871), .I1 (I12841), .I2 (I12842));
ND2X1 gate18570(.O (I15079), .I1 (g9827), .I2 (I15078));
ND2X1 gate18571(.O (g14677), .I1 (I16779), .I2 (I16780));
ND2X1 gate18572(.O (I12263), .I1 (g1448), .I2 (I12261));
ND2X1 gate18573(.O (g11545), .I1 (I14498), .I2 (I14499));
ND3X1 gate18574(.O (g11444), .I1 (g6905), .I2 (g6918), .I3 (g8733));
ND2X1 gate18575(.O (g13079), .I1 (g1312), .I2 (g11336));
ND2X1 gate18576(.O (I15078), .I1 (g9827), .I2 (g1968));
ND2X1 gate18577(.O (g12239), .I1 (I15106), .I2 (I15107));
ND2X1 gate18578(.O (g20201), .I1 (I20468), .I2 (I20469));
ND2X1 gate18579(.O (g8500), .I1 (g3431), .I2 (g3423));
ND2X1 gate18580(.O (g14937), .I1 (g12667), .I2 (g10421));
ND2X1 gate18581(.O (g26025), .I1 (g22405), .I2 (g24631));
ND4X1 gate18582(.O (g13086), .I1 (g6235), .I2 (g12101), .I3 (g6346), .I4 (g10003));
ND2X1 gate18583(.O (g16681), .I1 (I17884), .I2 (I17885));
ND4X1 gate18584(.O (g17578), .I1 (g5212), .I2 (g14399), .I3 (g5283), .I4 (g12497));
ND2X1 gate18585(.O (g12941), .I1 (g7167), .I2 (g10537));
ND2X1 gate18586(.O (g19795), .I1 (g13600), .I2 (g16275));
ND2X1 gate18587(.O (g12185), .I1 (g9905), .I2 (g799));
ND4X1 gate18588(.O (g21402), .I1 (g17757), .I2 (g14740), .I3 (g17716), .I4 (g14674));
ND2X1 gate18589(.O (g17586), .I1 (g14638), .I2 (g14601));
ND2X1 gate18590(.O (g11977), .I1 (g8373), .I2 (g2476));
ND2X1 gate18591(.O (g13977), .I1 (g11610), .I2 (g11729));
ND2X1 gate18592(.O (I14530), .I1 (g8840), .I2 (g8873));
ND2X1 gate18593(.O (g8737), .I1 (I12729), .I2 (I12730));
ND2X1 gate18594(.O (g15011), .I1 (g12716), .I2 (g12632));
ND2X1 gate18595(.O (g34227), .I1 (I32203), .I2 (I32204));
ND2X1 gate18596(.O (g14015), .I1 (g11658), .I2 (g11747));
ND2X1 gate18597(.O (g11561), .I1 (I14517), .I2 (I14518));
ND2X1 gate18598(.O (g25172), .I1 (g5052), .I2 (g23560));
ND2X1 gate18599(.O (I22872), .I1 (g12150), .I2 (I22871));
ND2X1 gate18600(.O (g25996), .I1 (g24601), .I2 (g22838));
ND4X1 gate18601(.O (g20170), .I1 (g16741), .I2 (g13897), .I3 (g16687), .I4 (g13866));
ND2X1 gate18602(.O (g10556), .I1 (g7971), .I2 (g8133));
ND2X1 gate18603(.O (g13823), .I1 (g11313), .I2 (g3774));
ND2X1 gate18604(.O (I13454), .I1 (g1959), .I2 (I13452));
ND2X1 gate18605(.O (I21992), .I1 (g7670), .I2 (g19638));
ND2X1 gate18606(.O (g14223), .I1 (g9092), .I2 (g11858));
ND2X1 gate18607(.O (g17493), .I1 (g8659), .I2 (g14367));
ND2X1 gate18608(.O (g15959), .I1 (I17405), .I2 (I17406));
ND4X1 gate18609(.O (g27577), .I1 (g25019), .I2 (g25002), .I3 (g24988), .I4 (g25765));
ND2X1 gate18610(.O (I15364), .I1 (g10182), .I2 (I15363));
ND3X1 gate18611(.O (g12577), .I1 (g7051), .I2 (g5990), .I3 (g6044));
ND2X1 gate18612(.O (g14110), .I1 (g11692), .I2 (g8906));
ND2X1 gate18613(.O (g9246), .I1 (g847), .I2 (g812));
ND4X1 gate18614(.O (g15742), .I1 (g5575), .I2 (g12093), .I3 (g5637), .I4 (g14669));
ND2X1 gate18615(.O (I23586), .I1 (g22409), .I2 (I23585));
ND2X1 gate18616(.O (g9203), .I1 (g3706), .I2 (g3752));
ND4X1 gate18617(.O (g14740), .I1 (g5913), .I2 (g12129), .I3 (g6031), .I4 (g12614));
ND2X1 gate18618(.O (I13382), .I1 (g269), .I2 (g246));
ND2X1 gate18619(.O (I15289), .I1 (g6697), .I2 (I15287));
ND2X1 gate18620(.O (g19358), .I1 (g15723), .I2 (g1399));
ND2X1 gate18621(.O (I13519), .I1 (g2514), .I2 (I13518));
ND3X1 gate18622(.O (g16299), .I1 (g8160), .I2 (g8112), .I3 (g13706));
ND3X1 gate18623(.O (g31003), .I1 (g27163), .I2 (g29497), .I3 (g19644));
ND2X1 gate18624(.O (g14953), .I1 (g12646), .I2 (g12405));
ND2X1 gate18625(.O (I15288), .I1 (g10061), .I2 (I15287));
ND2X1 gate18626(.O (I13518), .I1 (g2514), .I2 (g2518));
ND2X1 gate18627(.O (g12083), .I1 (g2217), .I2 (g8205));
ND2X1 gate18628(.O (I15308), .I1 (g2407), .I2 (I15306));
ND2X1 gate18629(.O (g11224), .I1 (I14290), .I2 (I14291));
ND2X1 gate18630(.O (g13288), .I1 (g10946), .I2 (g1442));
ND4X1 gate18631(.O (g15730), .I1 (g6609), .I2 (g14556), .I3 (g6711), .I4 (g10061));
ND2X1 gate18632(.O (g14800), .I1 (g7704), .I2 (g12443));
ND2X1 gate18633(.O (I24414), .I1 (g23751), .I2 (g14382));
ND2X1 gate18634(.O (g29046), .I1 (g27779), .I2 (g9640));
ND3X1 gate18635(.O (g13495), .I1 (g1008), .I2 (g11786), .I3 (g7972));
ND2X1 gate18636(.O (I29261), .I1 (g29485), .I2 (g12046));
ND2X1 gate18637(.O (g24809), .I1 (g19965), .I2 (g23132));
ND2X1 gate18638(.O (I22846), .I1 (g21228), .I2 (I22844));
ND2X1 gate18639(.O (g24808), .I1 (I23986), .I2 (I23987));
ND2X1 gate18640(.O (I13729), .I1 (g4534), .I2 (g4537));
ND2X1 gate18641(.O (g10587), .I1 (g2421), .I2 (g7456));
ND2X1 gate18642(.O (g11374), .I1 (g9536), .I2 (g1536));
ND2X1 gate18643(.O (g28391), .I1 (g27064), .I2 (g13637));
ND2X1 gate18644(.O (g12415), .I1 (g7496), .I2 (g5976));
ND2X1 gate18645(.O (g21287), .I1 (g14616), .I2 (g17571));
ND2X1 gate18646(.O (g19506), .I1 (g4087), .I2 (g15825));
ND2X1 gate18647(.O (g10909), .I1 (g7304), .I2 (g1116));
ND3X1 gate18648(.O (g20733), .I1 (g14406), .I2 (g17290), .I3 (g9509));
ND4X1 gate18649(.O (g21307), .I1 (g15719), .I2 (g13067), .I3 (g15709), .I4 (g13040));
ND2X1 gate18650(.O (g15002), .I1 (g12609), .I2 (g10312));
ND2X1 gate18651(.O (I25243), .I1 (g490), .I2 (I25242));
ND2X1 gate18652(.O (g13260), .I1 (g1116), .I2 (g10666));
ND2X1 gate18653(.O (g14908), .I1 (g7812), .I2 (g10491));
ND2X1 gate18654(.O (g10569), .I1 (g2287), .I2 (g7418));
ND2X1 gate18655(.O (I22929), .I1 (g12223), .I2 (g21228));
ND2X1 gate18656(.O (I15195), .I1 (g6005), .I2 (I15193));
ND2X1 gate18657(.O (I17405), .I1 (g13378), .I2 (I17404));
ND2X1 gate18658(.O (I12344), .I1 (g3106), .I2 (g3111));
ND4X1 gate18659(.O (g14569), .I1 (g3195), .I2 (g11194), .I3 (g3329), .I4 (g8481));
ND2X1 gate18660(.O (g11489), .I1 (g9661), .I2 (g3618));
ND2X1 gate18661(.O (g10568), .I1 (g7328), .I2 (g7374));
ND2X1 gate18662(.O (g25895), .I1 (g1259), .I2 (g24453));
ND2X1 gate18663(.O (g16316), .I1 (g9429), .I2 (g13518));
ND2X1 gate18664(.O (g11559), .I1 (I14509), .I2 (I14510));
ND2X1 gate18665(.O (g11424), .I1 (g9662), .I2 (g4012));
ND2X1 gate18666(.O (I13566), .I1 (g2652), .I2 (I13564));
ND2X1 gate18667(.O (g23655), .I1 (I22793), .I2 (I22794));
ND2X1 gate18668(.O (I29271), .I1 (g12050), .I2 (I29269));
ND2X1 gate18669(.O (g9883), .I1 (g5782), .I2 (g5774));
ND2X1 gate18670(.O (g14123), .I1 (g10685), .I2 (g10928));
ND4X1 gate18671(.O (g15737), .I1 (g13240), .I2 (g13115), .I3 (g7903), .I4 (g13210));
ND2X1 gate18672(.O (g14807), .I1 (g7738), .I2 (g12453));
ND3X1 gate18673(.O (g19903), .I1 (g13707), .I2 (g16319), .I3 (g8227));
ND2X1 gate18674(.O (g12115), .I1 (g1926), .I2 (g8249));
ND2X1 gate18675(.O (g14974), .I1 (g12744), .I2 (g12622));
ND4X1 gate18676(.O (g17790), .I1 (g6311), .I2 (g14575), .I3 (g6322), .I4 (g10003));
ND3X1 gate18677(.O (g17137), .I1 (g13727), .I2 (g13511), .I3 (g13527));
ND2X1 gate18678(.O (I13139), .I1 (g6154), .I2 (g6159));
ND3X1 gate18679(.O (g11544), .I1 (g8700), .I2 (g3990), .I3 (g4045));
ND4X1 gate18680(.O (g13544), .I1 (g7972), .I2 (g10521), .I3 (g7549), .I4 (g1008));
ND2X1 gate18681(.O (g24570), .I1 (g22957), .I2 (g2941));
ND2X1 gate18682(.O (g12052), .I1 (g7387), .I2 (g2465));
ND2X1 gate18683(.O (g14638), .I1 (g9626), .I2 (g12361));
ND2X1 gate18684(.O (I15042), .I1 (g9752), .I2 (I15041));
ND2X1 gate18685(.O (I15255), .I1 (g1848), .I2 (I15253));
ND2X1 gate18686(.O (I13852), .I1 (g7397), .I2 (I13850));
ND2X1 gate18687(.O (g14841), .I1 (g12593), .I2 (g12443));
ND3X1 gate18688(.O (g25385), .I1 (g22369), .I2 (g1783), .I3 (g8241));
ND2X1 gate18689(.O (g24567), .I1 (g22957), .I2 (g2917));
ND2X1 gate18690(.O (g11189), .I1 (I14248), .I2 (I14249));
ND2X1 gate18691(.O (g11679), .I1 (g8836), .I2 (g802));
ND2X1 gate18692(.O (I23600), .I1 (g22360), .I2 (g4322));
ND3X1 gate18693(.O (g29778), .I1 (g294), .I2 (g28444), .I3 (g23204));
ND4X1 gate18694(.O (g13124), .I1 (g10666), .I2 (g7661), .I3 (g979), .I4 (g1061));
ND2X1 gate18695(.O (g25888), .I1 (g914), .I2 (g24439));
ND2X1 gate18696(.O (g31971), .I1 (g30573), .I2 (g10511));
ND2X1 gate18697(.O (g23210), .I1 (g18957), .I2 (g2882));
ND4X1 gate18698(.O (g16696), .I1 (g13871), .I2 (g13855), .I3 (g14682), .I4 (g12340));
ND4X1 gate18699(.O (g20185), .I1 (g16772), .I2 (g13928), .I3 (g16723), .I4 (g13882));
ND2X1 gate18700(.O (g10578), .I1 (g7174), .I2 (g6058));
ND3X1 gate18701(.O (g20675), .I1 (g14377), .I2 (g17246), .I3 (g9442));
ND2X1 gate18702(.O (g20092), .I1 (g11373), .I2 (g17794));
ND4X1 gate18703(.O (g14014), .I1 (g3199), .I2 (g11217), .I3 (g3298), .I4 (g11519));
ND2X1 gate18704(.O (g11938), .I1 (g8259), .I2 (g2208));
ND2X1 gate18705(.O (g10586), .I1 (g7380), .I2 (g7418));
ND4X1 gate18706(.O (g13093), .I1 (g10649), .I2 (g7661), .I3 (g979), .I4 (g1061));
ND2X1 gate18707(.O (g8873), .I1 (I12849), .I2 (I12850));
ND2X1 gate18708(.O (g8632), .I1 (g1514), .I2 (g1500));
ND2X1 gate18709(.O (g9538), .I1 (g1792), .I2 (g1760));
ND2X1 gate18710(.O (I20221), .I1 (g16272), .I2 (g11170));
ND2X1 gate18711(.O (I12240), .I1 (g1111), .I2 (g1105));
ND2X1 gate18712(.O (g9509), .I1 (g5770), .I2 (g5774));
ND2X1 gate18713(.O (g23286), .I1 (g6875), .I2 (g20887));
ND2X1 gate18714(.O (g25426), .I1 (g12371), .I2 (g22369));
ND2X1 gate18715(.O (g29672), .I1 (g28376), .I2 (g13672));
ND2X1 gate18716(.O (g17593), .I1 (I18537), .I2 (I18538));
ND2X1 gate18717(.O (g14116), .I1 (g11697), .I2 (g11584));
ND2X1 gate18718(.O (I32185), .I1 (g33665), .I2 (g33661));
ND2X1 gate18719(.O (I14509), .I1 (g370), .I2 (I14508));
ND2X1 gate18720(.O (g10041), .I1 (I13565), .I2 (I13566));
ND2X1 gate18721(.O (g14720), .I1 (g12593), .I2 (g10266));
ND2X1 gate18722(.O (I32518), .I1 (g34422), .I2 (I32516));
ND3X1 gate18723(.O (g16259), .I1 (g4743), .I2 (g13908), .I3 (g12054));
ND2X1 gate18724(.O (I14508), .I1 (g370), .I2 (g8721));
ND3X1 gate18725(.O (g16225), .I1 (g13544), .I2 (g13528), .I3 (g13043));
ND2X1 gate18726(.O (g14041), .I1 (g11610), .I2 (g11473));
ND2X1 gate18727(.O (g21187), .I1 (g14616), .I2 (g17364));
ND2X1 gate18728(.O (I22710), .I1 (g11915), .I2 (g21434));
ND2X1 gate18729(.O (g12207), .I1 (g9887), .I2 (g5794));
ND2X1 gate18730(.O (g23975), .I1 (I23119), .I2 (I23120));
ND2X1 gate18731(.O (g12539), .I1 (I15341), .I2 (I15342));
ND2X1 gate18732(.O (I24463), .I1 (g14437), .I2 (I24461));
ND4X1 gate18733(.O (g15753), .I1 (g6239), .I2 (g14529), .I3 (g6351), .I4 (g10003));
ND2X1 gate18734(.O (g12538), .I1 (I15334), .I2 (I15335));
ND2X1 gate18735(.O (I12262), .I1 (g1454), .I2 (I12261));
ND2X1 gate18736(.O (I13184), .I1 (g6505), .I2 (I13182));
ND2X1 gate18737(.O (I14213), .I1 (g9295), .I2 (I14211));
ND4X1 gate18738(.O (g15736), .I1 (g6295), .I2 (g14575), .I3 (g6373), .I4 (g10003));
ND4X1 gate18739(.O (g17635), .I1 (g3542), .I2 (g13730), .I3 (g3654), .I4 (g8542));
ND2X1 gate18740(.O (g16069), .I1 (I17447), .I2 (I17448));
ND2X1 gate18741(.O (g13915), .I1 (g11566), .I2 (g11473));
ND2X1 gate18742(.O (I22945), .I1 (g9492), .I2 (I22944));
ND2X1 gate18743(.O (g14142), .I1 (g11715), .I2 (g8958));
ND3X1 gate18744(.O (g33925), .I1 (g33394), .I2 (g4462), .I3 (g4467));
ND4X1 gate18745(.O (g16657), .I1 (g3554), .I2 (g13730), .I3 (g3625), .I4 (g11576));
ND2X1 gate18746(.O (I14205), .I1 (g8508), .I2 (I14204));
ND3X1 gate18747(.O (g15843), .I1 (g7922), .I2 (g7503), .I3 (g13264));
ND4X1 gate18748(.O (g14517), .I1 (g3231), .I2 (g11217), .I3 (g3321), .I4 (g8481));
ND2X1 gate18749(.O (g24906), .I1 (g8743), .I2 (g23088));
ND2X1 gate18750(.O (g26714), .I1 (g9316), .I2 (g25175));
ND2X1 gate18751(.O (g23666), .I1 (g20875), .I2 (g11139));
ND2X1 gate18752(.O (I26417), .I1 (g26519), .I2 (g14247));
ND4X1 gate18753(.O (g21363), .I1 (g17708), .I2 (g14664), .I3 (g17640), .I4 (g14598));
ND2X1 gate18754(.O (I32439), .I1 (g34227), .I2 (g34220));
ND2X1 gate18755(.O (g12100), .I1 (I14956), .I2 (I14957));
ND2X1 gate18756(.O (I17380), .I1 (g13336), .I2 (I17379));
ND2X1 gate18757(.O (g24566), .I1 (g22755), .I2 (g22713));
ND2X1 gate18758(.O (g22711), .I1 (g19581), .I2 (g7888));
ND2X1 gate18759(.O (g14130), .I1 (g11621), .I2 (g8906));
ND2X1 gate18760(.O (I18682), .I1 (g14752), .I2 (I18680));
ND2X1 gate18761(.O (g17474), .I1 (g14547), .I2 (g14521));
ND3X1 gate18762(.O (g28516), .I1 (g10857), .I2 (g26105), .I3 (g27155));
ND2X1 gate18763(.O (g11419), .I1 (I14428), .I2 (I14429));
ND2X1 gate18764(.O (g29097), .I1 (g9700), .I2 (g27858));
ND4X1 gate18765(.O (g15709), .I1 (g5224), .I2 (g14399), .I3 (g5327), .I4 (g9780));
ND4X1 gate18766(.O (g27882), .I1 (g21228), .I2 (g25307), .I3 (g26424), .I4 (g26213));
ND3X1 gate18767(.O (g11155), .I1 (g4776), .I2 (g7892), .I3 (g9030));
ND2X1 gate18768(.O (I14350), .I1 (g8890), .I2 (g8848));
ND2X1 gate18769(.O (g15708), .I1 (g7340), .I2 (g13083));
ND3X1 gate18770(.O (g12414), .I1 (g7028), .I2 (g7041), .I3 (g10165));
ND2X1 gate18771(.O (g13822), .I1 (g8160), .I2 (g11306));
ND3X1 gate18772(.O (g13266), .I1 (g12440), .I2 (g9920), .I3 (g9843));
ND2X1 gate18773(.O (g25527), .I1 (g21294), .I2 (g23462));
ND2X1 gate18774(.O (I12098), .I1 (g1322), .I2 (I12096));
ND2X1 gate18775(.O (g14727), .I1 (g12604), .I2 (g12505));
ND2X1 gate18776(.O (I12251), .I1 (g1124), .I2 (g1129));
ND2X1 gate18777(.O (I22717), .I1 (g11916), .I2 (g21434));
ND2X1 gate18778(.O (g17492), .I1 (g8655), .I2 (g14367));
ND2X1 gate18779(.O (I17448), .I1 (g956), .I2 (I17446));
ND2X1 gate18780(.O (I15167), .I1 (g9904), .I2 (I15166));
ND2X1 gate18781(.O (I15194), .I1 (g9935), .I2 (I15193));
ND2X1 gate18782(.O (I17404), .I1 (g13378), .I2 (g1472));
ND2X1 gate18783(.O (I31985), .I1 (g33648), .I2 (I31983));
ND2X1 gate18784(.O (g21186), .I1 (g14616), .I2 (g17363));
ND2X1 gate18785(.O (g23685), .I1 (I22823), .I2 (I22824));
ND2X1 gate18786(.O (g7223), .I1 (I11878), .I2 (I11879));
ND2X1 gate18787(.O (g14600), .I1 (g9564), .I2 (g12311));
ND4X1 gate18788(.O (g14781), .I1 (g6259), .I2 (g12173), .I3 (g6377), .I4 (g12672));
ND2X1 gate18789(.O (g24576), .I1 (g22957), .I2 (g2902));
ND4X1 gate18790(.O (g13119), .I1 (g6625), .I2 (g12211), .I3 (g6715), .I4 (g10061));
ND2X1 gate18791(.O (g21417), .I1 (g11677), .I2 (g17157));
ND2X1 gate18792(.O (g11118), .I1 (I14170), .I2 (I14171));
ND2X1 gate18793(.O (g12114), .I1 (g8241), .I2 (g8146));
ND4X1 gate18794(.O (g13118), .I1 (g5897), .I2 (g12067), .I3 (g6031), .I4 (g9935));
ND2X1 gate18795(.O (g21334), .I1 (g14616), .I2 (g17596));
ND2X1 gate18796(.O (g24609), .I1 (g22850), .I2 (g22650));
ND2X1 gate18797(.O (g20200), .I1 (I20461), .I2 (I20462));
ND2X1 gate18798(.O (I29295), .I1 (g29495), .I2 (g12117));
ND2X1 gate18799(.O (g22663), .I1 (I21977), .I2 (I21978));
ND3X1 gate18800(.O (g33299), .I1 (g608), .I2 (g32296), .I3 (g12323));
ND2X1 gate18801(.O (g23762), .I1 (I22900), .I2 (I22901));
ND2X1 gate18802(.O (I15053), .I1 (g2259), .I2 (I15051));
ND2X1 gate18803(.O (I15254), .I1 (g10078), .I2 (I15253));
ND2X1 gate18804(.O (g27141), .I1 (I25846), .I2 (I25847));
ND2X1 gate18805(.O (I25909), .I1 (g24782), .I2 (I25907));
ND2X1 gate18806(.O (g24798), .I1 (I23962), .I2 (I23963));
ND4X1 gate18807(.O (g14422), .I1 (g3187), .I2 (g11194), .I3 (g3298), .I4 (g8481));
ND2X1 gate18808(.O (g24973), .I1 (g21272), .I2 (g23462));
ND4X1 gate18809(.O (g20184), .I1 (g16770), .I2 (g13918), .I3 (g16719), .I4 (g13896));
ND2X1 gate18810(.O (g23909), .I1 (g7028), .I2 (g20739));
ND2X1 gate18811(.O (I25908), .I1 (g26256), .I2 (I25907));
ND2X1 gate18812(.O (g22757), .I1 (g20114), .I2 (g7891));
ND2X1 gate18813(.O (g12332), .I1 (I15167), .I2 (I15168));
ND2X1 gate18814(.O (g25019), .I1 (g20055), .I2 (g23172));
ND2X1 gate18815(.O (g25018), .I1 (g20107), .I2 (g23154));
ND2X1 gate18816(.O (I18633), .I1 (g2504), .I2 (g14713));
ND4X1 gate18817(.O (g14542), .I1 (g3582), .I2 (g11238), .I3 (g3672), .I4 (g8542));
ND2X1 gate18818(.O (g14021), .I1 (g11697), .I2 (g8958));
ND2X1 gate18819(.O (g24934), .I1 (g21283), .I2 (g23462));
ND2X1 gate18820(.O (I25242), .I1 (g490), .I2 (g24744));
ND4X1 gate18821(.O (g17757), .I1 (g5909), .I2 (g14549), .I3 (g6005), .I4 (g12614));
ND4X1 gate18822(.O (g10726), .I1 (g7304), .I2 (g7661), .I3 (g979), .I4 (g1061));
ND2X1 gate18823(.O (g23747), .I1 (I22865), .I2 (I22866));
ND3X1 gate18824(.O (g10614), .I1 (g9024), .I2 (g8977), .I3 (g8928));
ND4X1 gate18825(.O (g27833), .I1 (g21228), .I2 (g25282), .I3 (g26424), .I4 (g26190));
ND2X1 gate18826(.O (g12049), .I1 (g2208), .I2 (g8150));
ND2X1 gate18827(.O (g10905), .I1 (g1116), .I2 (g7304));
ND2X1 gate18828(.O (I15166), .I1 (g9904), .I2 (g9823));
ND2X1 gate18829(.O (g14905), .I1 (g12785), .I2 (g7142));
ND2X1 gate18830(.O (g12048), .I1 (g7369), .I2 (g2040));
ND4X1 gate18831(.O (g20214), .I1 (g16854), .I2 (g13993), .I3 (g16776), .I4 (g13967));
ND2X1 gate18832(.O (g28109), .I1 (g27051), .I2 (g25783));
ND2X1 gate18833(.O (g12221), .I1 (I15079), .I2 (I15080));
ND4X1 gate18834(.O (g27613), .I1 (g24942), .I2 (g24933), .I3 (g25048), .I4 (g26871));
ND2X1 gate18835(.O (g11892), .I1 (g7777), .I2 (g9086));
ND2X1 gate18836(.O (g13892), .I1 (g11653), .I2 (g11473));
ND3X1 gate18837(.O (g13476), .I1 (g7503), .I2 (g11336), .I3 (g11869));
ND4X1 gate18838(.O (g21416), .I1 (g17775), .I2 (g14781), .I3 (g17744), .I4 (g14706));
ND2X1 gate18839(.O (I13141), .I1 (g6159), .I2 (I13139));
ND2X1 gate18840(.O (I14249), .I1 (g8091), .I2 (I14247));
ND2X1 gate18841(.O (I17379), .I1 (g13336), .I2 (g1129));
ND2X1 gate18842(.O (I17925), .I1 (g1478), .I2 (I17923));
ND2X1 gate18843(.O (I23949), .I1 (g23162), .I2 (g13603));
ND2X1 gate18844(.O (g14797), .I1 (g12593), .I2 (g12405));
ND3X1 gate18845(.O (g27273), .I1 (g10504), .I2 (g26131), .I3 (g26105));
ND2X1 gate18846(.O (I14482), .I1 (g655), .I2 (I14480));
ND4X1 gate18847(.O (g16687), .I1 (g3255), .I2 (g13700), .I3 (g3325), .I4 (g11519));
ND2X1 gate18848(.O (g13712), .I1 (g8984), .I2 (g11283));
ND4X1 gate18849(.O (g17634), .I1 (g3219), .I2 (g11217), .I3 (g3281), .I4 (g13877));
ND2X1 gate18850(.O (g11914), .I1 (g8187), .I2 (g1648));
ND4X1 gate18851(.O (g17872), .I1 (g6617), .I2 (g14602), .I3 (g6711), .I4 (g12721));
ND2X1 gate18852(.O (g12947), .I1 (g7184), .I2 (g10561));
ND2X1 gate18853(.O (I14248), .I1 (g1322), .I2 (I14247));
ND2X1 gate18854(.O (I22944), .I1 (g9492), .I2 (g19620));
ND4X1 gate18855(.O (g8728), .I1 (g3618), .I2 (g3661), .I3 (g3632), .I4 (g3654));
ND2X1 gate18856(.O (I14204), .I1 (g8508), .I2 (g3821));
ND2X1 gate18857(.O (g25300), .I1 (g22369), .I2 (g12018));
ND3X1 gate18858(.O (g27463), .I1 (g287), .I2 (g26330), .I3 (g23204));
ND4X1 gate18859(.O (g13907), .I1 (g3941), .I2 (g11225), .I3 (g4023), .I4 (g11631));
ND2X1 gate18860(.O (g28381), .I1 (g27074), .I2 (g13621));
ND2X1 gate18861(.O (g29057), .I1 (g27800), .I2 (g9649));
ND2X1 gate18862(.O (g12463), .I1 (g7513), .I2 (g6322));
ND2X1 gate18863(.O (g14136), .I1 (g11571), .I2 (g8906));
ND2X1 gate18864(.O (g14408), .I1 (g6069), .I2 (g11924));
ND2X1 gate18865(.O (g12972), .I1 (g7209), .I2 (g10578));
ND2X1 gate18866(.O (g28174), .I1 (g1270), .I2 (g27059));
ND3X1 gate18867(.O (g28796), .I1 (g27858), .I2 (g7418), .I3 (g7335));
ND2X1 gate18868(.O (g31753), .I1 (I29314), .I2 (I29315));
ND2X1 gate18869(.O (I22793), .I1 (g11956), .I2 (I22792));
ND3X1 gate18870(.O (g16260), .I1 (g4888), .I2 (g13910), .I3 (g12088));
ND2X1 gate18871(.O (g7823), .I1 (I12218), .I2 (I12219));
ND3X1 gate18872(.O (g28840), .I1 (g27858), .I2 (g7380), .I3 (g2287));
ND3X1 gate18873(.O (g11382), .I1 (g8644), .I2 (g6895), .I3 (g8663));
ND2X1 gate18874(.O (I15176), .I1 (g2661), .I2 (I15174));
ND2X1 gate18875(.O (I12203), .I1 (g1094), .I2 (g1135));
ND3X1 gate18876(.O (g19632), .I1 (g1413), .I2 (g1542), .I3 (g16047));
ND2X1 gate18877(.O (I24440), .I1 (g14411), .I2 (I24438));
ND2X1 gate18878(.O (g11675), .I1 (g8984), .I2 (g4912));
ND4X1 gate18879(.O (g13176), .I1 (g10715), .I2 (g7675), .I3 (g1322), .I4 (g1404));
ND2X1 gate18880(.O (g13092), .I1 (g1061), .I2 (g10761));
ND2X1 gate18881(.O (g26269), .I1 (I25243), .I2 (I25244));
ND3X1 gate18882(.O (g34550), .I1 (g626), .I2 (g34359), .I3 (g12323));
ND2X1 gate18883(.O (g11154), .I1 (I14212), .I2 (I14213));
ND2X1 gate18884(.O (g29737), .I1 (g28421), .I2 (g13779));
ND3X1 gate18885(.O (g28522), .I1 (g10857), .I2 (g26131), .I3 (g27142));
ND2X1 gate18886(.O (g8678), .I1 (g376), .I2 (g358));
ND2X1 gate18887(.O (g17592), .I1 (I18530), .I2 (I18531));
ND3X1 gate18888(.O (g16893), .I1 (g10685), .I2 (g13252), .I3 (g703));
ND2X1 gate18889(.O (g10537), .I1 (g7138), .I2 (g5366));
ND2X1 gate18890(.O (I14331), .I1 (g225), .I2 (I14330));
ND2X1 gate18891(.O (g8105), .I1 (g3068), .I2 (g3072));
ND2X1 gate18892(.O (I31984), .I1 (g33653), .I2 (I31983));
ND2X1 gate18893(.O (g16713), .I1 (I17924), .I2 (I17925));
ND2X1 gate18894(.O (I20462), .I1 (g14187), .I2 (I20460));
ND2X1 gate18895(.O (I29255), .I1 (g12017), .I2 (I29253));
ND2X1 gate18896(.O (I24462), .I1 (g23796), .I2 (I24461));
ND4X1 gate18897(.O (g17820), .I1 (g5925), .I2 (g14549), .I3 (g6019), .I4 (g12614));
ND2X1 gate18898(.O (g31709), .I1 (I29285), .I2 (I29286));
ND4X1 gate18899(.O (g15752), .I1 (g5921), .I2 (g12129), .I3 (g5983), .I4 (g14701));
ND2X1 gate18900(.O (I29270), .I1 (g29486), .I2 (I29269));
ND2X1 gate18901(.O (g28949), .I1 (g27903), .I2 (g14643));
ND2X1 gate18902(.O (I13463), .I1 (g2380), .I2 (I13462));
ND2X1 gate18903(.O (g31708), .I1 (I29278), .I2 (I29279));
ND4X1 gate18904(.O (g17846), .I1 (g6271), .I2 (g14575), .I3 (g6365), .I4 (g12672));
ND2X1 gate18905(.O (g17396), .I1 (g7345), .I2 (g14272));
ND4X1 gate18906(.O (g14750), .I1 (g6633), .I2 (g12137), .I3 (g6715), .I4 (g12721));
ND3X1 gate18907(.O (g24584), .I1 (g22852), .I2 (g22836), .I3 (g22715));
ND2X1 gate18908(.O (I14212), .I1 (g9252), .I2 (I14211));
ND2X1 gate18909(.O (g7167), .I1 (g5360), .I2 (g5406));
ND2X1 gate18910(.O (g10796), .I1 (g7537), .I2 (g7523));
ND2X1 gate18911(.O (g20107), .I1 (g11404), .I2 (g17794));
ND2X1 gate18912(.O (g11906), .I1 (I14713), .I2 (I14714));
ND2X1 gate18913(.O (I12403), .I1 (g3813), .I2 (I12401));
ND2X1 gate18914(.O (g16093), .I1 (I17461), .I2 (I17462));
ND3X1 gate18915(.O (g12344), .I1 (g10093), .I2 (g7041), .I3 (g10130));
ND3X1 gate18916(.O (g13083), .I1 (g4392), .I2 (g10590), .I3 (g4434));
ND2X1 gate18917(.O (I32441), .I1 (g34220), .I2 (I32439));
ND2X1 gate18918(.O (g13284), .I1 (g10695), .I2 (g1157));
ND2X1 gate18919(.O (g7549), .I1 (g1018), .I2 (g1030));
ND2X1 gate18920(.O (g25341), .I1 (g22417), .I2 (g12047));
ND2X1 gate18921(.O (g29722), .I1 (g28410), .I2 (g13742));
ND2X1 gate18922(.O (g25268), .I1 (g21124), .I2 (g23692));
ND4X1 gate18923(.O (g16875), .I1 (g3223), .I2 (g13765), .I3 (g3317), .I4 (g11519));
ND2X1 gate18924(.O (g7598), .I1 (I12075), .I2 (I12076));
ND2X1 gate18925(.O (I32758), .I1 (g25779), .I2 (I32756));
ND4X1 gate18926(.O (g14663), .I1 (g5236), .I2 (g12002), .I3 (g5290), .I4 (g12239));
ND2X1 gate18927(.O (g24804), .I1 (g19916), .I2 (g23105));
ND3X1 gate18928(.O (g24652), .I1 (g22712), .I2 (g22940), .I3 (g22757));
ND4X1 gate18929(.O (g13139), .I1 (g6589), .I2 (g12137), .I3 (g6723), .I4 (g10061));
ND4X1 gate18930(.O (g15713), .I1 (g5571), .I2 (g14425), .I3 (g5673), .I4 (g9864));
ND2X1 gate18931(.O (I14369), .I1 (g8481), .I2 (I14368));
ND2X1 gate18932(.O (g34469), .I1 (I32517), .I2 (I32518));
ND2X1 gate18933(.O (I15333), .I1 (g10152), .I2 (g2116));
ND3X1 gate18934(.O (g19546), .I1 (g15969), .I2 (g10841), .I3 (g10884));
ND2X1 gate18935(.O (g8227), .I1 (g3770), .I2 (g3774));
ND2X1 gate18936(.O (I14368), .I1 (g8481), .I2 (g3303));
ND2X1 gate18937(.O (g12028), .I1 (I14884), .I2 (I14885));
ND2X1 gate18938(.O (g15042), .I1 (g12806), .I2 (g10491));
ND2X1 gate18939(.O (g21253), .I1 (g6423), .I2 (g17482));
ND2X1 gate18940(.O (I29277), .I1 (g29488), .I2 (g12081));
ND2X1 gate18941(.O (g23781), .I1 (I22937), .I2 (I22938));
ND2X1 gate18942(.O (g13963), .I1 (g11715), .I2 (g11584));
ND4X1 gate18943(.O (g17640), .I1 (g5264), .I2 (g14399), .I3 (g5335), .I4 (g12497));
ND2X1 gate18944(.O (I14229), .I1 (g979), .I2 (I14228));
ND4X1 gate18945(.O (g21351), .I1 (g15729), .I2 (g13098), .I3 (g15720), .I4 (g13069));
ND2X1 gate18946(.O (g26666), .I1 (g9229), .I2 (g25144));
ND2X1 gate18947(.O (I14228), .I1 (g979), .I2 (g8055));
ND2X1 gate18948(.O (g15030), .I1 (g12716), .I2 (g12680));
ND4X1 gate18949(.O (g27903), .I1 (g21228), .I2 (g25316), .I3 (g26424), .I4 (g26218));
ND3X1 gate18950(.O (g13554), .I1 (g11336), .I2 (g7582), .I3 (g1351));
ND2X1 gate18951(.O (I17924), .I1 (g13378), .I2 (I17923));
ND3X1 gate18952(.O (g12491), .I1 (g7285), .I2 (g4462), .I3 (g6961));
ND3X1 gate18953(.O (g28780), .I1 (g27742), .I2 (g7308), .I3 (g1636));
ND2X1 gate18954(.O (I22753), .I1 (g11937), .I2 (g21434));
ND2X1 gate18955(.O (g11312), .I1 (g8565), .I2 (g3794));
ND2X1 gate18956(.O (g11200), .I1 (g8592), .I2 (g3798));
ND2X1 gate18957(.O (g25038), .I1 (g21331), .I2 (g23363));
ND3X1 gate18958(.O (g13115), .I1 (g1008), .I2 (g11786), .I3 (g11294));
ND2X1 gate18959(.O (I15052), .I1 (g9759), .I2 (I15051));
ND2X1 gate18960(.O (g14933), .I1 (g12700), .I2 (g12571));
ND2X1 gate18961(.O (I14925), .I1 (g5835), .I2 (I14923));
ND2X1 gate18962(.O (g16155), .I1 (I17495), .I2 (I17496));
ND2X1 gate18963(.O (g17662), .I1 (I18634), .I2 (I18635));
ND3X1 gate18964(.O (g28820), .I1 (g27742), .I2 (g1668), .I3 (g1592));
ND2X1 gate18965(.O (I12546), .I1 (g194), .I2 (I12544));
ND2X1 gate18966(.O (I17461), .I1 (g13378), .I2 (I17460));
ND2X1 gate18967(.O (g14851), .I1 (g7738), .I2 (g12505));
ND2X1 gate18968(.O (g27767), .I1 (I26367), .I2 (I26368));
ND2X1 gate18969(.O (g9775), .I1 (g4831), .I2 (g4681));
ND4X1 gate18970(.O (g20371), .I1 (g16956), .I2 (g14088), .I3 (g16694), .I4 (g16660));
ND2X1 gate18971(.O (g24951), .I1 (g199), .I2 (g23088));
ND2X1 gate18972(.O (g24972), .I1 (g19962), .I2 (g23172));
ND2X1 gate18973(.O (g12767), .I1 (g4467), .I2 (g6961));
ND2X1 gate18974(.O (g13798), .I1 (g11280), .I2 (g3423));
ND2X1 gate18975(.O (g11973), .I1 (g8365), .I2 (g2051));
ND2X1 gate18976(.O (g30580), .I1 (g29335), .I2 (g19666));
ND2X1 gate18977(.O (g29657), .I1 (g28363), .I2 (g13634));
ND4X1 gate18978(.O (g17779), .I1 (g6637), .I2 (g14556), .I3 (g6704), .I4 (g12471));
ND2X1 gate18979(.O (g11674), .I1 (g8676), .I2 (g4674));
ND2X1 gate18980(.O (g7879), .I1 (I12262), .I2 (I12263));
ND2X1 gate18981(.O (g23726), .I1 (g9559), .I2 (g21140));
ND2X1 gate18982(.O (I20203), .I1 (g16246), .I2 (g11147));
ND2X1 gate18983(.O (g16524), .I1 (g13822), .I2 (g13798));
ND2X1 gate18984(.O (g26685), .I1 (g9264), .I2 (g25160));
ND2X1 gate18985(.O (I14429), .I1 (g4005), .I2 (I14427));
ND2X1 gate18986(.O (g14574), .I1 (g12256), .I2 (g6120));
ND2X1 gate18987(.O (g12191), .I1 (I15052), .I2 (I15053));
ND4X1 gate18988(.O (g14452), .I1 (g3538), .I2 (g11207), .I3 (g3649), .I4 (g8542));
ND2X1 gate18989(.O (g11934), .I1 (g8139), .I2 (g8187));
ND2X1 gate18990(.O (g16119), .I1 (I17475), .I2 (I17476));
ND2X1 gate18991(.O (I14428), .I1 (g8595), .I2 (I14427));
ND2X1 gate18992(.O (g12521), .I1 (g7471), .I2 (g5969));
ND4X1 gate18993(.O (g17647), .I1 (g5905), .I2 (g14497), .I3 (g5976), .I4 (g12614));
ND2X1 gate18994(.O (I29313), .I1 (g29501), .I2 (g12154));
ND2X1 gate18995(.O (g8609), .I1 (g1171), .I2 (g1157));
ND2X1 gate18996(.O (g19450), .I1 (g11471), .I2 (g17794));
ND2X1 gate18997(.O (I14765), .I1 (g9808), .I2 (I14764));
ND2X1 gate18998(.O (g11761), .I1 (I14610), .I2 (I14611));
ND2X1 gate18999(.O (g22651), .I1 (g20114), .I2 (g2873));
ND2X1 gate19000(.O (I29285), .I1 (g29489), .I2 (I29284));
ND2X1 gate19001(.O (g14051), .I1 (g10323), .I2 (g11527));
ND2X1 gate19002(.O (g14072), .I1 (g11571), .I2 (g11483));
ND4X1 gate19003(.O (g16749), .I1 (g3957), .I2 (g13772), .I3 (g4027), .I4 (g11631));
ND2X1 gate19004(.O (g20163), .I1 (g16663), .I2 (g13938));
ND4X1 gate19005(.O (g15782), .I1 (g6585), .I2 (g14556), .I3 (g6697), .I4 (g10061));
ND2X1 gate19006(.O (I29254), .I1 (g29482), .I2 (I29253));
ND2X1 gate19007(.O (I15214), .I1 (g1714), .I2 (I15212));
ND4X1 gate19008(.O (g14780), .I1 (g6275), .I2 (g12101), .I3 (g6329), .I4 (g12423));
ND2X1 gate19009(.O (g12045), .I1 (g1783), .I2 (g8146));
ND3X1 gate19010(.O (g10820), .I1 (g9985), .I2 (g9920), .I3 (g9843));
ND4X1 gate19011(.O (g14820), .I1 (g6307), .I2 (g12173), .I3 (g6315), .I4 (g12423));
ND4X1 gate19012(.O (g17513), .I1 (g3247), .I2 (g13765), .I3 (g3325), .I4 (g8481));
ND3X1 gate19013(.O (g28827), .I1 (g27837), .I2 (g7362), .I3 (g1862));
ND2X1 gate19014(.O (g25531), .I1 (g22763), .I2 (g2868));
ND3X1 gate19015(.O (g15853), .I1 (g14714), .I2 (g9417), .I3 (g12337));
ND2X1 gate19016(.O (I15241), .I1 (g10003), .I2 (g6351));
ND3X1 gate19017(.O (g12462), .I1 (g7051), .I2 (g7064), .I3 (g10190));
ND2X1 gate19018(.O (g13241), .I1 (g7503), .I2 (g10544));
ND2X1 gate19019(.O (g25186), .I1 (g5396), .I2 (g23602));
ND2X1 gate19020(.O (g14691), .I1 (g12695), .I2 (g12505));
ND3X1 gate19021(.O (g25953), .I1 (g22756), .I2 (g24570), .I3 (g22688));
ND2X1 gate19022(.O (g8803), .I1 (g128), .I2 (g4646));
ND2X1 gate19023(.O (g9954), .I1 (g6128), .I2 (g6120));
ND2X1 gate19024(.O (I22792), .I1 (g11956), .I2 (g21434));
ND2X1 gate19025(.O (I22967), .I1 (g21228), .I2 (I22965));
ND4X1 gate19026(.O (g13100), .I1 (g6581), .I2 (g12137), .I3 (g6692), .I4 (g10061));
ND2X1 gate19027(.O (g23575), .I1 (I22711), .I2 (I22712));
ND2X1 gate19028(.O (g20173), .I1 (g16696), .I2 (g13972));
ND2X1 gate19029(.O (g10929), .I1 (g1099), .I2 (g7854));
ND2X1 gate19030(.O (g31669), .I1 (I29254), .I2 (I29255));
ND3X1 gate19031(.O (g15864), .I1 (g14833), .I2 (g12543), .I3 (g12487));
ND2X1 gate19032(.O (g33669), .I1 (g33378), .I2 (g862));
ND2X1 gate19033(.O (g25334), .I1 (g21253), .I2 (g23756));
ND4X1 gate19034(.O (g17723), .I1 (g6597), .I2 (g14556), .I3 (g6668), .I4 (g12721));
ND2X1 gate19035(.O (g10583), .I1 (g7475), .I2 (g862));
ND3X1 gate19036(.O (g10928), .I1 (g8181), .I2 (g8137), .I3 (g417));
ND4X1 gate19037(.O (g15748), .I1 (g13257), .I2 (g13130), .I3 (g7922), .I4 (g13241));
ND2X1 gate19038(.O (g21283), .I1 (g11291), .I2 (g17157));
ND2X1 gate19039(.O (g9912), .I1 (I13463), .I2 (I13464));
ND2X1 gate19040(.O (I13045), .I1 (g5120), .I2 (I13043));
ND4X1 gate19041(.O (g20134), .I1 (g17572), .I2 (g14542), .I3 (g17495), .I4 (g14452));
ND4X1 gate19042(.O (g13515), .I1 (g12628), .I2 (g12588), .I3 (g12524), .I4 (g12464));
ND4X1 gate19043(.O (g13882), .I1 (g3590), .I2 (g11207), .I3 (g3672), .I4 (g11576));
ND2X1 gate19044(.O (g24760), .I1 (I23918), .I2 (I23919));
ND2X1 gate19045(.O (I23961), .I1 (g23184), .I2 (g13631));
ND2X1 gate19046(.O (g25216), .I1 (g6088), .I2 (g23678));
ND2X1 gate19047(.O (g14113), .I1 (g11626), .I2 (g11537));
ND2X1 gate19048(.O (I24385), .I1 (g14347), .I2 (I24383));
ND2X1 gate19049(.O (g15036), .I1 (g12780), .I2 (g12581));
ND2X1 gate19050(.O (g19597), .I1 (g1199), .I2 (g15995));
ND2X1 gate19051(.O (g12629), .I1 (g7812), .I2 (g7142));
ND2X1 gate19052(.O (I12877), .I1 (g4200), .I2 (I12876));
ND2X1 gate19053(.O (I13462), .I1 (g2380), .I2 (g2384));
ND2X1 gate19054(.O (g8847), .I1 (g4831), .I2 (g4681));
ND3X1 gate19055(.O (g12628), .I1 (g7074), .I2 (g6336), .I3 (g6390));
ND3X1 gate19056(.O (g22850), .I1 (g1536), .I2 (g19581), .I3 (g10699));
ND2X1 gate19057(.O (g11441), .I1 (g9599), .I2 (g3267));
ND2X1 gate19058(.O (I13140), .I1 (g6154), .I2 (I13139));
ND2X1 gate19059(.O (I22901), .I1 (g21228), .I2 (I22899));
ND3X1 gate19060(.O (g28786), .I1 (g27837), .I2 (g7405), .I3 (g7322));
ND2X1 gate19061(.O (g11206), .I1 (I14276), .I2 (I14277));
ND3X1 gate19062(.O (g16238), .I1 (g4698), .I2 (g13883), .I3 (g12054));
ND2X1 gate19063(.O (I14499), .I1 (g8737), .I2 (I14497));
ND2X1 gate19064(.O (g17412), .I1 (g14520), .I2 (g14489));
ND2X1 gate19065(.O (I18625), .I1 (g2079), .I2 (g14712));
ND2X1 gate19066(.O (g14768), .I1 (g12662), .I2 (g12571));
ND2X1 gate19067(.O (g28945), .I1 (g27854), .I2 (g8211));
ND4X1 gate19068(.O (g14803), .I1 (g5208), .I2 (g12059), .I3 (g5308), .I4 (g12497));
ND2X1 gate19069(.O (I14498), .I1 (g9020), .I2 (I14497));
ND3X1 gate19070(.O (g33679), .I1 (g33394), .I2 (g10737), .I3 (g10308));
ND2X1 gate19071(.O (g12147), .I1 (g8302), .I2 (g8201));
ND2X1 gate19072(.O (I12402), .I1 (g3808), .I2 (I12401));
ND2X1 gate19073(.O (I15107), .I1 (g5313), .I2 (I15105));
ND2X1 gate19074(.O (I22823), .I1 (g11978), .I2 (I22822));
ND2X1 gate19075(.O (I14611), .I1 (g8678), .I2 (I14609));
ND2X1 gate19076(.O (I14924), .I1 (g9558), .I2 (I14923));
ND2X1 gate19077(.O (g12370), .I1 (I15213), .I2 (I15214));
ND2X1 gate19078(.O (g25974), .I1 (g24576), .I2 (g22837));
ND4X1 gate19079(.O (g17716), .I1 (g5957), .I2 (g14497), .I3 (g6027), .I4 (g12614));
ND2X1 gate19080(.O (g15008), .I1 (g12780), .I2 (g10341));
ND2X1 gate19081(.O (I23971), .I1 (g490), .I2 (I23969));
ND2X1 gate19082(.O (g25293), .I1 (g21190), .I2 (g23726));
ND2X1 gate19083(.O (g12151), .I1 (g8316), .I2 (g8211));
ND2X1 gate19084(.O (g19854), .I1 (I20222), .I2 (I20223));
ND4X1 gate19085(.O (g13940), .I1 (g11426), .I2 (g8889), .I3 (g11707), .I4 (g8829));
ND2X1 gate19086(.O (I22966), .I1 (g12288), .I2 (I22965));
ND2X1 gate19087(.O (g23949), .I1 (g7074), .I2 (g21012));
ND2X1 gate19088(.O (g28448), .I1 (g23975), .I2 (g27377));
ND2X1 gate19089(.O (I15263), .I1 (g10081), .I2 (I15262));
ND2X1 gate19090(.O (g10552), .I1 (g2153), .I2 (g7374));
ND4X1 gate19091(.O (g8751), .I1 (g3969), .I2 (g4012), .I3 (g3983), .I4 (g4005));
ND3X1 gate19092(.O (g15907), .I1 (g14833), .I2 (g9417), .I3 (g12487));
ND2X1 gate19093(.O (g22681), .I1 (I21993), .I2 (I21994));
ND2X1 gate19094(.O (g11135), .I1 (I14186), .I2 (I14187));
ND2X1 gate19095(.O (I14330), .I1 (g225), .I2 (g9966));
ND2X1 gate19096(.O (g19916), .I1 (g3029), .I2 (g16313));
ND4X1 gate19097(.O (g16728), .I1 (g13884), .I2 (g13870), .I3 (g14089), .I4 (g11639));
ND2X1 gate19098(.O (g12227), .I1 (g8418), .I2 (g8330));
ND2X1 gate19099(.O (I14764), .I1 (g9808), .I2 (g5821));
ND2X1 gate19100(.O (g11962), .I1 (I14789), .I2 (I14790));
ND2X1 gate19101(.O (I29284), .I1 (g29489), .I2 (g12085));
ND2X1 gate19102(.O (I31973), .I1 (g33641), .I2 (I31972));
ND2X1 gate19103(.O (I29304), .I1 (g12121), .I2 (I29302));
ND2X1 gate19104(.O (I18581), .I1 (g14678), .I2 (I18579));
ND2X1 gate19105(.O (I26051), .I1 (g13500), .I2 (I26049));
ND2X1 gate19106(.O (I25847), .I1 (g24799), .I2 (I25845));
ND2X1 gate19107(.O (I26072), .I1 (g13517), .I2 (I26070));
ND2X1 gate19108(.O (I11825), .I1 (g4593), .I2 (I11824));
ND2X1 gate19109(.O (I12876), .I1 (g4200), .I2 (g4180));
ND2X1 gate19110(.O (g14999), .I1 (g12739), .I2 (g12824));
ND3X1 gate19111(.O (g16304), .I1 (g4765), .I2 (g13970), .I3 (g12054));
ND2X1 gate19112(.O (g12044), .I1 (g1657), .I2 (g8139));
ND2X1 gate19113(.O (I15004), .I1 (g1700), .I2 (I15002));
ND4X1 gate19114(.O (g21509), .I1 (g17820), .I2 (g14898), .I3 (g17647), .I4 (g17608));
ND4X1 gate19115(.O (g17765), .I1 (g6649), .I2 (g14556), .I3 (g6719), .I4 (g12721));
ND2X1 gate19116(.O (I14259), .I1 (g3133), .I2 (I14257));
ND2X1 gate19117(.O (I17495), .I1 (g13378), .I2 (I17494));
ND2X1 gate19118(.O (g27377), .I1 (g10685), .I2 (g25930));
ND4X1 gate19119(.O (g24926), .I1 (g20172), .I2 (g20163), .I3 (g23357), .I4 (g13995));
ND2X1 gate19120(.O (g25275), .I1 (g22342), .I2 (g11991));
ND2X1 gate19121(.O (g12301), .I1 (I15148), .I2 (I15149));
ND2X1 gate19122(.O (I14258), .I1 (g8154), .I2 (I14257));
ND2X1 gate19123(.O (g12120), .I1 (g2476), .I2 (g8273));
ND4X1 gate19124(.O (g27738), .I1 (g21228), .I2 (g25243), .I3 (g26424), .I4 (g26148));
ND2X1 gate19125(.O (I32440), .I1 (g34227), .I2 (I32439));
ND2X1 gate19126(.O (g25237), .I1 (g6434), .I2 (g23711));
ND2X1 gate19127(.O (I15106), .I1 (g9780), .I2 (I15105));
ND2X1 gate19128(.O (g13273), .I1 (g1459), .I2 (g10699));
ND2X1 gate19129(.O (g19335), .I1 (g15717), .I2 (g1056));
ND2X1 gate19130(.O (g10961), .I1 (g1442), .I2 (g7876));
ND3X1 gate19131(.O (g29679), .I1 (g153), .I2 (g28353), .I3 (g23042));
ND4X1 gate19132(.O (g15729), .I1 (g5949), .I2 (g14549), .I3 (g6027), .I4 (g9935));
ND2X1 gate19133(.O (g14505), .I1 (g12073), .I2 (g9961));
ND2X1 gate19134(.O (I12287), .I1 (g1484), .I2 (g1300));
ND2X1 gate19135(.O (I14955), .I1 (g9620), .I2 (g6181));
ND2X1 gate19136(.O (g19965), .I1 (g3380), .I2 (g16424));
ND3X1 gate19137(.O (g11951), .I1 (g9166), .I2 (g847), .I3 (g703));
ND4X1 gate19138(.O (g15728), .I1 (g5200), .I2 (g14399), .I3 (g5313), .I4 (g9780));
ND2X1 gate19139(.O (g13951), .I1 (g10295), .I2 (g11729));
ND2X1 gate19140(.O (I12076), .I1 (g979), .I2 (I12074));
ND2X1 gate19141(.O (g23047), .I1 (g482), .I2 (g20000));
ND2X1 gate19142(.O (g13795), .I1 (g11216), .I2 (g401));
ND3X1 gate19143(.O (g28896), .I1 (g27837), .I2 (g1936), .I3 (g1862));
ND2X1 gate19144(.O (I14171), .I1 (g3119), .I2 (I14169));
ND2X1 gate19145(.O (g20871), .I1 (g14434), .I2 (g17396));
ND2X1 gate19146(.O (I22893), .I1 (g12189), .I2 (I22892));
ND2X1 gate19147(.O (I12269), .I1 (g1141), .I2 (g956));
ND2X1 gate19148(.O (I13044), .I1 (g5115), .I2 (I13043));
ND4X1 gate19149(.O (g17775), .I1 (g6255), .I2 (g14575), .I3 (g6351), .I4 (g12672));
ND2X1 gate19150(.O (I22865), .I1 (g12146), .I2 (I22864));
ND2X1 gate19151(.O (g23756), .I1 (g9621), .I2 (g21206));
ND2X1 gate19152(.O (g14723), .I1 (g7704), .I2 (g12772));
ND2X1 gate19153(.O (g23780), .I1 (I22930), .I2 (I22931));
ND2X1 gate19154(.O (g14433), .I1 (g12035), .I2 (g9890));
ND2X1 gate19155(.O (I24384), .I1 (g23721), .I2 (I24383));
ND4X1 gate19156(.O (g21350), .I1 (g15751), .I2 (g15742), .I3 (g15735), .I4 (g13108));
ND2X1 gate19157(.O (g16312), .I1 (g13580), .I2 (g13574));
ND2X1 gate19158(.O (g14104), .I1 (g11514), .I2 (g8864));
ND2X1 gate19159(.O (I25846), .I1 (g26212), .I2 (I25845));
ND2X1 gate19160(.O (g14343), .I1 (g11961), .I2 (g9670));
ND2X1 gate19161(.O (g10971), .I1 (g7867), .I2 (g7886));
ND2X1 gate19162(.O (g28958), .I1 (g27833), .I2 (g8249));
ND2X1 gate19163(.O (g14971), .I1 (g12667), .I2 (g12581));
ND4X1 gate19164(.O (g16745), .I1 (g3594), .I2 (g13730), .I3 (g3661), .I4 (g11389));
ND2X1 gate19165(.O (g31748), .I1 (I29303), .I2 (I29304));
ND2X1 gate19166(.O (g26208), .I1 (g7975), .I2 (g24751));
ND4X1 gate19167(.O (g16813), .I1 (g3614), .I2 (g13799), .I3 (g3625), .I4 (g8542));
ND2X1 gate19168(.O (I22938), .I1 (g21228), .I2 (I22936));
ND2X1 gate19169(.O (g27824), .I1 (I26394), .I2 (I26395));
ND2X1 gate19170(.O (g13920), .I1 (g11621), .I2 (g11483));
ND2X1 gate19171(.O (I17460), .I1 (g13378), .I2 (g1300));
ND2X1 gate19172(.O (g24591), .I1 (g22833), .I2 (g22642));
ND2X1 gate19173(.O (g24776), .I1 (g3040), .I2 (g23052));
ND2X1 gate19174(.O (I14817), .I1 (g9962), .I2 (I14816));
ND2X1 gate19175(.O (g25236), .I1 (I24415), .I2 (I24416));
ND2X1 gate19176(.O (I15121), .I1 (g9910), .I2 (g2102));
ND2X1 gate19177(.O (g34422), .I1 (I32432), .I2 (I32433));
ND3X1 gate19178(.O (g28857), .I1 (g27779), .I2 (g1802), .I3 (g1728));
ND2X1 gate19179(.O (g14133), .I1 (g11692), .I2 (g11747));
ND2X1 gate19180(.O (I12279), .I1 (g1472), .I2 (I12277));
ND2X1 gate19181(.O (I14532), .I1 (g8873), .I2 (I14530));
ND2X1 gate19182(.O (g13121), .I1 (g11117), .I2 (g8411));
ND3X1 gate19183(.O (g28793), .I1 (g27800), .I2 (g7328), .I3 (g2153));
ND2X1 gate19184(.O (I13403), .I1 (g2250), .I2 (I13401));
ND2X1 gate19185(.O (I12278), .I1 (g1467), .I2 (I12277));
ND2X1 gate19186(.O (g24950), .I1 (g19442), .I2 (g23154));
ND2X1 gate19187(.O (I12469), .I1 (g405), .I2 (I12468));
ND3X1 gate19188(.O (g27931), .I1 (g25425), .I2 (g25381), .I3 (g25780));
ND3X1 gate19189(.O (g28765), .I1 (g27800), .I2 (g7374), .I3 (g7280));
ND2X1 gate19190(.O (g7611), .I1 (g4057), .I2 (g4064));
ND2X1 gate19191(.O (g14011), .I1 (g10295), .I2 (g11473));
ND4X1 gate19192(.O (g20151), .I1 (g17598), .I2 (g14570), .I3 (g17514), .I4 (g14519));
ND2X1 gate19193(.O (g20172), .I1 (g16876), .I2 (g8131));
ND2X1 gate19194(.O (I12468), .I1 (g405), .I2 (g392));
ND2X1 gate19195(.O (g13291), .I1 (g10715), .I2 (g1500));
ND3X1 gate19196(.O (g11173), .I1 (g4966), .I2 (g7898), .I3 (g9064));
ND2X1 gate19197(.O (g12190), .I1 (g8365), .I2 (g8255));
ND2X1 gate19198(.O (g22753), .I1 (g1536), .I2 (g19632));
ND3X1 gate19199(.O (g28504), .I1 (g758), .I2 (g27528), .I3 (g11679));
ND4X1 gate19200(.O (g21357), .I1 (g15736), .I2 (g13109), .I3 (g15726), .I4 (g13086));
ND3X1 gate19201(.O (g31009), .I1 (g27187), .I2 (g29503), .I3 (g19644));
ND2X1 gate19202(.O (g14627), .I1 (g12553), .I2 (g12772));
ND2X1 gate19203(.O (g23357), .I1 (g20201), .I2 (g11231));
ND2X1 gate19204(.O (g14959), .I1 (g12695), .I2 (g12798));
ND2X1 gate19205(.O (g14379), .I1 (g5723), .I2 (g11907));
ND2X1 gate19206(.O (g22650), .I1 (g7888), .I2 (g19581));
ND3X1 gate19207(.O (g11134), .I1 (g8138), .I2 (g8240), .I3 (g8301));
ND2X1 gate19208(.O (g23105), .I1 (g8097), .I2 (g19887));
ND2X1 gate19209(.O (g13134), .I1 (g11134), .I2 (g8470));
ND2X1 gate19210(.O (g14378), .I1 (g11979), .I2 (g9731));
ND2X1 gate19211(.O (g7209), .I1 (g6052), .I2 (g6098));
ND2X1 gate19212(.O (g12024), .I1 (g8381), .I2 (g8418));
ND4X1 gate19213(.O (g17650), .I1 (g6299), .I2 (g12101), .I3 (g6315), .I4 (g14745));
ND2X1 gate19214(.O (g10603), .I1 (g10077), .I2 (g9751));
ND4X1 gate19215(.O (g17736), .I1 (g5563), .I2 (g14522), .I3 (g5659), .I4 (g12563));
ND4X1 gate19216(.O (g15798), .I1 (g6629), .I2 (g14602), .I3 (g6704), .I4 (g14786));
ND2X1 gate19217(.O (g25021), .I1 (g21417), .I2 (g23363));
ND2X1 gate19218(.O (I11824), .I1 (g4593), .I2 (g4601));
ND2X1 gate19219(.O (g15674), .I1 (g921), .I2 (g13110));
ND2X1 gate19220(.O (g9310), .I1 (I13078), .I2 (I13079));
ND2X1 gate19221(.O (I14289), .I1 (g8282), .I2 (g3835));
ND3X1 gate19222(.O (g28298), .I1 (g10533), .I2 (g26131), .I3 (g26990));
ND2X1 gate19223(.O (g9663), .I1 (g128), .I2 (g4646));
ND4X1 gate19224(.O (g13927), .I1 (g3578), .I2 (g11207), .I3 (g3632), .I4 (g11389));
ND2X1 gate19225(.O (I17494), .I1 (g13378), .I2 (g1448));
ND2X1 gate19226(.O (g29118), .I1 (g27886), .I2 (g9755));
ND2X1 gate19227(.O (I12217), .I1 (g1437), .I2 (g1478));
ND4X1 gate19228(.O (g14730), .I1 (g5615), .I2 (g12093), .I3 (g5623), .I4 (g12301));
ND2X1 gate19229(.O (g22709), .I1 (g1193), .I2 (g19611));
ND2X1 gate19230(.O (I22822), .I1 (g11978), .I2 (g21434));
ND2X1 gate19231(.O (g13240), .I1 (g1046), .I2 (g10521));
ND2X1 gate19232(.O (g24957), .I1 (g21359), .I2 (g23462));
ND2X1 gate19233(.O (g11491), .I1 (g9982), .I2 (g4000));
ND2X1 gate19234(.O (g12644), .I1 (g10233), .I2 (g4531));
ND2X1 gate19235(.O (g11903), .I1 (g9099), .I2 (g3712));
ND2X1 gate19236(.O (I14816), .I1 (g9962), .I2 (g6513));
ND2X1 gate19237(.O (I32203), .I1 (g33937), .I2 (I32202));
ND2X1 gate19238(.O (g23890), .I1 (g7004), .I2 (g20682));
ND3X1 gate19239(.O (g12969), .I1 (g4388), .I2 (g7178), .I3 (g10476));
ND2X1 gate19240(.O (I13520), .I1 (g2518), .I2 (I13518));
ND2X1 gate19241(.O (g20645), .I1 (g14344), .I2 (g17243));
ND2X1 gate19242(.O (g28856), .I1 (g27738), .I2 (g8093));
ND2X1 gate19243(.O (g14548), .I1 (g12208), .I2 (g5774));
ND2X1 gate19244(.O (g17225), .I1 (g8612), .I2 (g14367));
ND4X1 gate19245(.O (g17708), .I1 (g5216), .I2 (g14490), .I3 (g5313), .I4 (g12497));
ND2X1 gate19246(.O (g12197), .I1 (g7296), .I2 (g5290));
ND2X1 gate19247(.O (g8434), .I1 (g3080), .I2 (g3072));
ND3X1 gate19248(.O (g28512), .I1 (g10857), .I2 (g27155), .I3 (g27142));
ND2X1 gate19249(.O (g23552), .I1 (I22684), .I2 (I22685));
ND2X1 gate19250(.O (g15005), .I1 (g12667), .I2 (g12622));
ND2X1 gate19251(.O (g14317), .I1 (g5033), .I2 (g11862));
ND2X1 gate19252(.O (g12411), .I1 (g7393), .I2 (g5276));
ND3X1 gate19253(.O (g8347), .I1 (g4358), .I2 (g4349), .I3 (g4340));
ND2X1 gate19254(.O (I15262), .I1 (g10081), .I2 (g2273));
ND2X1 gate19255(.O (g23778), .I1 (I22922), .I2 (I22923));
ND2X1 gate19256(.O (g11395), .I1 (g9601), .I2 (g3983));
ND2X1 gate19257(.O (I13497), .I1 (g255), .I2 (g232));
ND2X1 gate19258(.O (g11990), .I1 (g9166), .I2 (g703));
ND2X1 gate19259(.O (g13990), .I1 (g11669), .I2 (g11584));
ND2X1 gate19260(.O (g23786), .I1 (I22945), .I2 (I22946));
ND2X1 gate19261(.O (I18487), .I1 (g14611), .I2 (I18485));
ND2X1 gate19262(.O (g13898), .I1 (g11621), .I2 (g11747));
ND2X1 gate19263(.O (I22864), .I1 (g12146), .I2 (g21228));
ND4X1 gate19264(.O (g21356), .I1 (g15780), .I2 (g15752), .I3 (g15743), .I4 (g13118));
ND2X1 gate19265(.O (I12373), .I1 (g3457), .I2 (I12372));
ND4X1 gate19266(.O (g14626), .I1 (g12232), .I2 (g9852), .I3 (g12159), .I4 (g9715));
ND3X1 gate19267(.O (g24661), .I1 (g23210), .I2 (g23195), .I3 (g22984));
ND3X1 gate19268(.O (g24547), .I1 (g22638), .I2 (g22643), .I3 (g22754));
ND2X1 gate19269(.O (I31972), .I1 (g33641), .I2 (g33631));
ND2X1 gate19270(.O (g12450), .I1 (g7738), .I2 (g10281));
ND3X1 gate19271(.O (g10775), .I1 (g7960), .I2 (g7943), .I3 (g8470));
ND2X1 gate19272(.O (g9295), .I1 (I13066), .I2 (I13067));
ND2X1 gate19273(.O (g12819), .I1 (g9848), .I2 (g6961));
ND2X1 gate19274(.O (g12910), .I1 (g11002), .I2 (g10601));
ND3X1 gate19275(.O (g34174), .I1 (g617), .I2 (g33851), .I3 (g12323));
ND4X1 gate19276(.O (g17792), .I1 (g6601), .I2 (g14602), .I3 (g6697), .I4 (g12721));
ND2X1 gate19277(.O (I22900), .I1 (g12193), .I2 (I22899));
ND2X1 gate19278(.O (g10737), .I1 (g6961), .I2 (g9848));
ND2X1 gate19279(.O (g25537), .I1 (g22763), .I2 (g2873));
ND2X1 gate19280(.O (g12111), .I1 (g847), .I2 (g9166));
ND3X1 gate19281(.O (g28271), .I1 (g10533), .I2 (g27004), .I3 (g26990));
ND2X1 gate19282(.O (g13861), .I1 (g1459), .I2 (g10671));
ND2X1 gate19283(.O (g21331), .I1 (g11402), .I2 (g17157));
ND4X1 gate19284(.O (g13573), .I1 (g8002), .I2 (g10544), .I3 (g7582), .I4 (g1351));
ND2X1 gate19285(.O (g23932), .I1 (g7051), .I2 (g20875));
ND2X1 gate19286(.O (I14713), .I1 (g9671), .I2 (I14712));
ND3X1 gate19287(.O (g12590), .I1 (g7097), .I2 (g7110), .I3 (g10229));
ND2X1 gate19288(.O (g33083), .I1 (g7805), .I2 (g32118));
ND2X1 gate19289(.O (g11389), .I1 (I14399), .I2 (I14400));
ND2X1 gate19290(.O (g25492), .I1 (g12479), .I2 (g22457));
ND2X1 gate19291(.O (g14697), .I1 (g12662), .I2 (g12824));
ND2X1 gate19292(.O (g9966), .I1 (I13498), .I2 (I13499));
ND2X1 gate19293(.O (g7184), .I1 (g5706), .I2 (g5752));
ND2X1 gate19294(.O (g9705), .I1 (g2619), .I2 (g2587));
ND2X1 gate19295(.O (I14610), .I1 (g8993), .I2 (I14609));
ND2X1 gate19296(.O (I26368), .I1 (g14211), .I2 (I26366));
ND2X1 gate19297(.O (I29263), .I1 (g12046), .I2 (I29261));
ND2X1 gate19298(.O (g11534), .I1 (g7121), .I2 (g8958));
ND2X1 gate19299(.O (I23602), .I1 (g4322), .I2 (I23600));
ND2X1 gate19300(.O (g20784), .I1 (g14616), .I2 (g17595));
ND3X1 gate19301(.O (g28736), .I1 (g27742), .I2 (g7308), .I3 (g7252));
ND4X1 gate19302(.O (g19265), .I1 (g15721), .I2 (g15715), .I3 (g13091), .I4 (g15710));
ND4X1 gate19303(.O (g13098), .I1 (g5933), .I2 (g12129), .I3 (g6023), .I4 (g9935));
ND2X1 gate19304(.O (I20487), .I1 (g16696), .I2 (I20486));
ND2X1 gate19305(.O (g11251), .I1 (g8438), .I2 (g3092));
ND2X1 gate19306(.O (g25381), .I1 (g538), .I2 (g23088));
ND2X1 gate19307(.O (I23970), .I1 (g22202), .I2 (I23969));
ND4X1 gate19308(.O (g13462), .I1 (g12449), .I2 (g12412), .I3 (g12342), .I4 (g12294));
ND3X1 gate19309(.O (g28843), .I1 (g27907), .I2 (g7456), .I3 (g7387));
ND3X1 gate19310(.O (g19510), .I1 (g15969), .I2 (g10841), .I3 (g10899));
ND2X1 gate19311(.O (g20181), .I1 (g13252), .I2 (g16846));
ND2X1 gate19312(.O (g12019), .I1 (g7322), .I2 (g1906));
ND4X1 gate19313(.O (g17598), .I1 (g3949), .I2 (g13824), .I3 (g4027), .I4 (g8595));
ND2X1 gate19314(.O (g12196), .I1 (g8764), .I2 (g4688));
ND2X1 gate19315(.O (g11997), .I1 (g2319), .I2 (g8316));
ND2X1 gate19316(.O (I20469), .I1 (g16728), .I2 (I20467));
ND2X1 gate19317(.O (I21994), .I1 (g19638), .I2 (I21992));
ND2X1 gate19318(.O (I12242), .I1 (g1105), .I2 (I12240));
ND3X1 gate19319(.O (g12526), .I1 (g10194), .I2 (g7110), .I3 (g10213));
ND4X1 gate19320(.O (g15725), .I1 (g5603), .I2 (g14522), .I3 (g5681), .I4 (g9864));
ND2X1 gate19321(.O (I20468), .I1 (g16663), .I2 (I20467));
ND2X1 gate19322(.O (g29154), .I1 (g27937), .I2 (g9835));
ND4X1 gate19323(.O (g21433), .I1 (g17792), .I2 (g14830), .I3 (g17765), .I4 (g14750));
ND2X1 gate19324(.O (I22892), .I1 (g12189), .I2 (g21228));
ND2X1 gate19325(.O (g19442), .I1 (g11431), .I2 (g17794));
ND2X1 gate19326(.O (g12402), .I1 (g7704), .I2 (g10266));
ND2X1 gate19327(.O (g10611), .I1 (g10115), .I2 (g9831));
ND2X1 gate19328(.O (I13111), .I1 (g5813), .I2 (I13109));
ND2X1 gate19329(.O (g13871), .I1 (g4955), .I2 (g11834));
ND2X1 gate19330(.O (I23919), .I1 (g9333), .I2 (I23917));
ND2X1 gate19331(.O (I18486), .I1 (g1677), .I2 (I18485));
ND3X1 gate19332(.O (g28259), .I1 (g10504), .I2 (g26987), .I3 (g26973));
ND2X1 gate19333(.O (g14924), .I1 (g12558), .I2 (g12505));
ND2X1 gate19334(.O (I22712), .I1 (g21434), .I2 (I22710));
ND2X1 gate19335(.O (g17656), .I1 (I18626), .I2 (I18627));
ND2X1 gate19336(.O (I20187), .I1 (g16272), .I2 (g1333));
ND4X1 gate19337(.O (g15744), .I1 (g6641), .I2 (g14602), .I3 (g6719), .I4 (g10061));
ND2X1 gate19338(.O (I17476), .I1 (g1105), .I2 (I17474));
ND2X1 gate19339(.O (I23918), .I1 (g23975), .I2 (I23917));
ND2X1 gate19340(.O (I18580), .I1 (g1945), .I2 (I18579));
ND2X1 gate19341(.O (I26050), .I1 (g25997), .I2 (I26049));
ND2X1 gate19342(.O (I13384), .I1 (g246), .I2 (I13382));
ND2X1 gate19343(.O (g12001), .I1 (I14854), .I2 (I14855));
ND2X1 gate19344(.O (I13067), .I1 (g4304), .I2 (I13065));
ND2X1 gate19345(.O (I12841), .I1 (g4222), .I2 (I12840));
ND2X1 gate19346(.O (I11877), .I1 (g4388), .I2 (g4430));
ND2X1 gate19347(.O (g10529), .I1 (g1592), .I2 (g7308));
ND2X1 gate19348(.O (g13628), .I1 (g3372), .I2 (g11107));
ND2X1 gate19349(.O (g23850), .I1 (g12185), .I2 (g19462));
ND2X1 gate19350(.O (g13911), .I1 (g11834), .I2 (g4917));
ND2X1 gate19351(.O (I18531), .I1 (g14640), .I2 (I18529));
ND2X1 gate19352(.O (g17364), .I1 (g8639), .I2 (g14367));
ND3X1 gate19353(.O (g28955), .I1 (g27837), .I2 (g1936), .I3 (g7362));
ND2X1 gate19354(.O (I14277), .I1 (g3484), .I2 (I14275));
ND2X1 gate19355(.O (I21977), .I1 (g7680), .I2 (I21976));
ND4X1 gate19356(.O (g14696), .I1 (g5567), .I2 (g12093), .I3 (g5685), .I4 (g12563));
ND2X1 gate19357(.O (I24363), .I1 (g23687), .I2 (g14320));
ND2X1 gate19358(.O (g8163), .I1 (g3419), .I2 (g3423));
ND3X1 gate19359(.O (g15962), .I1 (g14833), .I2 (g9417), .I3 (g9340));
ND2X1 gate19360(.O (g14764), .I1 (g7738), .I2 (g12798));
ND2X1 gate19361(.O (g11591), .I1 (I14531), .I2 (I14532));
ND3X1 gate19362(.O (g21011), .I1 (g14504), .I2 (g17399), .I3 (g9629));
ND2X1 gate19363(.O (I15147), .I1 (g9864), .I2 (g5659));
ND2X1 gate19364(.O (g12066), .I1 (I14924), .I2 (I14925));
ND2X1 gate19365(.O (I20486), .I1 (g16696), .I2 (g16757));
ND2X1 gate19366(.O (g24943), .I1 (g20068), .I2 (g23172));
ND3X1 gate19367(.O (g20644), .I1 (g14342), .I2 (g17220), .I3 (g9372));
ND2X1 gate19368(.O (g27876), .I1 (I26418), .I2 (I26419));
ND3X1 gate19369(.O (g15833), .I1 (g14714), .I2 (g12378), .I3 (g12337));
ND2X1 gate19370(.O (I13402), .I1 (g2246), .I2 (I13401));
ND2X1 gate19371(.O (g11355), .I1 (g9551), .I2 (g3310));
ND3X1 gate19372(.O (g28994), .I1 (g27907), .I2 (g2495), .I3 (g7424));
ND2X1 gate19373(.O (g14868), .I1 (g12755), .I2 (g12680));
ND2X1 gate19374(.O (g17571), .I1 (g8579), .I2 (g14367));
ND2X1 gate19375(.O (I11866), .I1 (g4401), .I2 (I11864));
ND4X1 gate19376(.O (g27854), .I1 (g21228), .I2 (g25283), .I3 (g26424), .I4 (g26195));
ND2X1 gate19377(.O (g25062), .I1 (g21403), .I2 (g23363));
ND2X1 gate19378(.O (I20223), .I1 (g11170), .I2 (I20221));
ND2X1 gate19379(.O (g16507), .I1 (g13797), .I2 (g13764));
ND2X1 gate19380(.O (g11858), .I1 (g9014), .I2 (g3010));
ND2X1 gate19381(.O (I14352), .I1 (g8848), .I2 (I14350));
ND2X1 gate19382(.O (I17883), .I1 (g13336), .I2 (g1135));
ND2X1 gate19383(.O (g11172), .I1 (g8478), .I2 (g3096));
ND3X1 gate19384(.O (g12511), .I1 (g7028), .I2 (g5644), .I3 (g5698));
ND2X1 gate19385(.O (g22687), .I1 (g19560), .I2 (g7870));
ND2X1 gate19386(.O (g7885), .I1 (I12270), .I2 (I12271));
ND2X1 gate19387(.O (g11996), .I1 (g7280), .I2 (g2197));
ND4X1 gate19388(.O (g17495), .I1 (g3566), .I2 (g13730), .I3 (g3668), .I4 (g8542));
ND2X1 gate19389(.O (g23379), .I1 (g20216), .I2 (g11248));
ND2X1 gate19390(.O (I14170), .I1 (g8389), .I2 (I14169));
ND2X1 gate19391(.O (I13077), .I1 (g5462), .I2 (g5467));
ND2X1 gate19392(.O (g23112), .I1 (g21024), .I2 (g10733));
ND3X1 gate19393(.O (g20870), .I1 (g14432), .I2 (g17315), .I3 (g9567));
ND4X1 gate19394(.O (g17816), .I1 (g6657), .I2 (g14602), .I3 (g6668), .I4 (g10061));
ND2X1 gate19395(.O (g14258), .I1 (g9203), .I2 (g11903));
ND2X1 gate19396(.O (g11394), .I1 (g9600), .I2 (g3661));
ND2X1 gate19397(.O (g22643), .I1 (g20136), .I2 (g18954));
ND2X1 gate19398(.O (g34051), .I1 (I31973), .I2 (I31974));
ND4X1 gate19399(.O (g21386), .I1 (g15798), .I2 (g15788), .I3 (g15782), .I4 (g13139));
ND2X1 gate19400(.O (I18587), .I1 (g2370), .I2 (g14679));
ND4X1 gate19401(.O (g21603), .I1 (g17872), .I2 (g14987), .I3 (g17723), .I4 (g17689));
ND2X1 gate19402(.O (I14853), .I1 (g9433), .I2 (g5142));
ND2X1 gate19403(.O (g27550), .I1 (g24943), .I2 (g25772));
ND2X1 gate19404(.O (g9485), .I1 (g1657), .I2 (g1624));
ND2X1 gate19405(.O (g14069), .I1 (g11653), .I2 (g8864));
ND2X1 gate19406(.O (g22668), .I1 (g20219), .I2 (g2912));
ND2X1 gate19407(.O (g10602), .I1 (g7411), .I2 (g7451));
ND3X1 gate19408(.O (g11446), .I1 (g8700), .I2 (g6941), .I3 (g8734));
ND2X1 gate19409(.O (g14810), .I1 (g12700), .I2 (g10312));
ND2X1 gate19410(.O (g15033), .I1 (g12806), .I2 (g7142));
ND2X1 gate19411(.O (g12287), .I1 (g8381), .I2 (g2587));
ND4X1 gate19412(.O (g21429), .I1 (g17788), .I2 (g14803), .I3 (g17578), .I4 (g17520));
ND4X1 gate19413(.O (g17669), .I1 (g3570), .I2 (g11238), .I3 (g3632), .I4 (g13902));
ND2X1 gate19414(.O (g12307), .I1 (g7395), .I2 (g5983));
ND2X1 gate19415(.O (g14879), .I1 (g12646), .I2 (g10266));
ND2X1 gate19416(.O (I13066), .I1 (g4308), .I2 (I13065));
ND4X1 gate19417(.O (g17668), .I1 (g3235), .I2 (g13765), .I3 (g3310), .I4 (g13877));
ND2X1 gate19418(.O (g23428), .I1 (g13945), .I2 (g20522));
ND2X1 gate19419(.O (g13058), .I1 (g10544), .I2 (g1312));
ND3X1 gate19420(.O (g28977), .I1 (g27937), .I2 (g2629), .I3 (g2555));
ND2X1 gate19421(.O (g12431), .I1 (I15254), .I2 (I15255));
ND2X1 gate19422(.O (g20979), .I1 (g5385), .I2 (g17309));
ND3X1 gate19423(.O (g28783), .I1 (g27779), .I2 (g7315), .I3 (g1728));
ND2X1 gate19424(.O (g20055), .I1 (g11269), .I2 (g17794));
ND4X1 gate19425(.O (g20111), .I1 (g17513), .I2 (g14517), .I3 (g17468), .I4 (g14422));
ND2X1 gate19426(.O (g17525), .I1 (g14600), .I2 (g14574));
ND2X1 gate19427(.O (I13511), .I1 (g2093), .I2 (I13509));
ND2X1 gate19428(.O (g12341), .I1 (g7512), .I2 (g5308));
ND2X1 gate19429(.O (g28823), .I1 (g27738), .I2 (g14565));
ND2X1 gate19430(.O (I14276), .I1 (g8218), .I2 (I14275));
ND2X1 gate19431(.O (I21976), .I1 (g7680), .I2 (g19620));
ND2X1 gate19432(.O (g16291), .I1 (g13551), .I2 (g13545));
ND2X1 gate19433(.O (I23985), .I1 (g22182), .I2 (g482));
ND2X1 gate19434(.O (g13281), .I1 (g10916), .I2 (g1099));
ND2X1 gate19435(.O (g27670), .I1 (g25172), .I2 (g26666));
ND2X1 gate19436(.O (g22713), .I1 (g20114), .I2 (g2890));
ND2X1 gate19437(.O (g11957), .I1 (g8205), .I2 (g8259));
ND4X1 gate19438(.O (g28336), .I1 (g27064), .I2 (g24756), .I3 (g27163), .I4 (g19644));
ND2X1 gate19439(.O (I32202), .I1 (g33937), .I2 (g33670));
ND2X1 gate19440(.O (g13739), .I1 (g11773), .I2 (g11261));
ND3X1 gate19441(.O (g25396), .I1 (g22384), .I2 (g2208), .I3 (g8259));
ND3X1 gate19442(.O (g28966), .I1 (g27858), .I2 (g2361), .I3 (g7380));
ND2X1 gate19443(.O (g14918), .I1 (g12646), .I2 (g12772));
ND4X1 gate19444(.O (g20150), .I1 (g17705), .I2 (g17669), .I3 (g17635), .I4 (g14590));
ND2X1 gate19445(.O (g14079), .I1 (g11626), .I2 (g11763));
ND4X1 gate19446(.O (g17705), .I1 (g3586), .I2 (g13799), .I3 (g3661), .I4 (g13902));
ND2X1 gate19447(.O (g8292), .I1 (g218), .I2 (g215));
ND2X1 gate19448(.O (g14599), .I1 (g12207), .I2 (g9739));
ND2X1 gate19449(.O (I12253), .I1 (g1129), .I2 (I12251));
ND4X1 gate19450(.O (g17679), .I1 (g5611), .I2 (g14425), .I3 (g5681), .I4 (g12563));
ND2X1 gate19451(.O (g7869), .I1 (I12252), .I2 (I12253));
ND2X1 gate19452(.O (g10598), .I1 (g7191), .I2 (g6404));
ND4X1 gate19453(.O (g15788), .I1 (g6613), .I2 (g12211), .I3 (g6675), .I4 (g14786));
ND2X1 gate19454(.O (I18579), .I1 (g1945), .I2 (g14678));
ND4X1 gate19455(.O (g14598), .I1 (g5248), .I2 (g12002), .I3 (g5331), .I4 (g12497));
ND2X1 gate19456(.O (I14733), .I1 (g9732), .I2 (g5475));
ND2X1 gate19457(.O (g15829), .I1 (g4112), .I2 (g13831));
ND4X1 gate19458(.O (g17686), .I1 (g6251), .I2 (g14529), .I3 (g6322), .I4 (g12672));
ND2X1 gate19459(.O (I12372), .I1 (g3457), .I2 (g3462));
ND2X1 gate19460(.O (g14817), .I1 (g12711), .I2 (g12622));
ND3X1 gate19461(.O (g28288), .I1 (g10533), .I2 (g26105), .I3 (g27004));
ND2X1 gate19462(.O (g19913), .I1 (g11430), .I2 (g17794));
ND2X1 gate19463(.O (g19614), .I1 (g1542), .I2 (g16047));
ND2X1 gate19464(.O (g22875), .I1 (g20516), .I2 (g2980));
ND2X1 gate19465(.O (g25020), .I1 (g21377), .I2 (g23462));
ND2X1 gate19466(.O (g7442), .I1 (g896), .I2 (g890));
ND2X1 gate19467(.O (g24917), .I1 (g19913), .I2 (g23172));
ND2X1 gate19468(.O (g10561), .I1 (g7157), .I2 (g5712));
ND4X1 gate19469(.O (g27468), .I1 (g24951), .I2 (g24932), .I3 (g24925), .I4 (g26852));
ND2X1 gate19470(.O (I22921), .I1 (g14677), .I2 (g21284));
ND2X1 gate19471(.O (g27306), .I1 (g24787), .I2 (g26235));
ND2X1 gate19472(.O (g19530), .I1 (g15829), .I2 (g10841));
ND2X1 gate19473(.O (g12286), .I1 (I15129), .I2 (I15130));
ND2X1 gate19474(.O (g14656), .I1 (g12553), .I2 (g12405));
ND2X1 gate19475(.O (g9177), .I1 (g3355), .I2 (g3401));
ND2X1 gate19476(.O (g22837), .I1 (g20219), .I2 (g2907));
ND2X1 gate19477(.O (g12306), .I1 (g7394), .I2 (g5666));
ND2X1 gate19478(.O (I26461), .I1 (g14306), .I2 (I26459));
ND2X1 gate19479(.O (I24416), .I1 (g14382), .I2 (I24414));
ND4X1 gate19480(.O (g16604), .I1 (g3251), .I2 (g11194), .I3 (g3267), .I4 (g13877));
ND2X1 gate19481(.O (I22799), .I1 (g11960), .I2 (g21434));
ND4X1 gate19482(.O (g13551), .I1 (g11812), .I2 (g7479), .I3 (g7903), .I4 (g10521));
ND2X1 gate19483(.O (g10336), .I1 (I13750), .I2 (I13751));
ND2X1 gate19484(.O (g28976), .I1 (g27903), .I2 (g8273));
ND2X1 gate19485(.O (I14712), .I1 (g9671), .I2 (g5128));
ND2X1 gate19486(.O (I13335), .I1 (g1687), .I2 (I13334));
ND4X1 gate19487(.O (g16770), .I1 (g3263), .I2 (g13765), .I3 (g3274), .I4 (g8481));
ND2X1 gate19488(.O (g8561), .I1 (g3782), .I2 (g3774));
ND2X1 gate19489(.O (I22973), .I1 (g9657), .I2 (I22972));
ND2X1 gate19490(.O (g26248), .I1 (I25220), .I2 (I25221));
ND2X1 gate19491(.O (g12187), .I1 (I15042), .I2 (I15043));
ND2X1 gate19492(.O (I29262), .I1 (g29485), .I2 (I29261));
ND3X1 gate19493(.O (g11490), .I1 (g8666), .I2 (g3639), .I3 (g3694));
ND2X1 gate19494(.O (I26393), .I1 (g26488), .I2 (g14227));
NR2X1 gate19495(.O (g30249), .I1 (g5297), .I2 (g28982));
NR2X1 gate19496(.O (g33141), .I1 (g32099), .I2 (g8400));
NR2X1 gate19497(.O (g13824), .I1 (g8623), .I2 (g11702));
NR2X1 gate19498(.O (g27479), .I1 (g9056), .I2 (g26616));
NR2X1 gate19499(.O (g12479), .I1 (g2028), .I2 (g8310));
NR2X1 gate19500(.O (g20854), .I1 (g5381), .I2 (g17243));
NR2X1 gate19501(.O (g33135), .I1 (g32090), .I2 (g8350));
NR4X1 gate19502(.O (g7675), .I1 (g1554), .I2 (g1559), .I3 (g1564), .I4 (g1548));
NR4X1 gate19503(.O (g12486), .I1 (g9055), .I2 (g9013), .I3 (g8957), .I4 (g8905));
NR2X1 gate19504(.O (g9694), .I1 (g1936), .I2 (g1862));
NR2X1 gate19505(.O (g8906), .I1 (g3530), .I2 (g3522));
NR2X1 gate19506(.O (g14816), .I1 (g10166), .I2 (g12252));
NR2X1 gate19507(.O (g12223), .I1 (g2051), .I2 (g8365));
NR2X1 gate19508(.O (g14687), .I1 (g5352), .I2 (g12166));
NR2X1 gate19509(.O (g14752), .I1 (g12540), .I2 (g10040));
NR2X1 gate19510(.O (g16272), .I1 (g13580), .I2 (g11189));
NR2X1 gate19511(.O (g22524), .I1 (g19720), .I2 (g1361));
NR2X1 gate19512(.O (g25778), .I1 (g25459), .I2 (g25420));
NR2X1 gate19513(.O (g26212), .I1 (g23837), .I2 (g25408));
NR2X1 gate19514(.O (g17194), .I1 (g11039), .I2 (g13480));
NR2X1 gate19515(.O (g14392), .I1 (g12114), .I2 (g9537));
NR2X1 gate19516(.O (g13700), .I1 (g3288), .I2 (g11615));
NR2X1 gate19517(.O (g11658), .I1 (g8021), .I2 (g3506));
NR2X1 gate19518(.O (g15718), .I1 (g13858), .I2 (g11330));
NR3X1 gate19519(.O (g10488), .I1 (g4616), .I2 (g7133), .I3 (g10336));
NR3X1 gate19520(.O (g29107), .I1 (g6203), .I2 (g7791), .I3 (g26977));
NR3X1 gate19521(.O (g10893), .I1 (g1189), .I2 (g7715), .I3 (g7749));
NR2X1 gate19522(.O (g25932), .I1 (g7680), .I2 (g24528));
NR2X1 gate19523(.O (g29141), .I1 (g9374), .I2 (g27999));
NR2X1 gate19524(.O (g14713), .I1 (g12483), .I2 (g9974));
NR2X1 gate19525(.O (g31507), .I1 (g9064), .I2 (g29556));
NR2X1 gate19526(.O (g15099), .I1 (g13191), .I2 (g12869));
NR2X1 gate19527(.O (g11527), .I1 (g8165), .I2 (g8114));
NR3X1 gate19528(.O (g32715), .I1 (g31327), .I2 (I30261), .I3 (I30262));
NR2X1 gate19529(.O (g15098), .I1 (g13191), .I2 (g6927));
NR2X1 gate19530(.O (g30148), .I1 (g28799), .I2 (g7335));
NR2X1 gate19531(.O (g23602), .I1 (g9672), .I2 (g20979));
NR2X1 gate19532(.O (g28470), .I1 (g8021), .I2 (g27617));
NR2X1 gate19533(.O (g16220), .I1 (g13499), .I2 (g4939));
NR2X1 gate19534(.O (g14679), .I1 (g12437), .I2 (g9911));
NR2X1 gate19535(.O (g23955), .I1 (g2823), .I2 (g18890));
NR2X1 gate19536(.O (g33163), .I1 (g32099), .I2 (g7809));
NR2X1 gate19537(.O (g24619), .I1 (g23554), .I2 (g23581));
NR2X1 gate19538(.O (g14188), .I1 (g9162), .I2 (g12259));
NR2X1 gate19539(.O (g14124), .I1 (g8830), .I2 (g11083));
NR2X1 gate19540(.O (g14678), .I1 (g12432), .I2 (g9907));
NR2X1 gate19541(.O (g16246), .I1 (g13551), .I2 (g11169));
NR2X1 gate19542(.O (g12117), .I1 (g10113), .I2 (g9755));
NR2X1 gate19543(.O (g29361), .I1 (g7553), .I2 (g28174));
NR2X1 gate19544(.O (g15140), .I1 (g12887), .I2 (g13680));
NR2X1 gate19545(.O (g14093), .I1 (g8833), .I2 (g11083));
NR2X1 gate19546(.O (g15061), .I1 (g6815), .I2 (g13394));
NR3X1 gate19547(.O (g13910), .I1 (g4899), .I2 (g4975), .I3 (g11173));
NR2X1 gate19548(.O (g13202), .I1 (g8347), .I2 (g10511));
NR2X1 gate19549(.O (g12123), .I1 (g6856), .I2 (g2748));
NR2X1 gate19550(.O (g27772), .I1 (g7297), .I2 (g25839));
NR2X1 gate19551(.O (g12772), .I1 (g5188), .I2 (g9300));
NR2X1 gate19552(.O (g31121), .I1 (g4776), .I2 (g29540));
NR2X1 gate19553(.O (g23918), .I1 (g2799), .I2 (g21382));
NR2X1 gate19554(.O (g15162), .I1 (g13809), .I2 (g12904));
NR2X1 gate19555(.O (g11384), .I1 (g8538), .I2 (g8540));
NR2X1 gate19556(.O (g23079), .I1 (g8390), .I2 (g19965));
NR2X1 gate19557(.O (g29106), .I1 (g9451), .I2 (g28020));
NR2X1 gate19558(.O (g13094), .I1 (g7487), .I2 (g10762));
NR2X1 gate19559(.O (g26603), .I1 (g24908), .I2 (g24900));
NR3X1 gate19560(.O (g29033), .I1 (g5511), .I2 (g7738), .I3 (g28010));
NR2X1 gate19561(.O (g15628), .I1 (g11907), .I2 (g14228));
NR3X1 gate19562(.O (g32520), .I1 (g31554), .I2 (I30054), .I3 (I30055));
NR2X1 gate19563(.O (g17239), .I1 (g11119), .I2 (g13518));
NR3X1 gate19564(.O (g31134), .I1 (g8033), .I2 (g29679), .I3 (g24732));
NR2X1 gate19565(.O (g33134), .I1 (g7686), .I2 (g32057));
NR2X1 gate19566(.O (g16227), .I1 (g1554), .I2 (g13574));
NR2X1 gate19567(.O (g27007), .I1 (g5706), .I2 (g25821));
NR2X1 gate19568(.O (g31506), .I1 (g4793), .I2 (g29540));
NR2X1 gate19569(.O (g15071), .I1 (g6831), .I2 (g13416));
NR2X1 gate19570(.O (g15147), .I1 (g13716), .I2 (g12892));
NR3X1 gate19571(.O (g15754), .I1 (g341), .I2 (g7440), .I3 (g13385));
NR2X1 gate19572(.O (g14037), .I1 (g8748), .I2 (g11083));
NR2X1 gate19573(.O (g15825), .I1 (g7666), .I2 (g13217));
NR2X1 gate19574(.O (g16044), .I1 (g10961), .I2 (g13861));
NR2X1 gate19575(.O (g27720), .I1 (g9253), .I2 (g25791));
NR2X1 gate19576(.O (g14419), .I1 (g12152), .I2 (g9546));
NR2X1 gate19577(.O (g29012), .I1 (g5863), .I2 (g28020));
NR2X1 gate19578(.O (g15151), .I1 (g13745), .I2 (g7027));
NR2X1 gate19579(.O (g14418), .I1 (g12151), .I2 (g9594));
NR2X1 gate19580(.O (g10266), .I1 (g5188), .I2 (g5180));
NR2X1 gate19581(.O (g25958), .I1 (g7779), .I2 (g24609));
NR3X1 gate19582(.O (g32296), .I1 (g9044), .I2 (g31509), .I3 (g12259));
NR2X1 gate19583(.O (g31491), .I1 (g8938), .I2 (g29725));
NR2X1 gate19584(.O (g11280), .I1 (g8647), .I2 (g3408));
NR2X1 gate19585(.O (g25944), .I1 (g7716), .I2 (g24591));
NR2X1 gate19586(.O (g29359), .I1 (g7528), .I2 (g28167));
NR2X1 gate19587(.O (g12806), .I1 (g9472), .I2 (g9407));
NR2X1 gate19588(.O (g14194), .I1 (g5029), .I2 (g10515));
NR2X1 gate19589(.O (g19413), .I1 (g17151), .I2 (g14221));
NR3X1 gate19590(.O (g24953), .I1 (g10262), .I2 (g23978), .I3 (g12259));
NR2X1 gate19591(.O (g15059), .I1 (g12839), .I2 (g13350));
NR2X1 gate19592(.O (g26298), .I1 (g8297), .I2 (g24825));
NR2X1 gate19593(.O (g30129), .I1 (g28739), .I2 (g14537));
NR2X1 gate19594(.O (g15058), .I1 (g12838), .I2 (g13350));
NR3X1 gate19595(.O (g11231), .I1 (g7928), .I2 (g4801), .I3 (g4793));
NR2X1 gate19596(.O (g17284), .I1 (g9253), .I2 (g14317));
NR2X1 gate19597(.O (g12193), .I1 (g2342), .I2 (g8316));
NR2X1 gate19598(.O (g11885), .I1 (g7153), .I2 (g7167));
NR3X1 gate19599(.O (g29173), .I1 (g9259), .I2 (g27999), .I3 (g7704));
NR2X1 gate19600(.O (g14313), .I1 (g12016), .I2 (g9250));
NR2X1 gate19601(.O (g28476), .I1 (g27627), .I2 (g26547));
NR2X1 gate19602(.O (g16226), .I1 (g8052), .I2 (g13545));
NR2X1 gate19603(.O (g11763), .I1 (g3881), .I2 (g8172));
NR2X1 gate19604(.O (g25504), .I1 (g22550), .I2 (g7222));
NR2X1 gate19605(.O (g15120), .I1 (g12873), .I2 (g13605));
NR3X1 gate19606(.O (g32910), .I1 (g31327), .I2 (I30468), .I3 (I30469));
NR2X1 gate19607(.O (g25317), .I1 (g9766), .I2 (g23782));
NR2X1 gate19608(.O (g10808), .I1 (g8509), .I2 (g7611));
NR2X1 gate19609(.O (g15146), .I1 (g13716), .I2 (g7003));
NR2X1 gate19610(.O (g14036), .I1 (g8725), .I2 (g11083));
NR2X1 gate19611(.O (g34737), .I1 (g34706), .I2 (g30003));
NR2X1 gate19612(.O (g12437), .I1 (g2319), .I2 (g8267));
NR2X1 gate19613(.O (g27703), .I1 (g9607), .I2 (g25791));
NR2X1 gate19614(.O (g20000), .I1 (g13661), .I2 (g16264));
NR2X1 gate19615(.O (g13480), .I1 (g3017), .I2 (g11858));
NR2X1 gate19616(.O (g14642), .I1 (g12374), .I2 (g9829));
NR2X1 gate19617(.O (g12347), .I1 (g9321), .I2 (g9274));
NR2X1 gate19618(.O (g14064), .I1 (g9214), .I2 (g12259));
NR2X1 gate19619(.O (g13076), .I1 (g7443), .I2 (g10741));
NR2X1 gate19620(.O (g33098), .I1 (g31997), .I2 (g4616));
NR3X1 gate19621(.O (g28519), .I1 (g8011), .I2 (g27602), .I3 (g10295));
NR4X1 gate19622(.O (g12821), .I1 (g7132), .I2 (g10223), .I3 (g7149), .I4 (g10261));
NR2X1 gate19623(.O (g27063), .I1 (g26485), .I2 (g26516));
NR2X1 gate19624(.O (g24751), .I1 (g3034), .I2 (g23105));
NR2X1 gate19625(.O (g29903), .I1 (g6928), .I2 (g28484));
NR2X1 gate19626(.O (g11773), .I1 (g8883), .I2 (g4785));
NR2X1 gate19627(.O (g27516), .I1 (g9180), .I2 (g26657));
NR2X1 gate19628(.O (g33140), .I1 (g7693), .I2 (g32072));
NR2X1 gate19629(.O (g13341), .I1 (g7863), .I2 (g10762));
NR2X1 gate19630(.O (g12137), .I1 (g6682), .I2 (g7097));
NR2X1 gate19631(.O (g13670), .I1 (g8123), .I2 (g10756));
NR3X1 gate19632(.O (g10555), .I1 (g7227), .I2 (g4601), .I3 (g4608));
NR2X1 gate19633(.O (g20841), .I1 (g17847), .I2 (g12027));
NR3X1 gate19634(.O (g23042), .I1 (g16581), .I2 (g19462), .I3 (g10685));
NR2X1 gate19635(.O (g14712), .I1 (g12479), .I2 (g9971));
NR2X1 gate19636(.O (g13335), .I1 (g7851), .I2 (g10741));
NR2X1 gate19637(.O (g19890), .I1 (g16987), .I2 (g8058));
NR2X1 gate19638(.O (g14914), .I1 (g12822), .I2 (g12797));
NR2X1 gate19639(.O (g24391), .I1 (g22190), .I2 (g14645));
NR2X1 gate19640(.O (g15127), .I1 (g12879), .I2 (g13605));
NR2X1 gate19641(.O (g30271), .I1 (g7041), .I2 (g29008));
NR2X1 gate19642(.O (g23124), .I1 (g8443), .I2 (g20011));
NR2X1 gate19643(.O (g23678), .I1 (g9809), .I2 (g21190));
NR2X1 gate19644(.O (g16024), .I1 (g14216), .I2 (g11890));
NR2X1 gate19645(.O (g12208), .I1 (g10096), .I2 (g5759));
NR2X1 gate19646(.O (g33447), .I1 (g31978), .I2 (g7643));
NR2X1 gate19647(.O (g26330), .I1 (g8631), .I2 (g24825));
NR2X1 gate19648(.O (g23686), .I1 (g2767), .I2 (g21066));
NR2X1 gate19649(.O (g20014), .I1 (g17096), .I2 (g11244));
NR2X1 gate19650(.O (g33162), .I1 (g4859), .I2 (g32072));
NR2X1 gate19651(.O (g29898), .I1 (g6895), .I2 (g28458));
NR2X1 gate19652(.O (g12453), .I1 (g9444), .I2 (g5527));
NR2X1 gate19653(.O (g15095), .I1 (g13177), .I2 (g12866));
NR2X1 gate19654(.O (g29191), .I1 (g7738), .I2 (g28010));
NR2X1 gate19655(.O (g19778), .I1 (g16268), .I2 (g1061));
NR2X1 gate19656(.O (g11618), .I1 (g8114), .I2 (g8070));
NR2X1 gate19657(.O (g14382), .I1 (g9390), .I2 (g11139));
NR2X1 gate19658(.O (g14176), .I1 (g9044), .I2 (g12259));
NR2X1 gate19659(.O (g14092), .I1 (g8774), .I2 (g11083));
NR2X1 gate19660(.O (g19999), .I1 (g16232), .I2 (g13742));
NR2X1 gate19661(.O (g22400), .I1 (g19345), .I2 (g15718));
NR2X1 gate19662(.O (g20720), .I1 (g17847), .I2 (g9299));
NR3X1 gate19663(.O (g11469), .I1 (g650), .I2 (g9903), .I3 (g645));
NR2X1 gate19664(.O (g12593), .I1 (g9234), .I2 (g5164));
NR2X1 gate19665(.O (g12346), .I1 (g9931), .I2 (g9933));
NR3X1 gate19666(.O (g24720), .I1 (g1322), .I2 (g23051), .I3 (g19793));
NR2X1 gate19667(.O (g11039), .I1 (g9056), .I2 (g9092));
NR2X1 gate19668(.O (g11306), .I1 (g3412), .I2 (g8647));
NR2X1 gate19669(.O (g30132), .I1 (g28789), .I2 (g7362));
NR2X1 gate19670(.O (g22539), .I1 (g1030), .I2 (g19699));
NR2X1 gate19671(.O (g8958), .I1 (g3881), .I2 (g3873));
NR2X1 gate19672(.O (g33147), .I1 (g32090), .I2 (g7788));
NR2X1 gate19673(.O (g9061), .I1 (g3401), .I2 (g3361));
NR2X1 gate19674(.O (g19932), .I1 (g3376), .I2 (g16296));
NR2X1 gate19675(.O (g25887), .I1 (g24984), .I2 (g11706));
NR2X1 gate19676(.O (g15089), .I1 (g13144), .I2 (g12861));
NR2X1 gate19677(.O (g15088), .I1 (g13144), .I2 (g6874));
NR3X1 gate19678(.O (g13937), .I1 (g8883), .I2 (g4785), .I3 (g11155));
NR3X1 gate19679(.O (g21277), .I1 (g9417), .I2 (g9340), .I3 (g17467));
NR2X1 gate19680(.O (g29032), .I1 (g9300), .I2 (g27999));
NR2X1 gate19681(.O (g15126), .I1 (g12878), .I2 (g13605));
NR2X1 gate19682(.O (g11666), .I1 (g8172), .I2 (g8125));
NR2X1 gate19683(.O (g16581), .I1 (g13756), .I2 (g8086));
NR2X1 gate19684(.O (g11363), .I1 (g8626), .I2 (g8751));
NR2X1 gate19685(.O (g11217), .I1 (g8531), .I2 (g6875));
NR2X1 gate19686(.O (g31318), .I1 (g4785), .I2 (g29697));
NR2X1 gate19687(.O (g12711), .I1 (g6209), .I2 (g9326));
NR3X1 gate19688(.O (g8177), .I1 (g4966), .I2 (g4991), .I3 (g4983));
NR2X1 gate19689(.O (g30171), .I1 (g28880), .I2 (g7431));
NR2X1 gate19690(.O (g17515), .I1 (g13221), .I2 (g10828));
NR2X1 gate19691(.O (g15060), .I1 (g13350), .I2 (g6814));
NR3X1 gate19692(.O (g12492), .I1 (g7704), .I2 (g5170), .I3 (g5164));
NR2X1 gate19693(.O (g26545), .I1 (g24881), .I2 (g24855));
NR2X1 gate19694(.O (g27982), .I1 (g7212), .I2 (g25856));
NR2X1 gate19695(.O (g27381), .I1 (g8075), .I2 (g26657));
NR2X1 gate19696(.O (g14415), .I1 (g12147), .I2 (g9590));
NR2X1 gate19697(.O (g13110), .I1 (g7841), .I2 (g10741));
NR3X1 gate19698(.O (g26598), .I1 (g8990), .I2 (g13756), .I3 (g24732));
NR2X1 gate19699(.O (g33146), .I1 (g4669), .I2 (g32057));
NR2X1 gate19700(.O (g29071), .I1 (g5873), .I2 (g28020));
NR2X1 gate19701(.O (g29370), .I1 (g28585), .I2 (g28599));
NR2X1 gate19702(.O (g33427), .I1 (g10278), .I2 (g31950));
NR2X1 gate19703(.O (g22399), .I1 (g1367), .I2 (g19720));
NR2X1 gate19704(.O (g10312), .I1 (g5881), .I2 (g5873));
NR2X1 gate19705(.O (g15055), .I1 (g6808), .I2 (g13350));
NR2X1 gate19706(.O (g15070), .I1 (g6829), .I2 (g13416));
NR2X1 gate19707(.O (g30159), .I1 (g28799), .I2 (g14589));
NR2X1 gate19708(.O (g23560), .I1 (g9607), .I2 (g20838));
NR2X1 gate19709(.O (g12483), .I1 (g2453), .I2 (g8324));
NR2X1 gate19710(.O (g11216), .I1 (g7998), .I2 (g8037));
NR2X1 gate19711(.O (g10799), .I1 (g347), .I2 (g7541));
NR2X1 gate19712(.O (g12553), .I1 (g5170), .I2 (g9206));
NR2X1 gate19713(.O (g23642), .I1 (g9733), .I2 (g21124));
NR2X1 gate19714(.O (g15067), .I1 (g12842), .I2 (g13394));
NR2X1 gate19715(.O (g15094), .I1 (g13177), .I2 (g12865));
NR2X1 gate19716(.O (g30144), .I1 (g28789), .I2 (g7322));
NR2X1 gate19717(.O (g24453), .I1 (g7446), .I2 (g22325));
NR2X1 gate19718(.O (g15150), .I1 (g12895), .I2 (g13745));
NR2X1 gate19719(.O (g31127), .I1 (g4966), .I2 (g29556));
NR3X1 gate19720(.O (g13908), .I1 (g4709), .I2 (g8796), .I3 (g11155));
NR2X1 gate19721(.O (g12252), .I1 (g9995), .I2 (g10185));
NR2X1 gate19722(.O (g26309), .I1 (g8575), .I2 (g24825));
NR2X1 gate19723(.O (g11747), .I1 (g3530), .I2 (g8114));
NR2X1 gate19724(.O (g13568), .I1 (g8046), .I2 (g12527));
NR2X1 gate19725(.O (g16066), .I1 (g10929), .I2 (g13307));
NR2X1 gate19726(.O (g16231), .I1 (g13515), .I2 (g4771));
NR2X1 gate19727(.O (g33103), .I1 (g32176), .I2 (g31212));
NR2X1 gate19728(.O (g19793), .I1 (g16292), .I2 (g1404));
NR2X1 gate19729(.O (g33095), .I1 (g31997), .I2 (g7236));
NR2X1 gate19730(.O (g12847), .I1 (g6838), .I2 (g10430));
NR2X1 gate19731(.O (g25144), .I1 (g5046), .I2 (g23623));
NR2X1 gate19732(.O (g13772), .I1 (g3990), .I2 (g11702));
NR2X1 gate19733(.O (g28515), .I1 (g3881), .I2 (g27635));
NR2X1 gate19734(.O (g28414), .I1 (g27467), .I2 (g26347));
NR2X1 gate19735(.O (g30288), .I1 (g7087), .I2 (g29073));
NR2X1 gate19736(.O (g26976), .I1 (g5016), .I2 (g25791));
NR2X1 gate19737(.O (g29146), .I1 (g6565), .I2 (g26994));
NR2X1 gate19738(.O (g12851), .I1 (g6846), .I2 (g10430));
NR2X1 gate19739(.O (g14539), .I1 (g11977), .I2 (g9833));
NR2X1 gate19740(.O (g9649), .I1 (g2227), .I2 (g2153));
NR2X1 gate19741(.O (g14538), .I1 (g11973), .I2 (g9828));
NR2X1 gate19742(.O (g28584), .I1 (g7121), .I2 (g27635));
NR2X1 gate19743(.O (g16287), .I1 (g13622), .I2 (g11144));
NR2X1 gate19744(.O (g33089), .I1 (g31978), .I2 (g4322));
NR2X1 gate19745(.O (g15102), .I1 (g14591), .I2 (g6954));
NR2X1 gate19746(.O (g15157), .I1 (g13782), .I2 (g12900));
NR2X1 gate19747(.O (g33088), .I1 (g31997), .I2 (g7224));
NR2X1 gate19748(.O (g22514), .I1 (g19699), .I2 (g1018));
NR2X1 gate19749(.O (g12311), .I1 (g6109), .I2 (g10136));
NR2X1 gate19750(.O (g15066), .I1 (g12841), .I2 (g13394));
NR2X1 gate19751(.O (g24575), .I1 (g23498), .I2 (g23514));
NR2X1 gate19752(.O (g30260), .I1 (g7018), .I2 (g28982));
NR2X1 gate19753(.O (g23883), .I1 (g2779), .I2 (g21067));
NR2X1 gate19754(.O (g26865), .I1 (g25328), .I2 (g25290));
NR2X1 gate19755(.O (g31126), .I1 (g7928), .I2 (g29540));
NR2X1 gate19756(.O (g16268), .I1 (g7913), .I2 (g13121));
NR2X1 gate19757(.O (g12780), .I1 (g9402), .I2 (g9326));
NR2X1 gate19758(.O (g14515), .I1 (g12225), .I2 (g9761));
NR2X1 gate19759(.O (g14414), .I1 (g12145), .I2 (g9639));
NR2X1 gate19760(.O (g11493), .I1 (g8964), .I2 (g8967));
NR2X1 gate19761(.O (g25954), .I1 (g7750), .I2 (g24591));
NR2X1 gate19762(.O (g23729), .I1 (g17482), .I2 (g21206));
NR2X1 gate19763(.O (g20982), .I1 (g17929), .I2 (g12065));
NR2X1 gate19764(.O (g19880), .I1 (g16201), .I2 (g13634));
NR2X1 gate19765(.O (g27731), .I1 (g9229), .I2 (g25791));
NR2X1 gate19766(.O (g12846), .I1 (g6837), .I2 (g10430));
NR2X1 gate19767(.O (g22535), .I1 (g19699), .I2 (g1030));
NR2X1 gate19768(.O (g13806), .I1 (g11245), .I2 (g4076));
NR2X1 gate19769(.O (g29889), .I1 (g6905), .I2 (g28471));
NR2X1 gate19770(.O (g26686), .I1 (g23678), .I2 (g25189));
NR2X1 gate19771(.O (g13517), .I1 (g8541), .I2 (g12692));
NR2X1 gate19772(.O (g20390), .I1 (g17182), .I2 (g14257));
NR2X1 gate19773(.O (g29181), .I1 (g6573), .I2 (g26994));
NR2X1 gate19774(.O (g21284), .I1 (g16646), .I2 (g9690));
NR2X1 gate19775(.O (g26267), .I1 (g8033), .I2 (g24732));
NR2X1 gate19776(.O (g12405), .I1 (g9374), .I2 (g5180));
NR2X1 gate19777(.O (g16210), .I1 (g13479), .I2 (g4894));
NR2X1 gate19778(.O (g15054), .I1 (g12837), .I2 (g13350));
NR2X1 gate19779(.O (g27046), .I1 (g7544), .I2 (g25888));
NR2X1 gate19780(.O (g15156), .I1 (g13782), .I2 (g7050));
NR2X1 gate19781(.O (g30294), .I1 (g7110), .I2 (g29110));
NR2X1 gate19782(.O (g12046), .I1 (g10036), .I2 (g9640));
NR2X1 gate19783(.O (g14399), .I1 (g5297), .I2 (g12598));
NR2X1 gate19784(.O (g11006), .I1 (g7686), .I2 (g7836));
NR2X1 gate19785(.O (g12113), .I1 (g1648), .I2 (g8187));
NR2X1 gate19786(.O (g28106), .I1 (g7812), .I2 (g26994));
NR2X1 gate19787(.O (g25189), .I1 (g6082), .I2 (g23726));
NR2X1 gate19788(.O (g27827), .I1 (g9456), .I2 (g25839));
NR2X1 gate19789(.O (g9586), .I1 (g1668), .I2 (g1592));
NR2X1 gate19790(.O (g19887), .I1 (g3025), .I2 (g16275));
NR2X1 gate19791(.O (g29497), .I1 (g22763), .I2 (g28241));
NR2X1 gate19792(.O (g27769), .I1 (g9434), .I2 (g25805));
NR2X1 gate19793(.O (g15131), .I1 (g12881), .I2 (g13638));
NR2X1 gate19794(.O (g27768), .I1 (g9264), .I2 (g25805));
NR2X1 gate19795(.O (g30160), .I1 (g28846), .I2 (g7387));
NR2X1 gate19796(.O (g33094), .I1 (g31950), .I2 (g4639));
NR2X1 gate19797(.O (g14361), .I1 (g12079), .I2 (g9413));
NR2X1 gate19798(.O (g20183), .I1 (g17152), .I2 (g14222));
NR2X1 gate19799(.O (g28514), .I1 (g8165), .I2 (g27617));
NR2X1 gate19800(.O (g22491), .I1 (g1361), .I2 (g19720));
NR2X1 gate19801(.O (g16479), .I1 (g14719), .I2 (g12490));
NR2X1 gate19802(.O (g27027), .I1 (g26398), .I2 (g26484));
NR2X1 gate19803(.O (g24508), .I1 (g23577), .I2 (g23618));
NR2X1 gate19804(.O (g23052), .I1 (g8334), .I2 (g19916));
NR2X1 gate19805(.O (g12662), .I1 (g5863), .I2 (g9274));
NR2X1 gate19806(.O (g25160), .I1 (g5390), .I2 (g23659));
NR2X1 gate19807(.O (g12249), .I1 (g5763), .I2 (g10096));
NR2X1 gate19808(.O (g11834), .I1 (g8938), .I2 (g8822));
NR2X1 gate19809(.O (g12204), .I1 (g9927), .I2 (g10160));
NR2X1 gate19810(.O (g15143), .I1 (g6998), .I2 (g13680));
NR2X1 gate19811(.O (g30170), .I1 (g28846), .I2 (g14615));
NR2X1 gate19812(.O (g29503), .I1 (g22763), .I2 (g28250));
NR2X1 gate19813(.O (g14033), .I1 (g8808), .I2 (g12259));
NR2X1 gate19814(.O (g12081), .I1 (g10079), .I2 (g9694));
NR2X1 gate19815(.O (g13021), .I1 (g7544), .I2 (g10741));
NR2X1 gate19816(.O (g22521), .I1 (g1036), .I2 (g19699));
NR2X1 gate19817(.O (g27647), .I1 (g3004), .I2 (g26616));
NR2X1 gate19818(.O (g11913), .I1 (g7197), .I2 (g9166));
NR2X1 gate19819(.O (g13913), .I1 (g8859), .I2 (g11083));
NR2X1 gate19820(.O (g27356), .I1 (g9429), .I2 (g26657));
NR2X1 gate19821(.O (g7601), .I1 (g1322), .I2 (g1333));
NR2X1 gate19822(.O (g15168), .I1 (g13835), .I2 (g12909));
NR2X1 gate19823(.O (g27826), .I1 (g9501), .I2 (g25821));
NR2X1 gate19824(.O (g29910), .I1 (g3990), .I2 (g28484));
NR3X1 gate19825(.O (g11607), .I1 (g8848), .I2 (g8993), .I3 (g376));
NR2X1 gate19826(.O (g14514), .I1 (g11959), .I2 (g9760));
NR2X1 gate19827(.O (g11346), .I1 (g7980), .I2 (g7964));
NR3X1 gate19828(.O (g29070), .I1 (g5857), .I2 (g7766), .I3 (g28020));
NR2X1 gate19829(.O (g12651), .I1 (g9269), .I2 (g5511));
NR2X1 gate19830(.O (g10421), .I1 (g6227), .I2 (g9518));
NR2X1 gate19831(.O (g30119), .I1 (g28761), .I2 (g7315));
NR2X1 gate19832(.O (g14163), .I1 (g8997), .I2 (g12259));
NR2X1 gate19833(.O (g11797), .I1 (g8883), .I2 (g8796));
NR2X1 gate19834(.O (g19919), .I1 (g16987), .I2 (g11205));
NR2X1 gate19835(.O (g30276), .I1 (g7074), .I2 (g29073));
NR2X1 gate19836(.O (g30285), .I1 (g7097), .I2 (g29110));
NR2X1 gate19837(.O (g19444), .I1 (g17192), .I2 (g14295));
NR2X1 gate19838(.O (g12505), .I1 (g9444), .I2 (g9381));
NR2X1 gate19839(.O (g27717), .I1 (g9492), .I2 (g26745));
NR2X1 gate19840(.O (g9100), .I1 (g3752), .I2 (g3712));
NR2X1 gate19841(.O (g12026), .I1 (g9417), .I2 (g9340));
NR2X1 gate19842(.O (g8984), .I1 (g4899), .I2 (g4975));
NR2X1 gate19843(.O (g14121), .I1 (g8891), .I2 (g12259));
NR2X1 gate19844(.O (g25022), .I1 (g714), .I2 (g23324));
NR2X1 gate19845(.O (g11891), .I1 (g812), .I2 (g9166));
NR2X1 gate19846(.O (g16242), .I1 (g13529), .I2 (g4961));
NR2X1 gate19847(.O (g28491), .I1 (g8114), .I2 (g27617));
NR2X1 gate19848(.O (g33085), .I1 (g31978), .I2 (g4311));
NR2X1 gate19849(.O (g14291), .I1 (g9839), .I2 (g12155));
NR2X1 gate19850(.O (g11537), .I1 (g8229), .I2 (g3873));
NR2X1 gate19851(.O (g27343), .I1 (g8005), .I2 (g26616));
NR2X1 gate19852(.O (g28981), .I1 (g9234), .I2 (g27999));
NR2X1 gate19853(.O (g29077), .I1 (g6555), .I2 (g26994));
NR2X1 gate19854(.O (g12646), .I1 (g9234), .I2 (g9206));
NR3X1 gate19855(.O (g11283), .I1 (g7953), .I2 (g4991), .I3 (g9064));
NR2X1 gate19856(.O (g10760), .I1 (g1046), .I2 (g7479));
NR2X1 gate19857(.O (g11303), .I1 (g8497), .I2 (g8500));
NR2X1 gate19858(.O (g31942), .I1 (g8977), .I2 (g30583));
NR2X1 gate19859(.O (g27368), .I1 (g8119), .I2 (g26657));
NR2X1 gate19860(.O (g21206), .I1 (g6419), .I2 (g17396));
NR2X1 gate19861(.O (g12850), .I1 (g10430), .I2 (g6845));
NR2X1 gate19862(.O (g13796), .I1 (g9158), .I2 (g12527));
NR2X1 gate19863(.O (g28521), .I1 (g27649), .I2 (g26604));
NR2X1 gate19864(.O (g31965), .I1 (g30583), .I2 (g4358));
NR2X1 gate19865(.O (g33131), .I1 (g4659), .I2 (g32057));
NR4X1 gate19866(.O (g12228), .I1 (g10222), .I2 (g10206), .I3 (g10184), .I4 (g10335));
NR2X1 gate19867(.O (g10649), .I1 (g1183), .I2 (g8407));
NR3X1 gate19868(.O (g12716), .I1 (g7812), .I2 (g6555), .I3 (g6549));
NR2X1 gate19869(.O (g15123), .I1 (g6975), .I2 (g13605));
NR2X1 gate19870(.O (g10491), .I1 (g6573), .I2 (g9576));
NR2X1 gate19871(.O (g20027), .I1 (g16242), .I2 (g13779));
NR2X1 gate19872(.O (g21652), .I1 (g17619), .I2 (g17663));
NR2X1 gate19873(.O (g27379), .I1 (g8492), .I2 (g26636));
NR2X1 gate19874(.O (g11483), .I1 (g8165), .I2 (g3522));
NR2X1 gate19875(.O (g31469), .I1 (g8822), .I2 (g29725));
NR2X1 gate19876(.O (g11862), .I1 (g7134), .I2 (g7150));
NR2X1 gate19877(.O (g12050), .I1 (g10038), .I2 (g9649));
NR2X1 gate19878(.O (g24779), .I1 (g3736), .I2 (g23167));
NR2X1 gate19879(.O (g16237), .I1 (g8088), .I2 (g13574));
NR3X1 gate19880(.O (g29916), .I1 (g8681), .I2 (g28504), .I3 (g11083));
NR2X1 gate19881(.O (g23135), .I1 (g16476), .I2 (g19981));
NR2X1 gate19882(.O (g15992), .I1 (g10929), .I2 (g13846));
NR2X1 gate19883(.O (g28462), .I1 (g3512), .I2 (g27617));
NR2X1 gate19884(.O (g13326), .I1 (g10929), .I2 (g10905));
NR2X1 gate19885(.O (g14767), .I1 (g10130), .I2 (g12204));
NR2X1 gate19886(.O (g14395), .I1 (g12118), .I2 (g9542));
NR2X1 gate19887(.O (g17420), .I1 (g9456), .I2 (g14408));
NR2X1 gate19888(.O (g10899), .I1 (g4064), .I2 (g8451));
NR2X1 gate19889(.O (g22540), .I1 (g19720), .I2 (g1373));
NR2X1 gate19890(.O (g11252), .I1 (g8620), .I2 (g3057));
NR2X1 gate19891(.O (g11621), .I1 (g3512), .I2 (g7985));
NR2X1 gate19892(.O (g15578), .I1 (g7216), .I2 (g14279));
NR2X1 gate19893(.O (g20998), .I1 (g18065), .I2 (g9450));
NR2X1 gate19894(.O (g33143), .I1 (g32293), .I2 (g31518));
NR4X1 gate19895(.O (g7661), .I1 (g1211), .I2 (g1216), .I3 (g1221), .I4 (g1205));
NR2X1 gate19896(.O (g29180), .I1 (g9569), .I2 (g26977));
NR2X1 gate19897(.O (g14247), .I1 (g9934), .I2 (g10869));
NR2X1 gate19898(.O (g13872), .I1 (g8745), .I2 (g11083));
NR2X1 gate19899(.O (g25501), .I1 (g23918), .I2 (g14645));
NR2X1 gate19900(.O (g20717), .I1 (g5037), .I2 (g17217));
NR2X1 gate19901(.O (g14272), .I1 (g6411), .I2 (g10598));
NR2X1 gate19902(.O (g12129), .I1 (g9992), .I2 (g7051));
NR2X1 gate19903(.O (g12002), .I1 (g5297), .I2 (g7004));
NR3X1 gate19904(.O (g11213), .I1 (g4776), .I2 (g7892), .I3 (g9030));
NR2X1 gate19905(.O (g15142), .I1 (g13680), .I2 (g12889));
NR2X1 gate19906(.O (g33084), .I1 (g31978), .I2 (g7655));
NR2X1 gate19907(.O (g20149), .I1 (g17091), .I2 (g14185));
NR2X1 gate19908(.O (g26609), .I1 (g146), .I2 (g24732));
NR2X1 gate19909(.O (g15130), .I1 (g13638), .I2 (g6985));
NR2X1 gate19910(.O (g24148), .I1 (g19268), .I2 (g19338));
NR2X1 gate19911(.O (g15165), .I1 (g12907), .I2 (g13835));
NR2X1 gate19912(.O (g31373), .I1 (g4975), .I2 (g29725));
NR2X1 gate19913(.O (g11780), .I1 (g4899), .I2 (g8822));
NR2X1 gate19914(.O (g14360), .I1 (g12078), .I2 (g9484));
NR2X1 gate19915(.O (g9835), .I1 (g2629), .I2 (g2555));
NR2X1 gate19916(.O (g14447), .I1 (g11938), .I2 (g9698));
NR2X1 gate19917(.O (g12856), .I1 (g10430), .I2 (g6855));
NR2X1 gate19918(.O (g29187), .I1 (g7704), .I2 (g27999));
NR3X1 gate19919(.O (g11846), .I1 (g7635), .I2 (g7518), .I3 (g7548));
NR2X1 gate19920(.O (g16209), .I1 (g13478), .I2 (g4749));
NR2X1 gate19921(.O (g14911), .I1 (g10213), .I2 (g12364));
NR2X1 gate19922(.O (g27499), .I1 (g9095), .I2 (g26636));
NR3X1 gate19923(.O (g28540), .I1 (g8125), .I2 (g27635), .I3 (g7121));
NR2X1 gate19924(.O (g15372), .I1 (g817), .I2 (g14279));
NR2X1 gate19925(.O (g14754), .I1 (g12821), .I2 (g2988));
NR2X1 gate19926(.O (g27722), .I1 (g7247), .I2 (g25805));
NR2X1 gate19927(.O (g31117), .I1 (g4991), .I2 (g29556));
NR2X1 gate19928(.O (g27924), .I1 (g9946), .I2 (g25839));
NR2X1 gate19929(.O (g33117), .I1 (g31261), .I2 (g32205));
NR2X1 gate19930(.O (g22190), .I1 (g2827), .I2 (g18949));
NR2X1 gate19931(.O (g8720), .I1 (g358), .I2 (g365));
NR2X1 gate19932(.O (g15063), .I1 (g6818), .I2 (g13394));
NR2X1 gate19933(.O (g30934), .I1 (g29836), .I2 (g29850));
NR2X1 gate19934(.O (g19984), .I1 (g17096), .I2 (g8171));
NR2X1 gate19935(.O (g15137), .I1 (g6992), .I2 (g13680));
NR2X1 gate19936(.O (g12432), .I1 (g1894), .I2 (g8249));
NR2X1 gate19937(.O (g24959), .I1 (g8858), .I2 (g23324));
NR2X1 gate19938(.O (g17190), .I1 (g723), .I2 (g14279));
NR2X1 gate19939(.O (g14394), .I1 (g12116), .I2 (g9414));
NR2X1 gate19940(.O (g14367), .I1 (g9547), .I2 (g12289));
NR2X1 gate19941(.O (g16292), .I1 (g7943), .I2 (g13134));
NR2X1 gate19942(.O (g11357), .I1 (g8558), .I2 (g8561));
NR3X1 gate19943(.O (g29179), .I1 (g9311), .I2 (g28010), .I3 (g7738));
NR2X1 gate19944(.O (g14420), .I1 (g12153), .I2 (g9490));
NR2X1 gate19945(.O (g12198), .I1 (g9797), .I2 (g9800));
NR2X1 gate19946(.O (g19853), .I1 (g15746), .I2 (g1052));
NR3X1 gate19947(.O (g27528), .I1 (g8770), .I2 (g26352), .I3 (g11083));
NR2X1 gate19948(.O (g10318), .I1 (g25), .I2 (g22));
NR2X1 gate19949(.O (g14446), .I1 (g12190), .I2 (g9644));
NR2X1 gate19950(.O (g14227), .I1 (g9863), .I2 (g10838));
NR2X1 gate19951(.O (g20857), .I1 (g17929), .I2 (g9380));
NR2X1 gate19952(.O (g27960), .I1 (g7134), .I2 (g25791));
NR2X1 gate19953(.O (g14540), .I1 (g12287), .I2 (g9834));
NR2X1 gate19954(.O (g19401), .I1 (g17193), .I2 (g14296));
NR2X1 gate19955(.O (g17700), .I1 (g14792), .I2 (g12983));
NR2X1 gate19956(.O (g17625), .I1 (g14541), .I2 (g12123));
NR2X1 gate19957(.O (g15073), .I1 (g12844), .I2 (g13416));
NR3X1 gate19958(.O (g28481), .I1 (g3506), .I2 (g10323), .I3 (g27617));
NR2X1 gate19959(.O (g10281), .I1 (g5535), .I2 (g5527));
NR2X1 gate19960(.O (g15122), .I1 (g6959), .I2 (g13605));
NR2X1 gate19961(.O (g26515), .I1 (g24843), .I2 (g24822));
NR2X1 gate19962(.O (g12708), .I1 (g9518), .I2 (g9462));
NR2X1 gate19963(.O (g25005), .I1 (g6811), .I2 (g23324));
NR2X1 gate19964(.O (g10699), .I1 (g8526), .I2 (g1514));
NR2X1 gate19965(.O (g15153), .I1 (g13745), .I2 (g12897));
NR2X1 gate19966(.O (g31116), .I1 (g7892), .I2 (g29540));
NR3X1 gate19967(.O (g11248), .I1 (g7953), .I2 (g4991), .I3 (g4983));
NR3X1 gate19968(.O (g32780), .I1 (g31327), .I2 (I30330), .I3 (I30331));
NR2X1 gate19969(.O (g15136), .I1 (g13680), .I2 (g12885));
NR2X1 gate19970(.O (g29908), .I1 (g6918), .I2 (g28471));
NR2X1 gate19971(.O (g27879), .I1 (g9523), .I2 (g25856));
NR2X1 gate19972(.O (g22450), .I1 (g19345), .I2 (g15724));
NR3X1 gate19973(.O (g12970), .I1 (g10555), .I2 (g10510), .I3 (g10488));
NR2X1 gate19974(.O (g27878), .I1 (g9559), .I2 (g25839));
NR2X1 gate19975(.O (g27337), .I1 (g8334), .I2 (g26616));
NR2X1 gate19976(.O (g15164), .I1 (g13835), .I2 (g12906));
NR2X1 gate19977(.O (g11945), .I1 (g7212), .I2 (g7228));
NR2X1 gate19978(.O (g11999), .I1 (g9654), .I2 (g7423));
NR2X1 gate19979(.O (g10715), .I1 (g8526), .I2 (g8466));
NR3X1 gate19980(.O (g21389), .I1 (g10143), .I2 (g17748), .I3 (g12259));
NR2X1 gate19981(.O (g20995), .I1 (g5727), .I2 (g17287));
NR2X1 gate19982(.O (g28520), .I1 (g8229), .I2 (g27635));
NR2X1 gate19983(.O (g25407), .I1 (g23871), .I2 (g14645));
NR2X1 gate19984(.O (g27010), .I1 (g6052), .I2 (g25839));
NR2X1 gate19985(.O (g11932), .I1 (g843), .I2 (g9166));
NR2X1 gate19986(.O (g33130), .I1 (g32265), .I2 (g31497));
NR2X1 gate19987(.O (g11448), .I1 (g4191), .I2 (g8790));
NR2X1 gate19988(.O (g14490), .I1 (g9853), .I2 (g12598));
NR2X1 gate19989(.O (g19907), .I1 (g16210), .I2 (g13676));
NR2X1 gate19990(.O (g21140), .I1 (g6073), .I2 (g17312));
NR2X1 gate19991(.O (g15091), .I1 (g13177), .I2 (g12863));
NR2X1 gate19992(.O (g33437), .I1 (g31997), .I2 (g10275));
NR2X1 gate19993(.O (g29007), .I1 (g9269), .I2 (g28010));
NR2X1 gate19994(.O (g10671), .I1 (g1526), .I2 (g8466));
NR2X1 gate19995(.O (g14181), .I1 (g9083), .I2 (g12259));
NR2X1 gate19996(.O (g23871), .I1 (g2811), .I2 (g21348));
NR2X1 gate19997(.O (g27353), .I1 (g8097), .I2 (g26616));
NR2X1 gate19998(.O (g16183), .I1 (g9223), .I2 (g13545));
NR2X1 gate19999(.O (g27823), .I1 (g9792), .I2 (g25805));
NR4X1 gate20000(.O (g11148), .I1 (g8052), .I2 (g9197), .I3 (g9174), .I4 (g9050));
NR2X1 gate20001(.O (g12680), .I1 (g9631), .I2 (g9576));
NR2X1 gate20002(.O (g19935), .I1 (g17062), .I2 (g8113));
NR2X1 gate20003(.O (g31372), .I1 (g8796), .I2 (g29697));
NR2X1 gate20004(.O (g25141), .I1 (g22228), .I2 (g10334));
NR2X1 gate20005(.O (g33175), .I1 (g32099), .I2 (g7828));
NR2X1 gate20006(.O (g24145), .I1 (g19402), .I2 (g19422));
NR2X1 gate20007(.O (g27966), .I1 (g7153), .I2 (g25805));
NR3X1 gate20008(.O (g13971), .I1 (g8938), .I2 (g4975), .I3 (g11173));
NR2X1 gate20009(.O (g29035), .I1 (g9321), .I2 (g28020));
NR2X1 gate20010(.O (g14211), .I1 (g9779), .I2 (g10823));
NR2X1 gate20011(.O (g27364), .I1 (g8426), .I2 (g26616));
NR2X1 gate20012(.O (g33137), .I1 (g4849), .I2 (g32072));
NR2X1 gate20013(.O (g12017), .I1 (g9969), .I2 (g9586));
NR2X1 gate20014(.O (g12364), .I1 (g10102), .I2 (g10224));
NR2X1 gate20015(.O (g30613), .I1 (g4507), .I2 (g29365));
NR2X1 gate20016(.O (g29142), .I1 (g5535), .I2 (g28010));
NR2X1 gate20017(.O (g14497), .I1 (g5990), .I2 (g12705));
NR2X1 gate20018(.O (g30273), .I1 (g5990), .I2 (g29036));
NR2X1 gate20019(.O (g30106), .I1 (g28739), .I2 (g7268));
NR2X1 gate20020(.O (g12288), .I1 (g2610), .I2 (g8418));
NR3X1 gate20021(.O (g29193), .I1 (g9529), .I2 (g26994), .I3 (g7812));
NR2X1 gate20022(.O (g19906), .I1 (g16209), .I2 (g13672));
NR2X1 gate20023(.O (g12571), .I1 (g9511), .I2 (g9451));
NR2X1 gate20024(.O (g12308), .I1 (g9951), .I2 (g9954));
NR2X1 gate20025(.O (g25004), .I1 (g676), .I2 (g23324));
NR2X1 gate20026(.O (g28496), .I1 (g3179), .I2 (g27602));
NR2X1 gate20027(.O (g29165), .I1 (g5881), .I2 (g28020));
NR2X1 gate20028(.O (g14339), .I1 (g12289), .I2 (g2735));
NR2X1 gate20029(.O (g16072), .I1 (g10961), .I2 (g13273));
NR2X1 gate20030(.O (g10338), .I1 (g5062), .I2 (g5022));
NR2X1 gate20031(.O (g15062), .I1 (g6817), .I2 (g13394));
NR2X1 gate20032(.O (g28986), .I1 (g5517), .I2 (g28010));
NR2X1 gate20033(.O (g29006), .I1 (g5180), .I2 (g27999));
NR2X1 gate20034(.O (g25947), .I1 (g1199), .I2 (g24591));
NR2X1 gate20035(.O (g15508), .I1 (g10320), .I2 (g14279));
NR2X1 gate20036(.O (g13959), .I1 (g3698), .I2 (g11309));
NR2X1 gate20037(.O (g27954), .I1 (g10014), .I2 (g25856));
NR2X1 gate20038(.O (g12752), .I1 (g9576), .I2 (g9529));
NR2X1 gate20039(.O (g11958), .I1 (g9543), .I2 (g7327));
NR2X1 gate20040(.O (g12374), .I1 (g2185), .I2 (g8205));
NR2X1 gate20041(.O (g13378), .I1 (g11374), .I2 (g11017));
NR2X1 gate20042(.O (g14411), .I1 (g9460), .I2 (g11160));
NR2X1 gate20043(.O (g13603), .I1 (g8009), .I2 (g10721));
NR2X1 gate20044(.O (g13944), .I1 (g10262), .I2 (g12259));
NR2X1 gate20045(.O (g14867), .I1 (g10191), .I2 (g12314));
NR2X1 gate20046(.O (g14450), .I1 (g12195), .I2 (g9598));
NR2X1 gate20047(.O (g29175), .I1 (g6227), .I2 (g26977));
NR2X1 gate20048(.O (g10819), .I1 (g7479), .I2 (g1041));
NR2X1 gate20049(.O (g13730), .I1 (g3639), .I2 (g11663));
NR3X1 gate20050(.O (g34359), .I1 (g9162), .I2 (g34174), .I3 (g12259));
NR2X1 gate20051(.O (g14707), .I1 (g10143), .I2 (g12259));
NR2X1 gate20052(.O (g28457), .I1 (g7980), .I2 (g27602));
NR3X1 gate20053(.O (g32212), .I1 (g8859), .I2 (g31262), .I3 (g11083));
NR3X1 gate20054(.O (g12558), .I1 (g7738), .I2 (g5517), .I3 (g5511));
NR2X1 gate20055(.O (g13765), .I1 (g8531), .I2 (g11615));
NR2X1 gate20056(.O (g15051), .I1 (g6801), .I2 (g13350));
NR2X1 gate20057(.O (g15072), .I1 (g13416), .I2 (g12843));
NR2X1 gate20058(.O (g7192), .I1 (g6444), .I2 (g6404));
NR2X1 gate20059(.O (g29873), .I1 (g6875), .I2 (g28458));
NR2X1 gate20060(.O (g17180), .I1 (g1559), .I2 (g13574));
NR3X1 gate20061(.O (g22993), .I1 (g1322), .I2 (g16292), .I3 (g19873));
NR2X1 gate20062(.O (g14094), .I1 (g8770), .I2 (g11083));
NR2X1 gate20063(.O (g15152), .I1 (g13745), .I2 (g12896));
NR2X1 gate20064(.O (g33109), .I1 (g31997), .I2 (g4584));
NR2X1 gate20065(.O (g12189), .I1 (g1917), .I2 (g8302));
NR2X1 gate20066(.O (g13129), .I1 (g7553), .I2 (g10762));
NR2X1 gate20067(.O (g10801), .I1 (g1041), .I2 (g7479));
NR2X1 gate20068(.O (g17694), .I1 (g12435), .I2 (g12955));
NR2X1 gate20069(.O (g33108), .I1 (g32183), .I2 (g31228));
NR2X1 gate20070(.O (g30134), .I1 (g28768), .I2 (g7280));
NR3X1 gate20071(.O (g11626), .I1 (g7121), .I2 (g3863), .I3 (g3857));
NR2X1 gate20072(.O (g10695), .I1 (g8462), .I2 (g8407));
NR2X1 gate20073(.O (g27093), .I1 (g26712), .I2 (g26749));
NR2X1 gate20074(.O (g17619), .I1 (g10179), .I2 (g12955));
NR2X1 gate20075(.O (g12093), .I1 (g9924), .I2 (g7028));
NR2X1 gate20076(.O (g26649), .I1 (g9037), .I2 (g24732));
NR2X1 gate20077(.O (g27875), .I1 (g9875), .I2 (g25821));
NR2X1 gate20078(.O (g33174), .I1 (g8714), .I2 (g32072));
NR3X1 gate20079(.O (g11232), .I1 (g4966), .I2 (g7898), .I3 (g9064));
NR2X1 gate20080(.O (g29034), .I1 (g5527), .I2 (g28010));
NR2X1 gate20081(.O (g19400), .I1 (g17139), .I2 (g14206));
NR2X1 gate20082(.O (g21127), .I1 (g18065), .I2 (g12099));
NR2X1 gate20083(.O (g11697), .I1 (g8080), .I2 (g3857));
NR2X1 gate20084(.O (g11995), .I1 (g9645), .I2 (g7410));
NR2X1 gate20085(.O (g16027), .I1 (g10929), .I2 (g13260));
NR3X1 gate20086(.O (g11261), .I1 (g7928), .I2 (g4801), .I3 (g9030));
NR2X1 gate20087(.O (g14001), .I1 (g739), .I2 (g11083));
NR2X1 gate20088(.O (g30240), .I1 (g7004), .I2 (g28982));
NR4X1 gate20089(.O (g24631), .I1 (g20516), .I2 (g20436), .I3 (g20219), .I4 (g22957));
NR2X1 gate20090(.O (g12160), .I1 (g9721), .I2 (g9724));
NR2X1 gate20091(.O (g13512), .I1 (g9077), .I2 (g12527));
NR2X1 gate20092(.O (g28480), .I1 (g8059), .I2 (g27602));
NR4X1 gate20093(.O (g23956), .I1 (g18957), .I2 (g18918), .I3 (g20136), .I4 (g20114));
NR2X1 gate20094(.O (g8933), .I1 (g4709), .I2 (g4785));
NR2X1 gate20095(.O (g31483), .I1 (g4899), .I2 (g29725));
NR2X1 gate20096(.O (g13831), .I1 (g11245), .I2 (g7666));
NR2X1 gate20097(.O (g12201), .I1 (g5417), .I2 (g10047));
NR2X1 gate20098(.O (g29164), .I1 (g9444), .I2 (g28010));
NR2X1 gate20099(.O (g12467), .I1 (g9472), .I2 (g9407));
NR2X1 gate20100(.O (g30262), .I1 (g5644), .I2 (g29008));
NR2X1 gate20101(.O (g13989), .I1 (g8697), .I2 (g11309));
NR2X1 gate20102(.O (g13056), .I1 (g7400), .I2 (g10741));
NR2X1 gate20103(.O (g16090), .I1 (g10961), .I2 (g13315));
NR2X1 gate20104(.O (g26573), .I1 (g24897), .I2 (g24884));
NR2X1 gate20105(.O (g11924), .I1 (g7187), .I2 (g7209));
NR2X1 gate20106(.O (g29109), .I1 (g9472), .I2 (g26994));
NR2X1 gate20107(.O (g27352), .I1 (g7975), .I2 (g26616));
NR2X1 gate20108(.O (g26247), .I1 (g7995), .I2 (g24732));
NR2X1 gate20109(.O (g7781), .I1 (g4064), .I2 (g4057));
NR2X1 gate20110(.O (g12419), .I1 (g9402), .I2 (g9326));
NR2X1 gate20111(.O (g25770), .I1 (g25417), .I2 (g25377));
NR2X1 gate20112(.O (g29108), .I1 (g6219), .I2 (g26977));
NR2X1 gate20113(.O (g24976), .I1 (g671), .I2 (g23324));
NR2X1 gate20114(.O (g12418), .I1 (g9999), .I2 (g10001));
NR2X1 gate20115(.O (g12170), .I1 (g10047), .I2 (g5413));
NR2X1 gate20116(.O (g26098), .I1 (g9073), .I2 (g24732));
NR2X1 gate20117(.O (g23024), .I1 (g7936), .I2 (g19407));
NR2X1 gate20118(.O (g13342), .I1 (g10961), .I2 (g10935));
NR2X1 gate20119(.O (g13031), .I1 (g7301), .I2 (g10741));
NR2X1 gate20120(.O (g12853), .I1 (g6848), .I2 (g10430));
NR3X1 gate20121(.O (g33851), .I1 (g8854), .I2 (g33299), .I3 (g12259));
NR2X1 gate20122(.O (g29174), .I1 (g9511), .I2 (g28020));
NR3X1 gate20123(.O (g21250), .I1 (g9417), .I2 (g9340), .I3 (g17494));
NR2X1 gate20124(.O (g21658), .I1 (g17694), .I2 (g17727));
NR2X1 gate20125(.O (g22654), .I1 (g7733), .I2 (g19506));
NR2X1 gate20126(.O (g25521), .I1 (g23955), .I2 (g14645));
NR3X1 gate20127(.O (g11869), .I1 (g7649), .I2 (g7534), .I3 (g7581));
NR2X1 gate20128(.O (g15647), .I1 (g11924), .I2 (g14248));
NR2X1 gate20129(.O (g28469), .I1 (g3171), .I2 (g27602));
NR2X1 gate20130(.O (g15090), .I1 (g13144), .I2 (g12862));
NR3X1 gate20131(.O (g28468), .I1 (g3155), .I2 (g10295), .I3 (g27602));
NR2X1 gate20132(.O (g10341), .I1 (g6227), .I2 (g6219));
NR2X1 gate20133(.O (g25247), .I1 (g23763), .I2 (g14645));
NR2X1 gate20134(.O (g27704), .I1 (g7239), .I2 (g25791));
NR2X1 gate20135(.O (g11225), .I1 (g3990), .I2 (g6928));
NR2X1 gate20136(.O (g26162), .I1 (g23052), .I2 (g24751));
NR3X1 gate20137(.O (g16646), .I1 (g13437), .I2 (g11020), .I3 (g11372));
NR2X1 gate20138(.O (g12466), .I1 (g10057), .I2 (g10059));
NR2X1 gate20139(.O (g25777), .I1 (g25482), .I2 (g25456));
NR2X1 gate20140(.O (g14335), .I1 (g12045), .I2 (g9283));
NR2X1 gate20141(.O (g12101), .I1 (g6336), .I2 (g7074));
NR2X1 gate20142(.O (g26628), .I1 (g8990), .I2 (g24732));
NR2X1 gate20143(.O (g29040), .I1 (g6209), .I2 (g26977));
NR2X1 gate20144(.O (g30162), .I1 (g28880), .I2 (g7462));
NR2X1 gate20145(.O (g8864), .I1 (g3179), .I2 (g3171));
NR2X1 gate20146(.O (g24383), .I1 (g22409), .I2 (g22360));
NR2X1 gate20147(.O (g27733), .I1 (g9305), .I2 (g25805));
NR3X1 gate20148(.O (g13970), .I1 (g8883), .I2 (g8796), .I3 (g11155));
NR4X1 gate20149(.O (g11171), .I1 (g8088), .I2 (g9226), .I3 (g9200), .I4 (g9091));
NR3X1 gate20150(.O (g29183), .I1 (g9392), .I2 (g28020), .I3 (g7766));
NR3X1 gate20151(.O (g24875), .I1 (g8725), .I2 (g23850), .I3 (g11083));
NR2X1 gate20152(.O (g12166), .I1 (g9856), .I2 (g10124));
NR3X1 gate20153(.O (g14278), .I1 (g562), .I2 (g12259), .I3 (g9217));
NR2X1 gate20154(.O (g13994), .I1 (g4049), .I2 (g11363));
NR2X1 gate20155(.O (g15149), .I1 (g13745), .I2 (g12894));
NR2X1 gate20156(.O (g25447), .I1 (g23883), .I2 (g14645));
NR2X1 gate20157(.O (g14306), .I1 (g10060), .I2 (g10887));
NR3X1 gate20158(.O (g29933), .I1 (g8808), .I2 (g28500), .I3 (g12259));
NR2X1 gate20159(.O (g15148), .I1 (g13716), .I2 (g12893));
NR2X1 gate20160(.O (g15097), .I1 (g12868), .I2 (g13191));
NR2X1 gate20161(.O (g30147), .I1 (g28768), .I2 (g14567));
NR2X1 gate20162(.O (g13919), .I1 (g3347), .I2 (g11276));
NR2X1 gate20163(.O (g9755), .I1 (g2070), .I2 (g1996));
NR2X1 gate20164(.O (g13078), .I1 (g7446), .I2 (g10762));
NR2X1 gate20165(.O (g23695), .I1 (g17420), .I2 (g21140));
NR2X1 gate20166(.O (g19951), .I1 (g16219), .I2 (g13709));
NR3X1 gate20167(.O (g25776), .I1 (g7166), .I2 (g24380), .I3 (g24369));
NR2X1 gate20168(.O (g25785), .I1 (g25488), .I2 (g25462));
NR2X1 gate20169(.O (g10884), .I1 (g7650), .I2 (g8451));
NR2X1 gate20170(.O (g27382), .I1 (g8219), .I2 (g26657));
NR2X1 gate20171(.O (g28953), .I1 (g5170), .I2 (g27999));
NR2X1 gate20172(.O (g24494), .I1 (g23513), .I2 (g23532));
NR2X1 gate20173(.O (g15133), .I1 (g12883), .I2 (g13638));
NR3X1 gate20174(.O (g32650), .I1 (g31579), .I2 (I30192), .I3 (I30193));
NR2X1 gate20175(.O (g13125), .I1 (g7863), .I2 (g10762));
NR2X1 gate20176(.O (g10666), .I1 (g8462), .I2 (g1171));
NR2X1 gate20177(.O (g25950), .I1 (g1070), .I2 (g24591));
NR2X1 gate20178(.O (g7142), .I1 (g6573), .I2 (g6565));
NR2X1 gate20179(.O (g12154), .I1 (g10155), .I2 (g9835));
NR2X1 gate20180(.O (g29072), .I1 (g9402), .I2 (g26977));
NR4X1 gate20181(.O (g9602), .I1 (g4688), .I2 (g4681), .I3 (g4674), .I4 (g4646));
NR2X1 gate20182(.O (g14556), .I1 (g6682), .I2 (g12790));
NR2X1 gate20183(.O (g26645), .I1 (g23602), .I2 (g25160));
NR2X1 gate20184(.O (g13336), .I1 (g11330), .I2 (g11011));
NR2X1 gate20185(.O (g21256), .I1 (g15483), .I2 (g12179));
NR3X1 gate20186(.O (g22983), .I1 (g979), .I2 (g16268), .I3 (g19853));
NR2X1 gate20187(.O (g9015), .I1 (g3050), .I2 (g3010));
NR2X1 gate20188(.O (g15050), .I1 (g12834), .I2 (g13350));
NR2X1 gate20189(.O (g12729), .I1 (g1657), .I2 (g8139));
NR2X1 gate20190(.O (g13631), .I1 (g8068), .I2 (g10733));
NR2X1 gate20191(.O (g10922), .I1 (g7650), .I2 (g4057));
NR2X1 gate20192(.O (g25446), .I1 (g23686), .I2 (g14645));
NR2X1 gate20193(.O (g22517), .I1 (g19720), .I2 (g1345));
NR4X1 gate20194(.O (g10179), .I1 (g2098), .I2 (g1964), .I3 (g1830), .I4 (g1696));
NR4X1 gate20195(.O (g9664), .I1 (g4878), .I2 (g4871), .I3 (g4864), .I4 (g4836));
NR2X1 gate20196(.O (g15096), .I1 (g13191), .I2 (g12867));
NR2X1 gate20197(.O (g30146), .I1 (g28833), .I2 (g7411));
NR2X1 gate20198(.O (g25540), .I1 (g22409), .I2 (g22360));
NR2X1 gate20199(.O (g14178), .I1 (g8899), .I2 (g11083));
NR2X1 gate20200(.O (g31482), .I1 (g8883), .I2 (g29697));
NR2X1 gate20201(.O (g30290), .I1 (g6682), .I2 (g29110));
NR2X1 gate20202(.O (g28568), .I1 (g10323), .I2 (g27617));
NR2X1 gate20203(.O (g25203), .I1 (g6428), .I2 (g23756));
NR2X1 gate20204(.O (g11309), .I1 (g8587), .I2 (g8728));
NR3X1 gate20205(.O (g11571), .I1 (g10323), .I2 (g3512), .I3 (g3506));
NR2X1 gate20206(.O (g22523), .I1 (g1345), .I2 (g19720));
NR2X1 gate20207(.O (g14417), .I1 (g12149), .I2 (g9648));
NR2X1 gate20208(.O (g12622), .I1 (g9569), .I2 (g9518));
NR2X1 gate20209(.O (g26715), .I1 (g23711), .I2 (g25203));
NR2X1 gate20210(.O (g23763), .I1 (g2795), .I2 (g21276));
NR2X1 gate20211(.O (g14334), .I1 (g12044), .I2 (g9337));
NR2X1 gate20212(.O (g16232), .I1 (g13516), .I2 (g4950));
NR2X1 gate20213(.O (g11976), .I1 (g9595), .I2 (g7379));
NR2X1 gate20214(.O (g33090), .I1 (g31997), .I2 (g4593));
NR3X1 gate20215(.O (g31233), .I1 (g8522), .I2 (g29778), .I3 (g24825));
NR2X1 gate20216(.O (g17727), .I1 (g12486), .I2 (g12983));
NR2X1 gate20217(.O (g11954), .I1 (g9538), .I2 (g7314));
NR2X1 gate20218(.O (g13954), .I1 (g8663), .I2 (g11276));
NR2X1 gate20219(.O (g28510), .I1 (g3530), .I2 (g27617));
NR2X1 gate20220(.O (g12333), .I1 (g1624), .I2 (g8139));
NR2X1 gate20221(.O (g26297), .I1 (g8519), .I2 (g24825));
NR2X1 gate20222(.O (g15129), .I1 (g6984), .I2 (g13638));
NR2X1 gate20223(.O (g12852), .I1 (g6847), .I2 (g10430));
NR2X1 gate20224(.O (g15057), .I1 (g6810), .I2 (g13350));
NR2X1 gate20225(.O (g11669), .I1 (g3863), .I2 (g8026));
NR2X1 gate20226(.O (g15128), .I1 (g13638), .I2 (g12880));
NR2X1 gate20227(.O (g14000), .I1 (g8766), .I2 (g12259));
NR2X1 gate20228(.O (g33449), .I1 (g10311), .I2 (g31950));
NR2X1 gate20229(.O (g33448), .I1 (g7785), .I2 (g31950));
NR2X1 gate20230(.O (g14568), .I1 (g12000), .I2 (g9915));
NR2X1 gate20231(.O (g17175), .I1 (g1216), .I2 (g13545));
NR2X1 gate20232(.O (g10123), .I1 (g4294), .I2 (g4297));
NR2X1 gate20233(.O (g21655), .I1 (g17657), .I2 (g17700));
NR3X1 gate20234(.O (g34354), .I1 (g9003), .I2 (g34162), .I3 (g11083));
NR3X1 gate20235(.O (g12609), .I1 (g7766), .I2 (g5863), .I3 (g5857));
NR4X1 gate20236(.O (g14751), .I1 (g10622), .I2 (g10617), .I3 (g10609), .I4 (g10603));
NR2X1 gate20237(.O (g14772), .I1 (g6044), .I2 (g12252));
NR2X1 gate20238(.O (g8182), .I1 (g405), .I2 (g392));
NR2X1 gate20239(.O (g28493), .I1 (g3873), .I2 (g27635));
NR2X1 gate20240(.O (g26546), .I1 (g24858), .I2 (g24846));
NR2X1 gate20241(.O (g19981), .I1 (g3727), .I2 (g16316));
NR2X1 gate20242(.O (g28340), .I1 (g27439), .I2 (g26339));
NR2X1 gate20243(.O (g14416), .I1 (g12148), .I2 (g9541));
NR2X1 gate20244(.O (g11610), .I1 (g7980), .I2 (g3155));
NR2X1 gate20245(.O (g25784), .I1 (g25507), .I2 (g25485));
NR2X1 gate20246(.O (g27973), .I1 (g7187), .I2 (g25839));
NR2X1 gate20247(.O (g33148), .I1 (g4854), .I2 (g32072));
NR2X1 gate20248(.O (g25956), .I1 (g1413), .I2 (g24609));
NR2X1 gate20249(.O (g11255), .I1 (g8623), .I2 (g6928));
NR2X1 gate20250(.O (g33097), .I1 (g31950), .I2 (g4628));
NR2X1 gate20251(.O (g14391), .I1 (g12112), .I2 (g9585));
NR2X1 gate20252(.O (g12798), .I1 (g5535), .I2 (g9381));
NR3X1 gate20253(.O (g10510), .I1 (g7183), .I2 (g4593), .I3 (g4584));
NR2X1 gate20254(.O (g11270), .I1 (g8431), .I2 (g8434));
NR2X1 gate20255(.O (g16198), .I1 (g9247), .I2 (g13574));
NR2X1 gate20256(.O (g7352), .I1 (g1526), .I2 (g1514));
NR2X1 gate20257(.O (g26625), .I1 (g23560), .I2 (g25144));
NR2X1 gate20258(.O (g27732), .I1 (g9364), .I2 (g25791));
NR3X1 gate20259(.O (g13939), .I1 (g4899), .I2 (g8822), .I3 (g11173));
NR2X1 gate20260(.O (g32017), .I1 (g31504), .I2 (g23475));
NR2X1 gate20261(.O (g26296), .I1 (g8287), .I2 (g24732));
NR2X1 gate20262(.O (g26338), .I1 (g8458), .I2 (g24825));
NR2X1 gate20263(.O (g15056), .I1 (g6809), .I2 (g13350));
NR2X1 gate20264(.O (g27400), .I1 (g8553), .I2 (g26657));
NR2X1 gate20265(.O (g10615), .I1 (g1636), .I2 (g7308));
NR2X1 gate20266(.O (g31133), .I1 (g7953), .I2 (g29556));
NR2X1 gate20267(.O (g33133), .I1 (g32278), .I2 (g31503));
NR2X1 gate20268(.O (g28475), .I1 (g3863), .I2 (g27635));
NR2X1 gate20269(.O (g21143), .I1 (g15348), .I2 (g9517));
NR2X1 gate20270(.O (g19388), .I1 (g17181), .I2 (g14256));
NR2X1 gate20271(.O (g15145), .I1 (g12891), .I2 (g13716));
NR2X1 gate20272(.O (g24439), .I1 (g7400), .I2 (g22312));
NR2X1 gate20273(.O (g9700), .I1 (g2361), .I2 (g2287));
NR2X1 gate20274(.O (g11201), .I1 (g4125), .I2 (g7765));
NR2X1 gate20275(.O (g33112), .I1 (g31240), .I2 (g32194));
NR2X1 gate20276(.O (g27771), .I1 (g9809), .I2 (g25839));
NR2X1 gate20277(.O (g19140), .I1 (g7939), .I2 (g15695));
NR2X1 gate20278(.O (g19997), .I1 (g16231), .I2 (g13739));
NR2X1 gate20279(.O (g15132), .I1 (g12882), .I2 (g13638));
NR2X1 gate20280(.O (g12235), .I1 (g9234), .I2 (g9206));
NR2X1 gate20281(.O (g33096), .I1 (g31997), .I2 (g4608));
NR2X1 gate20282(.O (g14362), .I1 (g12080), .I2 (g9338));
NR2X1 gate20283(.O (g22537), .I1 (g19720), .I2 (g1367));
NR2X1 gate20284(.O (g15161), .I1 (g13809), .I2 (g7073));
NR2X1 gate20285(.O (g14165), .I1 (g8951), .I2 (g11083));
NR2X1 gate20286(.O (g29104), .I1 (g5188), .I2 (g27999));
NR2X1 gate20287(.O (g12515), .I1 (g9511), .I2 (g5873));
NR2X1 gate20288(.O (g15087), .I1 (g12860), .I2 (g13144));
NR2X1 gate20289(.O (g32424), .I1 (g8721), .I2 (g31294));
NR2X1 gate20290(.O (g34496), .I1 (g34370), .I2 (g27648));
NR2X1 gate20291(.O (g14437), .I1 (g9527), .I2 (g11178));
NR2X1 gate20292(.O (g11194), .I1 (g3288), .I2 (g6875));
NR2X1 gate20293(.O (g15069), .I1 (g6828), .I2 (g13416));
NR2X1 gate20294(.O (g14347), .I1 (g9309), .I2 (g11123));
NR3X1 gate20295(.O (g14253), .I1 (g10032), .I2 (g12259), .I3 (g9217));
NR2X1 gate20296(.O (g15068), .I1 (g6826), .I2 (g13416));
NR2X1 gate20297(.O (g17174), .I1 (g9194), .I2 (g14279));
NR2X1 gate20298(.O (g34067), .I1 (g33859), .I2 (g11772));
NR2X1 gate20299(.O (g11119), .I1 (g9180), .I2 (g9203));
NR2X1 gate20300(.O (g30150), .I1 (g28846), .I2 (g7424));
NR2X1 gate20301(.O (g33129), .I1 (g8630), .I2 (g32072));
NR2X1 gate20302(.O (g10821), .I1 (g7503), .I2 (g1384));
NR4X1 gate20303(.O (g12435), .I1 (g9012), .I2 (g8956), .I3 (g8904), .I4 (g8863));
NR2X1 gate20304(.O (g33128), .I1 (g4653), .I2 (g32057));
NR2X1 gate20305(.O (g14821), .I1 (g6390), .I2 (g12314));
NR2X1 gate20306(.O (g22522), .I1 (g19699), .I2 (g1024));
NR2X1 gate20307(.O (g11313), .I1 (g8669), .I2 (g3759));
NR2X1 gate20308(.O (g27345), .I1 (g9360), .I2 (g26636));
NR2X1 gate20309(.O (g12744), .I1 (g9402), .I2 (g6203));
NR2X1 gate20310(.O (g14516), .I1 (g12227), .I2 (g9704));
NR2X1 gate20311(.O (g11276), .I1 (g8534), .I2 (g8691));
NR2X1 gate20312(.O (g12849), .I1 (g6840), .I2 (g10430));
NR2X1 gate20313(.O (g17663), .I1 (g10205), .I2 (g12983));
NR2X1 gate20314(.O (g12848), .I1 (g6839), .I2 (g10430));
NR2X1 gate20315(.O (g27652), .I1 (g3355), .I2 (g26636));
NR2X1 gate20316(.O (g26256), .I1 (g23873), .I2 (g25479));
NR2X1 gate20317(.O (g22536), .I1 (g1379), .I2 (g19720));
NR2X1 gate20318(.O (g15086), .I1 (g13144), .I2 (g12859));
NR2X1 gate20319(.O (g12361), .I1 (g6455), .I2 (g10172));
NR2X1 gate20320(.O (g14726), .I1 (g10090), .I2 (g12166));
NR2X1 gate20321(.O (g30280), .I1 (g7064), .I2 (g29036));
NR3X1 gate20322(.O (g32455), .I1 (g31566), .I2 (I29985), .I3 (I29986));
NR2X1 gate20323(.O (g15159), .I1 (g13809), .I2 (g12902));
NR2X1 gate20324(.O (g16288), .I1 (g13794), .I2 (g417));
NR2X1 gate20325(.O (g14320), .I1 (g9257), .I2 (g11111));
NR2X1 gate20326(.O (g15158), .I1 (g13782), .I2 (g12901));
NR2X1 gate20327(.O (g30157), .I1 (g28833), .I2 (g7369));
NR2X1 gate20328(.O (g14122), .I1 (g8895), .I2 (g12259));
NR2X1 gate20329(.O (g15144), .I1 (g13716), .I2 (g12890));
NR2X1 gate20330(.O (g31498), .I1 (g9030), .I2 (g29540));
NR3X1 gate20331(.O (g28492), .I1 (g3857), .I2 (g7121), .I3 (g27635));
NR3X1 gate20332(.O (g8086), .I1 (g168), .I2 (g174), .I3 (g182));
NR2X1 gate20333(.O (g11907), .I1 (g7170), .I2 (g7184));
NR2X1 gate20334(.O (g33432), .I1 (g31997), .I2 (g6978));
NR2X1 gate20335(.O (g26314), .I1 (g24808), .I2 (g24802));
NR2X1 gate20336(.O (g12371), .I1 (g1760), .I2 (g8195));
NR2X1 gate20337(.O (g23835), .I1 (g2791), .I2 (g21303));
NR2X1 gate20338(.O (g11238), .I1 (g8584), .I2 (g6905));
NR2X1 gate20339(.O (g17213), .I1 (g11107), .I2 (g13501));
NR2X1 gate20340(.O (g12234), .I1 (g9776), .I2 (g9778));
NR2X1 gate20341(.O (g23586), .I1 (g17284), .I2 (g20717));
NR2X1 gate20342(.O (g33145), .I1 (g8677), .I2 (g32072));
NR2X1 gate20343(.O (g14164), .I1 (g9000), .I2 (g12259));
NR3X1 gate20344(.O (g11185), .I1 (g8038), .I2 (g8183), .I3 (g6804));
NR2X1 gate20345(.O (g13518), .I1 (g3719), .I2 (g11903));
NR2X1 gate20346(.O (g16488), .I1 (g13697), .I2 (g13656));
NR2X1 gate20347(.O (g16424), .I1 (g8064), .I2 (g13628));
NR2X1 gate20348(.O (g26268), .I1 (g283), .I2 (g24825));
NR2X1 gate20349(.O (g14575), .I1 (g10050), .I2 (g12749));
NR2X1 gate20350(.O (g11935), .I1 (g9485), .I2 (g7267));
NR3X1 gate20351(.O (g8131), .I1 (g4776), .I2 (g4801), .I3 (g4793));
NR2X1 gate20352(.O (g27012), .I1 (g6398), .I2 (g25856));
NR3X1 gate20353(.O (g13883), .I1 (g4709), .I2 (g4785), .I3 (g11155));
NR2X1 gate20354(.O (g33132), .I1 (g4843), .I2 (g32072));
NR2X1 gate20355(.O (g12163), .I1 (g5073), .I2 (g9989));
NR2X1 gate20356(.O (g28483), .I1 (g8080), .I2 (g27635));
NR2X1 gate20357(.O (g26993), .I1 (g5360), .I2 (g25805));
NR2X1 gate20358(.O (g33161), .I1 (g32090), .I2 (g7806));
NR2X1 gate20359(.O (g26667), .I1 (g23642), .I2 (g25175));
NR2X1 gate20360(.O (g30156), .I1 (g28789), .I2 (g14587));
NR2X1 gate20361(.O (g11729), .I1 (g3179), .I2 (g8059));
NR2X1 gate20362(.O (g13501), .I1 (g3368), .I2 (g11881));
NR2X1 gate20363(.O (g27829), .I1 (g7345), .I2 (g25856));
NR2X1 gate20364(.O (g14091), .I1 (g8854), .I2 (g12259));
NR2X1 gate20365(.O (g27828), .I1 (g9892), .I2 (g25856));
NR3X1 gate20366(.O (g22405), .I1 (g18957), .I2 (g20136), .I3 (g20114));
NR2X1 gate20367(.O (g15669), .I1 (g11945), .I2 (g14272));
NR2X1 gate20368(.O (g12358), .I1 (g10019), .I2 (g10022));
NR2X1 gate20369(.O (g27344), .I1 (g8390), .I2 (g26636));
NR2X1 gate20370(.O (g12121), .I1 (g10117), .I2 (g9762));
NR2X1 gate20371(.O (g21193), .I1 (g15348), .I2 (g12135));
NR2X1 gate20372(.O (g22929), .I1 (g19773), .I2 (g12970));
NR2X1 gate20373(.O (g31068), .I1 (g4801), .I2 (g29540));
NR2X1 gate20374(.O (g11566), .I1 (g3161), .I2 (g7964));
NR2X1 gate20375(.O (g13622), .I1 (g278), .I2 (g11166));
NR2X1 gate20376(.O (g31970), .I1 (g9024), .I2 (g30583));
NR2X1 gate20377(.O (g12173), .I1 (g10050), .I2 (g7074));
NR2X1 gate20378(.O (g28509), .I1 (g8107), .I2 (g27602));
NR2X1 gate20379(.O (g16219), .I1 (g13498), .I2 (g4760));
NR2X1 gate20380(.O (g14522), .I1 (g9924), .I2 (g12656));
NR2X1 gate20381(.O (g11653), .I1 (g7980), .I2 (g7964));
NR2X1 gate20382(.O (g22357), .I1 (g1024), .I2 (g19699));
NR3X1 gate20383(.O (g29145), .I1 (g6549), .I2 (g7812), .I3 (g26994));
NR2X1 gate20384(.O (g12029), .I1 (g5644), .I2 (g7028));
NR2X1 gate20385(.O (g10862), .I1 (g7701), .I2 (g7840));
NR2X1 gate20386(.O (g11415), .I1 (g8080), .I2 (g8026));
NR2X1 gate20387(.O (g29198), .I1 (g7766), .I2 (g28020));
NR2X1 gate20388(.O (g13852), .I1 (g11320), .I2 (g8347));
NR2X1 gate20389(.O (g30601), .I1 (g16279), .I2 (g29718));
NR2X1 gate20390(.O (g28452), .I1 (g3161), .I2 (g27602));
NR2X1 gate20391(.O (g27927), .I1 (g9621), .I2 (g25856));
NR2X1 gate20392(.O (g16201), .I1 (g13462), .I2 (g4704));
NR2X1 gate20393(.O (g15093), .I1 (g13177), .I2 (g6904));
NR2X1 gate20394(.O (g30143), .I1 (g28761), .I2 (g14566));
NR2X1 gate20395(.O (g23063), .I1 (g16313), .I2 (g19887));
NR2X1 gate20396(.O (g15065), .I1 (g13394), .I2 (g12840));
NR2X1 gate20397(.O (g30169), .I1 (g28833), .I2 (g14613));
NR2X1 gate20398(.O (g14397), .I1 (g12120), .I2 (g9416));
NR2X1 gate20399(.O (g12604), .I1 (g5517), .I2 (g9239));
NR2X1 gate20400(.O (g27770), .I1 (g9386), .I2 (g25821));
NR2X1 gate20401(.O (g19338), .I1 (g16031), .I2 (g1306));
NR2X1 gate20402(.O (g12755), .I1 (g6555), .I2 (g9407));
NR2X1 gate20403(.O (g33125), .I1 (g8606), .I2 (g32057));
NR2X1 gate20404(.O (g21209), .I1 (g15483), .I2 (g9575));
NR2X1 gate20405(.O (g14872), .I1 (g6736), .I2 (g12364));
NR2X1 gate20406(.O (g19968), .I1 (g17062), .I2 (g11223));
NR2X1 gate20407(.O (g23208), .I1 (g20035), .I2 (g16324));
NR2X1 gate20408(.O (g15160), .I1 (g12903), .I2 (g13809));
NR2X1 gate20409(.O (g13799), .I1 (g8584), .I2 (g11663));
NR2X1 gate20410(.O (g17482), .I1 (g9523), .I2 (g14434));
NR2X1 gate20411(.O (g33144), .I1 (g4664), .I2 (g32057));
NR3X1 gate20412(.O (g33823), .I1 (g8774), .I2 (g33306), .I3 (g11083));
NR2X1 gate20413(.O (g20234), .I1 (g17140), .I2 (g14207));
NR2X1 gate20414(.O (g29069), .I1 (g9381), .I2 (g28010));
NR2X1 gate20415(.O (g11184), .I1 (g513), .I2 (g9040));
NR2X1 gate20416(.O (g7158), .I1 (g5752), .I2 (g5712));
NR4X1 gate20417(.O (g10205), .I1 (g2657), .I2 (g2523), .I3 (g2389), .I4 (g2255));
NR2X1 gate20418(.O (g24514), .I1 (g23619), .I2 (g23657));
NR2X1 gate20419(.O (g30922), .I1 (g16662), .I2 (g29810));
NR2X1 gate20420(.O (g29886), .I1 (g3288), .I2 (g28458));
NR2X1 gate20421(.O (g11692), .I1 (g8021), .I2 (g7985));
NR2X1 gate20422(.O (g16313), .I1 (g8005), .I2 (g13600));
NR2X1 gate20423(.O (g27926), .I1 (g9467), .I2 (g25856));
NR2X1 gate20424(.O (g13013), .I1 (g7957), .I2 (g10762));
NR2X1 gate20425(.O (g19070), .I1 (g16957), .I2 (g11720));
NR2X1 gate20426(.O (g22513), .I1 (g1002), .I2 (g19699));
NR2X1 gate20427(.O (g15155), .I1 (g12899), .I2 (g13782));
NR2X1 gate20428(.O (g11207), .I1 (g3639), .I2 (g6905));
NR2X1 gate20429(.O (g15170), .I1 (g7118), .I2 (g14279));
NR2X1 gate20430(.O (g22448), .I1 (g1018), .I2 (g19699));
NR2X1 gate20431(.O (g13539), .I1 (g8594), .I2 (g12735));
NR2X1 gate20432(.O (g13005), .I1 (g7939), .I2 (g10762));
NR2X1 gate20433(.O (g25321), .I1 (g23835), .I2 (g14645));
NR2X1 gate20434(.O (g14396), .I1 (g12119), .I2 (g9489));
NR2X1 gate20435(.O (g14731), .I1 (g5698), .I2 (g12204));
NR2X1 gate20436(.O (g15167), .I1 (g13835), .I2 (g12908));
NR2X1 gate20437(.O (g14413), .I1 (g11914), .I2 (g9638));
NR2X1 gate20438(.O (g28803), .I1 (g27730), .I2 (g22763));
NR2X1 gate20439(.O (g11771), .I1 (g8921), .I2 (g4185));
NR2X1 gate20440(.O (g25800), .I1 (g25518), .I2 (g25510));
NR2X1 gate20441(.O (g27766), .I1 (g9716), .I2 (g25791));
NR2X1 gate20442(.O (g23711), .I1 (g9892), .I2 (g21253));
NR2X1 gate20443(.O (g30117), .I1 (g28739), .I2 (g7252));
NR2X1 gate20444(.O (g29144), .I1 (g9518), .I2 (g26977));
NR2X1 gate20445(.O (g19402), .I1 (g15979), .I2 (g13133));
NR2X1 gate20446(.O (g23108), .I1 (g16424), .I2 (g19932));
NR2X1 gate20447(.O (g17148), .I1 (g827), .I2 (g14279));
NR2X1 gate20448(.O (g11414), .I1 (g8591), .I2 (g8593));
NR2X1 gate20449(.O (g16476), .I1 (g8119), .I2 (g13667));
NR3X1 gate20450(.O (g32585), .I1 (g31542), .I2 (I30123), .I3 (I30124));
NR2X1 gate20451(.O (g15053), .I1 (g12836), .I2 (g13350));
NR2X1 gate20452(.O (g28482), .I1 (g3522), .I2 (g27617));
NR2X1 gate20453(.O (g30123), .I1 (g28768), .I2 (g7328));
NR3X1 gate20454(.O (g27629), .I1 (g8891), .I2 (g26382), .I3 (g12259));
NR2X1 gate20455(.O (g28552), .I1 (g10295), .I2 (g27602));
NR2X1 gate20456(.O (g15101), .I1 (g12871), .I2 (g14591));
NR2X1 gate20457(.O (g12246), .I1 (g9880), .I2 (g9883));
NR2X1 gate20458(.O (g11584), .I1 (g8229), .I2 (g8172));
NR2X1 gate20459(.O (g30265), .I1 (g7051), .I2 (g29036));
NR2X1 gate20460(.O (g14640), .I1 (g12371), .I2 (g9824));
NR2X1 gate20461(.O (g15064), .I1 (g6820), .I2 (g13394));
NR2X1 gate20462(.O (g10803), .I1 (g1384), .I2 (g7503));
NR2X1 gate20463(.O (g12591), .I1 (g504), .I2 (g9040));
NR2X1 gate20464(.O (g12785), .I1 (g9472), .I2 (g6549));
NR2X1 gate20465(.O (g27355), .I1 (g8443), .I2 (g26657));
NR2X1 gate20466(.O (g13114), .I1 (g7528), .I2 (g10741));
NR2X1 gate20467(.O (g27825), .I1 (g9316), .I2 (g25821));
NR2X1 gate20468(.O (g11435), .I1 (g8107), .I2 (g3171));
NR2X1 gate20469(.O (g11107), .I1 (g9095), .I2 (g9177));
NR2X1 gate20470(.O (g15166), .I1 (g13835), .I2 (g7096));
NR2X1 gate20471(.O (g12858), .I1 (g10365), .I2 (g10430));
NR2X1 gate20472(.O (g11345), .I1 (g8477), .I2 (g8479));
NR2X1 gate20473(.O (g33093), .I1 (g31997), .I2 (g4601));
NR2X1 gate20474(.O (g31294), .I1 (g11326), .I2 (g29660));
NR2X1 gate20475(.O (g11940), .I1 (g2712), .I2 (g10084));
NR2X1 gate20476(.O (g27367), .I1 (g8155), .I2 (g26636));
NR2X1 gate20477(.O (g14027), .I1 (g8734), .I2 (g11363));
NR2X1 gate20478(.O (g11804), .I1 (g8938), .I2 (g4975));
NR2X1 gate20479(.O (g15570), .I1 (g822), .I2 (g14279));
NR2X1 gate20480(.O (g14248), .I1 (g6065), .I2 (g10578));
NR2X1 gate20481(.O (g16215), .I1 (g1211), .I2 (g13545));
NR2X1 gate20482(.O (g24990), .I1 (g8898), .I2 (g23324));
NR2X1 gate20483(.O (g14003), .I1 (g9003), .I2 (g11083));
NR2X1 gate20484(.O (g15074), .I1 (g12845), .I2 (g13416));
NR2X1 gate20485(.O (g12318), .I1 (g10172), .I2 (g6451));
NR2X1 gate20486(.O (g27059), .I1 (g7577), .I2 (g25895));
NR3X1 gate20487(.O (g15594), .I1 (g10614), .I2 (g13026), .I3 (g7285));
NR2X1 gate20488(.O (g12059), .I1 (g9853), .I2 (g7004));
NR2X1 gate20489(.O (g12025), .I1 (g9705), .I2 (g7461));
NR2X1 gate20490(.O (g33160), .I1 (g8672), .I2 (g32057));
NR2X1 gate20491(.O (g12540), .I1 (g2587), .I2 (g8381));
NR2X1 gate20492(.O (g13500), .I1 (g8480), .I2 (g12641));
NR2X1 gate20493(.O (g15092), .I1 (g12864), .I2 (g13177));
NR2X1 gate20494(.O (g28149), .I1 (g27598), .I2 (g27612));
NR2X1 gate20495(.O (g15154), .I1 (g13782), .I2 (g12898));
NR2X1 gate20496(.O (g21062), .I1 (g9547), .I2 (g17297));
NR2X1 gate20497(.O (g14090), .I1 (g8851), .I2 (g12259));
NR2X1 gate20498(.O (g13004), .I1 (g7933), .I2 (g10741));
NR2X1 gate20499(.O (g33075), .I1 (g31997), .I2 (g7163));
NR2X1 gate20500(.O (g19268), .I1 (g15979), .I2 (g962));
NR3X1 gate20501(.O (g12377), .I1 (g6856), .I2 (g2748), .I3 (g9708));
NR2X1 gate20502(.O (g12739), .I1 (g9321), .I2 (g9274));
NR2X1 gate20503(.O (g30130), .I1 (g28761), .I2 (g7275));
NR3X1 gate20504(.O (g24701), .I1 (g979), .I2 (g23024), .I3 (g19778));
NR2X1 gate20505(.O (g12146), .I1 (g1783), .I2 (g8241));
NR2X1 gate20506(.O (g12645), .I1 (g4467), .I2 (g6961));
NR2X1 gate20507(.O (g13947), .I1 (g8948), .I2 (g11083));
NR2X1 gate20508(.O (g11273), .I1 (g3061), .I2 (g8620));
NR2X1 gate20509(.O (g14513), .I1 (g12222), .I2 (g9754));
NR3X1 gate20510(.O (g29705), .I1 (g28399), .I2 (g8284), .I3 (g8404));
NR2X1 gate20511(.O (g14449), .I1 (g12194), .I2 (g9653));
NR3X1 gate20512(.O (g29189), .I1 (g9462), .I2 (g26977), .I3 (g7791));
NR2X1 gate20513(.O (g33419), .I1 (g31978), .I2 (g7627));
NR2X1 gate20514(.O (g14448), .I1 (g12192), .I2 (g9699));
NR2X1 gate20515(.O (g11972), .I1 (g9591), .I2 (g7361));
NR2X1 gate20516(.O (g27366), .I1 (g8016), .I2 (g26636));
NR2X1 gate20517(.O (g7567), .I1 (g979), .I2 (g990));
NR2X1 gate20518(.O (g14212), .I1 (g5373), .I2 (g10537));
NR2X1 gate20519(.O (g12632), .I1 (g9631), .I2 (g6565));
NR2X1 gate20520(.O (g24766), .I1 (g3385), .I2 (g23132));
NR2X1 gate20521(.O (g23051), .I1 (g7960), .I2 (g19427));
NR3X1 gate20522(.O (g34703), .I1 (g8899), .I2 (g34545), .I3 (g11083));
NR3X1 gate20523(.O (g11514), .I1 (g10295), .I2 (g3161), .I3 (g3155));
NR2X1 gate20524(.O (g12226), .I1 (g2476), .I2 (g8373));
NR2X1 gate20525(.O (g31119), .I1 (g7898), .I2 (g29556));
NR2X1 gate20526(.O (g26873), .I1 (g25374), .I2 (g25331));
NR2X1 gate20527(.O (g11012), .I1 (g7693), .I2 (g7846));
NR2X1 gate20528(.O (g15139), .I1 (g12886), .I2 (g13680));
NR2X1 gate20529(.O (g26209), .I1 (g23124), .I2 (g24779));
NR2X1 gate20530(.O (g15138), .I1 (g13680), .I2 (g6993));
NR2X1 gate20531(.O (g11473), .I1 (g8107), .I2 (g8059));
NR2X1 gate20532(.O (g29915), .I1 (g6941), .I2 (g28484));
NR2X1 gate20533(.O (g27354), .I1 (g8064), .I2 (g26636));
NR2X1 gate20534(.O (g12297), .I1 (g9269), .I2 (g9239));
NR2X1 gate20535(.O (g13325), .I1 (g7841), .I2 (g10741));
NR2X1 gate20536(.O (g12980), .I1 (g7909), .I2 (g10741));
NR2X1 gate20537(.O (g12824), .I1 (g5881), .I2 (g9451));
NR2X1 gate20538(.O (g25952), .I1 (g1542), .I2 (g24609));
NR2X1 gate20539(.O (g13946), .I1 (g8651), .I2 (g11083));
NR2X1 gate20540(.O (g25175), .I1 (g5736), .I2 (g23692));
NR2X1 gate20541(.O (g14228), .I1 (g5719), .I2 (g10561));
NR2X1 gate20542(.O (g15585), .I1 (g11862), .I2 (g14194));
NR2X1 gate20543(.O (g26346), .I1 (g8522), .I2 (g24825));
NR2X1 gate20544(.O (g15608), .I1 (g11885), .I2 (g14212));
NR2X1 gate20545(.O (g15052), .I1 (g12835), .I2 (g13350));
NR2X1 gate20546(.O (g12211), .I1 (g10099), .I2 (g7097));
NR2X1 gate20547(.O (g31008), .I1 (g30004), .I2 (g30026));
NR2X1 gate20548(.O (g31476), .I1 (g4709), .I2 (g29697));
NR2X1 gate20549(.O (g29167), .I1 (g9576), .I2 (g26994));
NR2X1 gate20550(.O (g17198), .I1 (g9282), .I2 (g14279));
NR2X1 gate20551(.O (g27659), .I1 (g3706), .I2 (g26657));
NR2X1 gate20552(.O (g17393), .I1 (g9386), .I2 (g14379));
NR2X1 gate20553(.O (g12700), .I1 (g9321), .I2 (g5857));
NR2X1 gate20554(.O (g12659), .I1 (g9451), .I2 (g9392));
NR2X1 gate20555(.O (g12126), .I1 (g9989), .I2 (g5069));
NR2X1 gate20556(.O (g30136), .I1 (g28799), .I2 (g7380));
NR2X1 gate20557(.O (g19953), .I1 (g16220), .I2 (g13712));
NR2X1 gate20558(.O (g10793), .I1 (g1389), .I2 (g7503));
NR2X1 gate20559(.O (g14793), .I1 (g2988), .I2 (g12228));
NR2X1 gate20560(.O (g27338), .I1 (g9291), .I2 (g26616));
NR2X1 gate20561(.O (g12296), .I1 (g9860), .I2 (g9862));
NR2X1 gate20562(.O (g9762), .I1 (g2495), .I2 (g2421));
NR2X1 gate20563(.O (g23662), .I1 (g17393), .I2 (g20995));
NR2X1 gate20564(.O (g27969), .I1 (g7170), .I2 (g25821));
NR2X1 gate20565(.O (g14549), .I1 (g9992), .I2 (g12705));
NR2X1 gate20566(.O (g11755), .I1 (g4709), .I2 (g8796));
NR2X1 gate20567(.O (g29900), .I1 (g3639), .I2 (g28471));
NR2X1 gate20568(.O (g33092), .I1 (g31978), .I2 (g4332));
NR2X1 gate20569(.O (g11563), .I1 (g8059), .I2 (g8011));
NR2X1 gate20570(.O (g12855), .I1 (g10430), .I2 (g6854));
NR2X1 gate20571(.O (g31935), .I1 (g30583), .I2 (g4349));
NR3X1 gate20572(.O (g23204), .I1 (g10685), .I2 (g19462), .I3 (g16488));
NR2X1 gate20573(.O (g14002), .I1 (g8681), .I2 (g11083));
NR2X1 gate20574(.O (g17657), .I1 (g14751), .I2 (g12955));
NR3X1 gate20575(.O (g11191), .I1 (g4776), .I2 (g4801), .I3 (g9030));
NR2X1 gate20576(.O (g28498), .I1 (g8172), .I2 (g27635));
NR2X1 gate20577(.O (g15100), .I1 (g13191), .I2 (g12870));
NR2X1 gate20578(.O (g12581), .I1 (g9569), .I2 (g6219));
NR2X1 gate20579(.O (g33439), .I1 (g31950), .I2 (g4633));
NR2X1 gate20580(.O (g7175), .I1 (g6098), .I2 (g6058));
NR2X1 gate20581(.O (g33438), .I1 (g31950), .I2 (g4621));
NR2X1 gate20582(.O (g7139), .I1 (g5406), .I2 (g5366));
NR2X1 gate20583(.O (g22545), .I1 (g1373), .I2 (g19720));
NR3X1 gate20584(.O (g28031), .I1 (g21209), .I2 (I26522), .I3 (I26523));
NR2X1 gate20585(.O (g12067), .I1 (g5990), .I2 (g7051));
NR2X1 gate20586(.O (g14512), .I1 (g11955), .I2 (g9753));
NR2X1 gate20587(.O (g27735), .I1 (g7262), .I2 (g25821));
NR2X1 gate20588(.O (g27877), .I1 (g9397), .I2 (g25839));
NR3X1 gate20589(.O (g28529), .I1 (g8070), .I2 (g27617), .I3 (g10323));
NR2X1 gate20590(.O (g12150), .I1 (g2208), .I2 (g8259));
NR2X1 gate20591(.O (g33139), .I1 (g8650), .I2 (g32057));
NR2X1 gate20592(.O (g10831), .I1 (g7690), .I2 (g7827));
NR2X1 gate20593(.O (g13032), .I1 (g7577), .I2 (g10762));
NR2X1 gate20594(.O (g33138), .I1 (g32287), .I2 (g31514));
NR2X1 gate20595(.O (g14445), .I1 (g12188), .I2 (g9693));
NR2X1 gate20596(.O (g12695), .I1 (g9269), .I2 (g9239));
NR3X1 gate20597(.O (g29675), .I1 (g28380), .I2 (g8236), .I3 (g8354));
NR2X1 gate20598(.O (g26183), .I1 (g23079), .I2 (g24766));
NR2X1 gate20599(.O (g30252), .I1 (g7028), .I2 (g29008));
NR2X1 gate20600(.O (g7304), .I1 (g1183), .I2 (g1171));
NR2X1 gate20601(.O (g14611), .I1 (g12333), .I2 (g9749));
NR2X1 gate20602(.O (g7499), .I1 (g333), .I2 (g355));
NR3X1 gate20603(.O (g14988), .I1 (g10816), .I2 (g10812), .I3 (g10805));
NR2X1 gate20604(.O (g11360), .I1 (g3763), .I2 (g8669));
NR2X1 gate20605(.O (g26872), .I1 (g25411), .I2 (g25371));
NR2X1 gate20606(.O (g14271), .I1 (g10002), .I2 (g10874));
NR2X1 gate20607(.O (g30183), .I1 (g28880), .I2 (g14644));
NR2X1 gate20608(.O (g19430), .I1 (g17150), .I2 (g14220));
NR2X1 gate20609(.O (g15141), .I1 (g12888), .I2 (g13680));
NR2X1 gate20610(.O (g14145), .I1 (g8945), .I2 (g12259));
NR2X1 gate20611(.O (g12256), .I1 (g10136), .I2 (g6105));
NR2X1 gate20612(.O (g25948), .I1 (g7752), .I2 (g24609));
NR2X1 gate20613(.O (g24497), .I1 (g23533), .I2 (g23553));
NR2X1 gate20614(.O (g14529), .I1 (g6336), .I2 (g12749));
NR2X1 gate20615(.O (g27102), .I1 (g26750), .I2 (g26779));
NR2X1 gate20616(.O (g15135), .I1 (g6990), .I2 (g13638));
NR2X1 gate20617(.O (g26574), .I1 (g24887), .I2 (g24861));
NR2X1 gate20618(.O (g14393), .I1 (g12115), .I2 (g9488));
NR2X1 gate20619(.O (g14365), .I1 (g12084), .I2 (g9339));
NR3X1 gate20620(.O (g32845), .I1 (g30673), .I2 (I30399), .I3 (I30400));
NR2X1 gate20621(.O (g17309), .I1 (g9305), .I2 (g14344));
NR2X1 gate20622(.O (g15049), .I1 (g13350), .I2 (g6799));
NR2X1 gate20623(.O (g11950), .I1 (g9220), .I2 (g9166));
NR2X1 gate20624(.O (g10709), .I1 (g7499), .I2 (g351));
NR3X1 gate20625(.O (g27511), .I1 (g22137), .I2 (g26866), .I3 (g20277));
NR2X1 gate20626(.O (g12854), .I1 (g6849), .I2 (g10430));
NR2X1 gate20627(.O (g28425), .I1 (g27493), .I2 (g26351));
NR4X1 gate20628(.O (g34912), .I1 (g34883), .I2 (g20277), .I3 (g20242), .I4 (g21370));
NR3X1 gate20629(.O (g25851), .I1 (g4311), .I2 (g24380), .I3 (g24369));
NR3X1 gate20630(.O (g13996), .I1 (g8938), .I2 (g8822), .I3 (g11173));
NR3X1 gate20631(.O (g28444), .I1 (g8575), .I2 (g27463), .I3 (g24825));
NR2X1 gate20632(.O (g15106), .I1 (g12872), .I2 (g10430));
NR2X1 gate20633(.O (g17954), .I1 (g832), .I2 (g14279));
NR2X1 gate20634(.O (g12550), .I1 (g9300), .I2 (g9259));
NR2X1 gate20635(.O (g12314), .I1 (g10053), .I2 (g10207));
NR2X1 gate20636(.O (g14602), .I1 (g10099), .I2 (g12790));
NR2X1 gate20637(.O (g27721), .I1 (g9672), .I2 (g25805));
NR2X1 gate20638(.O (g12085), .I1 (g10082), .I2 (g9700));
NR2X1 gate20639(.O (g22488), .I1 (g19699), .I2 (g1002));
NR2X1 gate20640(.O (g14337), .I1 (g12049), .I2 (g9284));
NR3X1 gate20641(.O (g11203), .I1 (g4966), .I2 (g4991), .I3 (g9064));
NR2X1 gate20642(.O (g13044), .I1 (g7349), .I2 (g10762));
NR4X1 gate20643(.O (g14792), .I1 (g10653), .I2 (g10623), .I3 (g10618), .I4 (g10611));
NR3X1 gate20644(.O (g28353), .I1 (g9073), .I2 (g27654), .I3 (g24732));
NR2X1 gate20645(.O (g29200), .I1 (g7791), .I2 (g26977));
NR2X1 gate20646(.O (g9640), .I1 (g1802), .I2 (g1728));
NR2X1 gate20647(.O (g19063), .I1 (g7909), .I2 (g15674));
NR2X1 gate20648(.O (g33100), .I1 (g32172), .I2 (g31188));
NR2X1 gate20649(.O (g13377), .I1 (g7873), .I2 (g10762));
NR2X1 gate20650(.O (g14425), .I1 (g5644), .I2 (g12656));
NR2X1 gate20651(.O (g27734), .I1 (g9733), .I2 (g25821));
NR2X1 gate20652(.O (g15163), .I1 (g13809), .I2 (g12905));
NR2X1 gate20653(.O (g30929), .I1 (g29803), .I2 (g29835));
NR2X1 gate20654(.O (g19873), .I1 (g15755), .I2 (g1395));
NR3X1 gate20655(.O (g10918), .I1 (g1532), .I2 (g7751), .I3 (g7778));
NR2X1 gate20656(.O (g19422), .I1 (g16031), .I2 (g13141));
NR2X1 gate20657(.O (g14444), .I1 (g11936), .I2 (g9692));
NR3X1 gate20658(.O (g12667), .I1 (g7791), .I2 (g6209), .I3 (g6203));
NR3X1 gate20659(.O (g19209), .I1 (g12971), .I2 (g15614), .I3 (g11320));
NR3X1 gate20660(.O (g13698), .I1 (g528), .I2 (g12527), .I3 (g11185));
NR2X1 gate20661(.O (g31515), .I1 (g4983), .I2 (g29556));
NR2X1 gate20662(.O (g29184), .I1 (g9631), .I2 (g26994));
NR2X1 gate20663(.O (g23626), .I1 (g17309), .I2 (g20854));
NR2X1 gate20664(.O (g15724), .I1 (g13858), .I2 (g11374));
NR2X1 gate20665(.O (g24018), .I1 (I23162), .I2 (I23163));
NR2X1 gate20666(.O (g30282), .I1 (g6336), .I2 (g29073));
NR2X1 gate20667(.O (g19453), .I1 (g17199), .I2 (g14316));
NR2X1 gate20668(.O (g15121), .I1 (g12874), .I2 (g13605));
NR2X1 gate20669(.O (g12443), .I1 (g9374), .I2 (g9300));
NR2X1 gate20670(.O (g19436), .I1 (g17176), .I2 (g14233));
NR2X1 gate20671(.O (g13661), .I1 (g528), .I2 (g11185));
NR2X1 gate20672(.O (g11715), .I1 (g8080), .I2 (g8026));
NR3X1 gate20673(.O (g29005), .I1 (g5164), .I2 (g7704), .I3 (g27999));
NR2X1 gate20674(.O (g33107), .I1 (g32180), .I2 (g31223));
NR2X1 gate20675(.O (g12601), .I1 (g9381), .I2 (g9311));
NR2X1 gate20676(.O (g15134), .I1 (g13638), .I2 (g12884));
NR2X1 gate20677(.O (g14364), .I1 (g12083), .I2 (g9415));
NR2X1 gate20678(.O (g25769), .I1 (g25453), .I2 (g25414));
NR2X1 gate20679(.O (g11385), .I1 (g8021), .I2 (g7985));
endmodule