module s5378_0(clk, n3065gat, n3066gat, n3067gat, n3068gat, n3069gat, n3070gat, n3071gat, n3072gat, n3073gat, n3074gat, n3075gat, n3076gat, n3077gat, n3078gat, n3079gat, n3080gat, n3081gat, n3082gat, n3083gat, n3084gat, n3085gat, n3086gat, n3087gat, n3088gat, n3089gat, n3090gat, n3091gat, n3092gat, n3093gat, n3094gat, n3095gat, n3097gat, n3098gat, n3099gat, n3100gat, n3104gat, n3105gat, n3106gat, n3107gat, n3108gat, n3109gat, n3110gat, n3111gat, n3112gat, n3113gat, n3114gat, n3115gat, n3116gat, n3117gat, n3118gat, n3119gat, n3120gat, n3121gat, n3122gat, n3123gat, n3124gat, n3125gat, n3126gat, n3127gat, n3128gat, n3129gat, n3130gat, n3131gat, n3132gat, n3133gat, n3134gat, n3135gat, n3136gat, n3137gat, n3138gat, n3139gat, n3140gat, n3141gat, n3142gat, n3143gat, n3144gat, n3145gat, n3146gat, n3147gat, n3148gat, n3149gat, n3150gat, n3151gat, n3152gat);
input clk, n3065gat, n3066gat, n3067gat, n3068gat, n3069gat, n3070gat, n3071gat, n3072gat, n3073gat, n3074gat, n3075gat, n3076gat, n3077gat, n3078gat, n3079gat, n3080gat, n3081gat, n3082gat, n3083gat, n3084gat, n3085gat, n3086gat, n3087gat, n3088gat, n3089gat, n3090gat, n3091gat, n3092gat, n3093gat, n3094gat, n3095gat, n3097gat, n3098gat, n3099gat, n3100gat;
output n3104gat, n3105gat, n3106gat, n3107gat, n3108gat, n3109gat, n3110gat, n3111gat, n3112gat, n3113gat, n3114gat, n3115gat, n3116gat, n3117gat, n3118gat, n3119gat, n3120gat, n3121gat, n3122gat, n3123gat, n3124gat, n3125gat, n3126gat, n3127gat, n3128gat, n3129gat, n3130gat, n3131gat, n3132gat, n3133gat, n3134gat, n3135gat, n3136gat, n3137gat, n3138gat, n3139gat, n3140gat, n3141gat, n3142gat, n3143gat, n3144gat, n3145gat, n3146gat, n3147gat, n3148gat, n3149gat, n3150gat, n3151gat, n3152gat;
wire clk, n3065gat, n3066gat, n3067gat, n3068gat, n3069gat, n3070gat, n3071gat, n3072gat, n3073gat, n3074gat, n3075gat, n3076gat, n3077gat, n3078gat, n3079gat, n3080gat, n3081gat, n3082gat, n3083gat, n3084gat, n3085gat, n3086gat, n3087gat, n3088gat, n3089gat, n3090gat, n3091gat, n3092gat, n3093gat, n3094gat, n3095gat, n3097gat, n3098gat, n3099gat, n3100gat;
wire n673gat, n398gat, n402gat, n919gat, n846gat, n394gat, n703gat, n722gat, n726gat, n2510gat, n271gat;
wire n160gat, n337gat, n842gat, n341gat, n2522gat, n2472gat, n2319gat, n1821gat, n1825gat, n2029gat, n1829gat;
wire n283gat, n165gat, n279gat, n1026gat, n275gat, n2476gat, n1068gat, n957gat, n861gat, n1294gat, n1241gat;
wire n1298gat, n865gat, n1080gat, n1148gat, n2468gat, n618gat, n491gat, n622gat, n626gat, n834gat, n707gat;
wire n838gat, n830gat, n614gat, n2526gat, n680gat, n816gat, n580gat, n824gat, n820gat, n883gat, n584gat;
wire n684gat, n699gat, n2464gat, n2399gat, n2343gat, n2203gat, n2562gat, n2207gat, n2626gat, n2490gat, n2622gat;
wire n2630gat, n2543gat, n2102gat, n1880gat, n1763gat, n2155gat, n1035gat, n1121gat, n1072gat, n1282gat, n1226gat;
wire n931gat, n1135gat, n1045gat, n1197gat, n2518gat, n667gat, n659gat, n553gat, n777gat, n561gat, n366gat;
wire n322gat, n318gat, n314gat, n2599gat, n2588gat, n2640gat, n2658gat, n2495gat, n2390gat, n2270gat, n2339gat;
wire n2502gat, n2634gat, n2506gat, n1834gat, n1767gat, n2084gat, n2143gat, n2061gat, n2139gat, n1899gat, n1850gat;
wire n2403gat, n2394gat, n2440gat, n2407gat, n2347gat, n1389gat, n2021gat, n1394gat, n1496gat, n2091gat, n1332gat;
wire n1740gat, n2179gat, n2190gat, n2135gat, n2262gat, n2182gat, n1433gat, n1316gat, n1363gat, n1312gat, n1775gat;
wire n1871gat, n2592gat, n1508gat, n1678gat, n2309gat, n2450gat, n2446gat, n2095gat, n2176gat, n2169gat, n2454gat;
wire n2040gat, n2044gat, n2037gat, n2025gat, n2099gat, n2266gat, n2033gat, n2110gat, n2125gat, n2121gat, n2117gat;
wire n1975gat, n2644gat, n156gat, n152gat, n331gat, n388gat, n463gat, n327gat, n384gat, n256gat, n470gat;
wire n148gat, n2458gat, n2514gat, n1771gat, n1336gat, n1748gat, n1675gat, n1807gat, n1340gat, n1456gat, n1525gat;
wire n1462gat, n1596gat, n1588gat, I1, n2717gat, n2715gat, I5, n2725gat, n2723gat, n296gat, I11;
wire n2768gat, I14, n2767gat, n373gat, I18, n2671gat, n2669gat, I23, n2845gat, n2844gat, I27;
wire n2668gat, I30, n2667gat, n856gat, I44, n672gat, I47, n2783gat, I50, n2782gat, n396gat;
wire I62, n2791gat, I65, n2790gat, I76, n401gat, n1645gat, I81, n2670gat, I92, n918gat;
wire n1553gat, I97, n2794gat, I100, n2793gat, I111, n845gat, n1559gat, n1643gat, n1651gat, n1562gat;
wire n1560gat, n1640gat, n1566gat, n1554gat, n1722gat, n392gat, I149, n702gat, n1319gat, n720gat, I171;
wire n725gat, n1447gat, n1627gat, I178, n721gat, n1380gat, n1628gat, n701gat, n1446gat, n1705gat, n1706gat;
wire I192, n2856gat, n2854gat, I196, n1218gat, I199, n2861gat, n2859gat, I203, n1219gat, I206;
wire n2864gat, n2862gat, I210, n1220gat, I214, n2860gat, I217, n1221gat, I220, n2863gat, I223;
wire n1222gat, I227, n2855gat, I230, n1223gat, n640gat, I237, n753gat, I240, n2716gat, I243;
wire n2869gat, n2867gat, I248, n2868gat, I253, n754gat, I256, n2724gat, I259, n2728gat, n2726gat;
wire I264, n2727gat, n422gat, I270, n755gat, n747gat, I275, n756gat, I278, n757gat, I282;
wire n758gat, n2508gat, I297, n2733gat, I300, n2732gat, I311, n270gat, I314, n263gat, I317;
wire n2777gat, I320, n2776gat, I331, n159gat, I334, n264gat, I337, n2736gat, I340, n2735gat;
wire I351, n336gat, I354, n265gat, n158gat, I359, n266gat, n335gat, I363, n267gat, n269gat;
wire I368, n268gat, n41gat, I375, n48gat, I378, n1018gat, I381, n2674gat, I384, n2673gat;
wire I395, n841gat, I398, n1019gat, I401, n1020gat, n840gat, I406, n1021gat, I409, n1022gat;
wire n724gat, I414, n1023gat, I420, n49gat, I423, n2780gat, I426, n2779gat, I437, n340gat;
wire I440, n480gat, I443, n481gat, I446, n393gat, I449, n482gat, I453, n483gat, I456;
wire n484gat, n339gat, I461, n485gat, n42gat, I468, n50gat, n162gat, I473, n51gat, I476;
wire n52gat, I480, n53gat, n2520gat, n1448gat, n1701gat, n1379gat, n1615gat, n1500gat, n1503gat, n1779gat;
wire I509, n2730gat, I512, n2729gat, n2470gat, n2317gat, n1819gat, n1823gat, n1816gat, n2027gat, I572;
wire n1828gat, I576, n2851gat, I579, n2850gat, I583, n2785gat, n92gat, n637gat, n293gat, I591;
wire n2722gat, I594, n2721gat, n297gat, I606, n282gat, I609, n172gat, I620, n164gat, I623;
wire n173gat, I634, n278gat, I637, n174gat, n163gat, I642, n175gat, n277gat, I646, n176gat;
wire n281gat, I651, n177gat, n54gat, I658, n60gat, I661, n911gat, I672, n1025gat, I675;
wire n912gat, I678, n913gat, n1024gat, I683, n914gat, n917gat, I687, n915gat, n844gat, I692;
wire n916gat, I698, n61gat, I709, n274gat, I712, n348gat, I715, n349gat, I718, n397gat;
wire I721, n350gat, n400gat, I726, n351gat, I729, n352gat, n273gat, I734, n353gat, n178gat;
wire I741, n62gat, n66gat, I746, n63gat, I749, n64gat, I753, n65gat, n2474gat, I768;
wire n2832gat, I771, n2831gat, n2731gat, I776, n2719gat, n2718gat, I790, n1067gat, I793, n949gat;
wire I796, n2839gat, n2838gat, n2775gat, I812, n956gat, I815, n950gat, I818, n2712gat, n2711gat;
wire n2734gat, I834, n860gat, I837, n951gat, n955gat, I842, n952gat, n859gat, I846, n953gat;
wire n1066gat, I851, n954gat, n857gat, I858, n938gat, n2792gat, I863, n2847gat, n2846gat, I877;
wire n1293gat, I880, n1233gat, n2672gat, I885, n2853gat, n2852gat, I899, n1240gat, I902, n1234gat;
wire I913, n1297gat, I916, n1235gat, n1239gat, I921, n1236gat, n1296gat, I925, n1237gat, n1292gat;
wire I930, n1238gat, I936, n939gat, n2778gat, I941, n2837gat, n2836gat, I955, n864gat, I958;
wire n1055gat, n2789gat, I963, n2841gat, n2840gat, I977, n1079gat, I980, n1056gat, n2781gat, I985;
wire n2843gat, n2842gat, I999, n1147gat, I1002, n1057gat, n1078gat, I1007, n1058gat, n1146gat, I1011;
wire n1059gat, n863gat, I1016, n1060gat, n928gat, I1023, n940gat, n858gat, I1028, n941gat, I1031;
wire n942gat, I1035, n943gat, n2466gat, n2720gat, n740gat, n2784gat, n743gat, n294gat, n374gat, n616gat;
wire I1067, n501gat, n489gat, I1079, n502gat, I1082, n617gat, I1085, n499gat, I1088, n490gat;
wire I1091, n500gat, n620gat, I1103, n738gat, n624gat, I1115, n737gat, I1118, n621gat, I1121;
wire n733gat, I1124, n625gat, I1127, n735gat, I1138, n833gat, I1141, n714gat, I1152, n706gat;
wire I1155, n715gat, I1166, n837gat, I1169, n716gat, n705gat, I1174, n717gat, n836gat, I1178;
wire n718gat, n832gat, I1183, n719gat, n515gat, I1190, n509gat, I1201, n829gat, I1204, n734gat;
wire n828gat, I1209, n736gat, I1216, n510gat, I1227, n613gat, I1230, n498gat, n612gat, I1236;
wire n503gat, n404gat, I1243, n511gat, n405gat, I1248, n512gat, I1251, n513gat, I1255, n514gat;
wire n2524gat, n17gat, n79gat, n219gat, n563gat, n289gat, n179gat, n188gat, n72gat, n111gat, I1302;
wire n679gat, I1305, n808gat, I1319, n815gat, I1322, n809gat, I1336, n579gat, I1339, n810gat;
wire n814gat, I1344, n811gat, n578gat, I1348, n812gat, n678gat, I1353, n813gat, n677gat, I1360;
wire n572gat, I1371, n823gat, I1374, n591gat, I1385, n819gat, I1388, n592gat, I1399, n882gat;
wire I1402, n593gat, n818gat, I1407, n594gat, n881gat, I1411, n595gat, n822gat, I1416, n596gat;
wire I1422, n573gat, I1436, n583gat, I1439, n691gat, I1450, n683gat, I1453, n692gat, I1464;
wire n698gat, I1467, n693gat, n682gat, I1472, n694gat, n697gat, I1476, n695gat, n582gat, I1481;
wire n696gat, n456gat, I1488, n574gat, n565gat, I1493, n575gat, I1496, n576gat, I1500, n577gat;
wire n2462gat, n2665gat, n2596gat, n189gat, n194gat, n21gat, I1538, n2398gat, n2353gat, I1550, n2342gat;
wire n2284gat, n2201gat, n2354gat, n2560gat, n2356gat, n2205gat, n2214gat, n2286gat, n2624gat, I1606, n2489gat;
wire I1617, n2621gat, n2533gat, I1630, n2629gat, n2486gat, n2541gat, n2429gat, n2432gat, I1655, n2101gat;
wire n1693gat, I1667, n1879gat, n1698gat, n1543gat, I1683, n1762gat, n1673gat, n1858gat, I1698, n2154gat;
wire n2488gat, I1703, n2625gat, n2530gat, I1708, n2542gat, n2482gat, n2426gat, n2153gat, n2341gat, n2355gat;
wire I1719, n2561gat, n2443gat, n2289gat, n2148gat, n855gat, n759gat, I1749, n1034gat, I1752, n1189gat;
wire n1075gat, I1766, n1120gat, I1769, n1190gat, n760gat, I1783, n1071gat, I1786, n1191gat, n1119gat;
wire I1791, n1192gat, n1070gat, I1795, n1193gat, n1033gat, I1800, n1194gat, n1183gat, I1807, n1274gat;
wire n644gat, n1280gat, n641gat, I1833, n1225gat, I1837, n1281gat, n1224gat, I1843, n1275gat, n761gat;
wire I1857, n930gat, I1860, n1206gat, n762gat, I1874, n1134gat, I1877, n1207gat, n643gat, I1891;
wire n1044gat, I1894, n1208gat, n1133gat, I1899, n1209gat, n1043gat, I1903, n1210gat, n929gat, I1908;
wire n1211gat, n1268gat, I1915, n1276gat, n1329gat, I1920, n1277gat, I1923, n1278gat, I1927, n1279gat;
wire n1284gat, n642gat, n1195gat, I1947, n1196gat, n2516gat, I1961, n3017gat, n851gat, n1725gat, n664gat;
wire n852gat, I1981, n666gat, n368gat, I1996, n658gat, I1999, n784gat, n662gat, I2014, n552gat;
wire I2017, n785gat, n661gat, I2032, n776gat, I2035, n786gat, n551gat, I2040, n787gat, n775gat;
wire I2044, n788gat, n657gat, I2049, n789gat, n35gat, I2056, n125gat, n558gat, n559gat, n371gat;
wire I2084, n365gat, I2088, n560gat, n364gat, I2094, n126gat, n663gat, I2109, n321gat, I2112;
wire n226gat, n370gat, I2127, n317gat, I2130, n227gat, n369gat, I2145, n313gat, I2148, n228gat;
wire n316gat, I2153, n229gat, n312gat, I2157, n230gat, n320gat, I2162, n231gat, n34gat, I2169;
wire n127gat, n133gat, I2174, n128gat, I2177, n129gat, I2181, n130gat, n665gat, n1601gat, n2597gat;
wire n2595gat, n2586gat, I2213, n2573gat, n2638gat, I2225, n2574gat, I2228, n2575gat, I2232, n2639gat;
wire I2235, n2576gat, I2238, n2577gat, I2242, n2578gat, I2248, n2582gat, I2251, n2206gat, I2254;
wire n2414gat, I2257, n2415gat, I2260, n2202gat, I2263, n2416gat, n2397gat, I2268, n2417gat, I2271;
wire n2418gat, I2275, n2419gat, I2281, n2585gat, n2656gat, n2493gat, n2388gat, I2316, n2389gat, I2319;
wire n2494gat, I2324, n2649gat, n2268gat, I2344, n2338gat, n2337gat, I2349, n2269gat, I2354, n2652gat;
wire n2500gat, n2620gat, n2612gat, I2372, n2606gat, n2532gat, I2376, n2607gat, n2540gat, I2380, n2608gat;
wire n2536gat, I2385, n2609gat, n2487gat, I2389, n2610gat, n2557gat, I2394, n2611gat, I2400, n2616gat;
wire I2403, n2550gat, I2414, n2633gat, I2417, n2551gat, I2420, n2552gat, n2632gat, I2425, n2553gat;
wire I2428, n2554gat, n2628gat, I2433, n2555gat, I2439, n2619gat, n2504gat, n2660gat, n1528gat, n1523gat;
wire n1592gat, n2666gat, n2422gat, n2290gat, n2081gat, n2285gat, n2359gat, n1414gat, n566gat, n1480gat, n1301gat;
wire n1150gat, n873gat, n2011gat, n1478gat, n875gat, n1410gat, n876gat, n1160gat, n1084gat, n983gat, n1482gat;
wire n1157gat, n985gat, n1530gat, n1307gat, n1085gat, n1479gat, n1348gat, n2217gat, n1591gat, n1437gat, n1832gat;
wire n1765gat, n1878gat, n1442gat, n1444gat, n1378gat, n1322gat, n1439gat, n1370gat, n1369gat, n1366gat, n1374gat;
wire n2162gat, n1450gat, n1427gat, n1603gat, n2082gat, n1449gat, n1590gat, n1248gat, n1418gat, n1306gat, n1353gat;
wire n1247gat, n1355gat, n1300gat, n1487gat, n1164gat, n1356gat, n1436gat, n1106gat, n1425gat, n1105gat, n1424gat;
wire n1309gat, I2672, n2142gat, n1788gat, I2684, n2060gat, n1786gat, I2696, n2138gat, n1839gat, n1897gat;
wire n1884gat, n1848gat, n1783gat, n1548gat, n1719gat, n2137gat, n1633gat, n2059gat, n1785gat, I2731, n1849gat;
wire n1784gat, n1716gat, n1635gat, n2401gat, n1989gat, n2392gat, n1918gat, I2771, n2439gat, n1986gat, n1866gat;
wire I2785, n2406gat, n2216gat, n2345gat, n1988gat, n1735gat, n1387gat, n1694gat, n1777gat, n1781gat, n2019gat;
wire n1549gat, n1551gat, I2837, n2346gat, n2152gat, n2405gat, n2351gat, I2843, n2402gat, n2212gat, I2847;
wire n2393gat, n1991gat, n1665gat, n1517gat, n1392gat, I2873, n1495gat, n1685gat, I2885, n2090gat, n1550gat;
wire n1552gat, n1330gat, n1738gat, I2915, n1739gat, n1925gat, n1917gat, n2141gat, n1787gat, n1717gat, n1859gat;
wire n1922gat, n1713gat, n1743gat, n1923gat, n1945gat, I2953, n2178gat, n1661gat, n1572gat, n2438gat, n2283gat;
wire n1520gat, n1580gat, n1990gat, I2978, n2189gat, I2989, n2134gat, I3000, n2261gat, n2128gat, n1836gat;
wire I3016, n2181gat, n1431gat, n1314gat, n1361gat, I3056, n1311gat, n1707gat, n1773gat, n1659gat, n1515gat;
wire n1736gat, n1658gat, n1724gat, n1662gat, n1656gat, n1670gat, n1569gat, n1568gat, n1727gat, n1797gat, n1730gat;
wire n1561gat, n1668gat, n1742gat, n1671gat, n1652gat, n1648gat, n1790gat, n2004gat, n1869gat, I3143, n2591gat;
wire n1584gat, n1714gat, n1718gat, I3163, n1507gat, n1396gat, I3168, n1393gat, n1409gat, I3174, n1898gat;
wire n1838gat, n1712gat, I3191, n1677gat, n2000gat, n2001gat, n1999gat, n2307gat, I3211, n3018gat, n2448gat;
wire n2661gat, n2444gat, I3235, n3019gat, n1310gat, n199gat, n195gat, n827gat, n2093gat, n2174gat, I3273;
wire n2168gat, n2452gat, n1691gat, I3287, n3020gat, I3290, n3021gat, I3293, n3022gat, n1699gat, I3297;
wire n3023gat, I3300, n3024gat, I3303, n3025gat, I3306, n3026gat, I3309, n3027gat, I3312, n3028gat;
wire I3315, n3029gat, I3318, n3030gat, n2260gat, n2257gat, n2188gat, n2187gat, I3336, n2039gat, I3339;
wire n1774gat, I3342, n1315gat, n2042gat, n2035gat, n2023gat, n2097gat, n1855gat, I3387, n3031gat, I3390;
wire n3032gat, n2256gat, I3394, n3033gat, n2251gat, n2184gat, I3401, n3034gat, n2133gat, n2131gat, n2049gat;
wire I3412, n3035gat, n2253gat, n2252gat, n2248gat, n2264gat, I3429, n2265gat, n2492gat, I3436, n3036gat;
wire n1709gat, n1845gat, n1891gat, n1963gat, n1886gat, n1968gat, n1629gat, n1631gat, n1711gat, n2200gat, n2437gat;
wire I3457, n3037gat, n1956gat, I3461, n3038gat, n1954gat, I3465, n3039gat, n1888gat, n2048gat, I3472;
wire n3040gat, n1969gat, n1893gat, n1892gat, I3483, n3041gat, n2056gat, I3491, n3042gat, I3494, n3043gat;
wire n1960gat, n1887gat, n1961gat, I3504, n3044gat, n2199gat, I3509, n3045gat, n2332gat, I3513, n3046gat;
wire n2259gat, n2328gat, I3520, n3047gat, n2151gat, n2209gat, I3530, n3048gat, n2052gat, n2058gat, I3539;
wire n3049gat, n2349gat, n2281gat, I3549, n3050gat, n2146gat, I3558, n3051gat, n2031gat, n2108gat, I3587;
wire n2124gat, n2123gat, n2119gat, n2115gat, I3610, n3052gat, I3621, n1974gat, n1955gat, n1970gat, n1973gat;
wire n2558gat, I3635, n3053gat, I3646, n2643gat, n2333gat, n2564gat, n2642gat, n2636gat, I3660, n3054gat;
wire n88gat, n375gat, I3677, n155gat, n253gat, n150gat, I3691, n151gat, n243gat, n233gat, n154gat;
wire n800gat, I3703, n3055gat, n235gat, I3713, n3056gat, n372gat, n329gat, I3736, n387gat, n334gat;
wire n386gat, I3742, n330gat, n1430gat, n1490gat, n452gat, I3754, n3057gat, n333gat, I3765, n3058gat;
wire I3777, n462gat, n325gat, n457gat, n461gat, n458gat, I3801, n3059gat, n144gat, I3808, n326gat;
wire n878gat, I3817, n3060gat, n382gat, I3831, n383gat, n134gat, I3841, n3061gat, n254gat, n252gat;
wire n468gat, I3867, n469gat, n381gat, I3876, n3062gat, n241gat, I3882, n255gat, n802gat, I3891;
wire n3063gat, n146gat, I3904, n147gat, n380gat, I3914, n3064gat, n69gat, n1885gat, I3923, n2707gat;
wire n16gat, n295gat, n11gat, n1889gat, I3935, n2700gat, n2051gat, I3941, n2680gat, n1350gat, I3945;
wire n2696gat, I3948, n2692gat, I3951, n2683gat, I3954, n2679gat, I3957, n2449gat, n1754gat, I3962;
wire n2827gat, n2590gat, n2456gat, n2512gat, n1544gat, n1769gat, n1683gat, n2167gat, n2013gat, n1791gat, n2691gat;
wire n1518gat, n2699gat, n2159gat, n2478gat, I4014, n2740gat, n2158gat, n2186gat, I4020, n2797gat, n2288gat;
wire n1513gat, n2537gat, n2442gat, n1334gat, I4055, n1747gat, I4067, n1674gat, n1403gat, I4081, n1806gat;
wire n1634gat, n1338gat, I4105, n1455gat, I4108, n1339gat, n1505gat, I4117, n2758gat, n2755gat, n1546gat;
wire I4122, n2752gat, n2748gat, n2012gat, n2002gat, I4129, n2858gat, n2857gat, I4135, n2766gat, I4138;
wire n2765gat, n1684gat, n1632gat, I4157, n1524gat, n1862gat, n1919gat, n1460gat, I4185, n1595gat, n1454gat;
wire n1468gat, I4194, n1461gat, n1477gat, n1594gat, I4212, n1587gat, n1681gat, I4222, n2751gat, n2747gat;
wire I4227, n2743gat, n2739gat, n1978gat, I4233, n2808gat, I4236, n2804gat, n517gat, n417gat, n413gat;
wire n412gat, n406gat, n407gat, n290gat, n527gat, n416gat, n528gat, n358gat, n639gat, n1111gat, n524gat;
wire n1112gat, n741gat, n633gat, n926gat, n670gat, n1123gat, n1007gat, n1006gat, I4309, n2814gat, I4312;
wire n2811gat, n1002gat, I4329, n2813gat, I4332, n2810gat, n888gat, I4349, n2818gat, I4352, n2816gat;
wire n898gat, I4369, n2817gat, I4372, n2815gat, n1179gat, I4389, n2824gat, I4392, n2821gat, n897gat;
wire I4409, n2823gat, I4412, n2820gat, n894gat, I4429, n2829gat, I4432, n2826gat, n1180gat, I4449;
wire n2828gat, I4452, n2825gat, n671gat, n628gat, n976gat, I4475, n2807gat, I4478, n2803gat, n2127gat;
wire I4482, n2682gat, I4485, n2678gat, n2046gat, I4489, n2681gat, I4492, n2677gat, n1708gat, I4496;
wire n2688gat, I4499, n2686gat, n455gat, n2237gat, I4506, n2763gat, n1782gat, I4512, n2760gat, n2325gat;
wire I4518, n2759gat, n2245gat, I4524, n2754gat, n2244gat, I4530, n2753gat, n2243gat, I4536, n2746gat;
wire n2246gat, I4542, n2745gat, n2384gat, I4548, n2738gat, n2385gat, I4554, n2737gat, n1286gat, I4558;
wire n2687gat, n2685gat, n1328gat, n1381gat, n1384gat, I4566, n2690gat, n1382gat, n1451gat, n1453gat, I4573;
wire n2689gat, n927gat, n925gat, n1452gat, I4580, n2698gat, n923gat, n921gat, n1890gat, I4587, n2697gat;
wire n850gat, n739gat, n1841gat, I4594, n2706gat, n922gat, n848gat, n2047gat, I4601, n2705gat, n924gat;
wire n849gat, n2050gat, I4608, n2796gat, n1118gat, n1032gat, n2054gat, I4615, n2795gat, I4620, n2806gat;
wire I4623, n2802gat, I4626, n1870gat, n1086gat, I4630, n2805gat, I4633, n2801gat, n67gat, n71gat;
wire n1840gat, I4642, n2809gat, n76gat, n14gat, n1842gat, I4651, n2819gat, I4654, n3104gat, I4657;
wire n3105gat, I4660, n3106gat, I4663, n3107gat, I4666, n3108gat, I4669, n3109gat, I4672, n3110gat;
wire I4675, n3111gat, I4678, n3112gat, I4681, n3113gat, I4684, n3114gat, I4687, n3115gat, I4690;
wire n3116gat, I4693, n3117gat, I4696, n3118gat, I4699, n3119gat, I4702, n3120gat, I4705, n3121gat;
wire I4708, n3122gat, I4711, n3123gat, I4714, n3124gat, I4717, n3125gat, I4720, n3126gat, I4723;
wire n3127gat, I4726, n3128gat, I4729, n3129gat, I4732, n3130gat, I4735, n3131gat, I4738, n3132gat;
wire I4741, n3133gat, I4744, n3134gat, I4747, n3135gat, I4750, n3136gat, I4753, n3137gat, I4756;
wire n3138gat, I4759, n3139gat, I4762, n3140gat, I4765, n3141gat, I4768, n3142gat, I4771, n3143gat;
wire I4774, n3144gat, I4777, n3145gat, I4780, n3146gat, I4783, n3147gat, I4786, n3148gat, I4789;
wire n3149gat, I4792, n3150gat, I4795, n3151gat, I4798, n3152gat, n2897gat, n1213gat, n2906gat, n2889gat;
wire n748gat, n258gat, n1013gat, n475gat, n43gat, n2786gat, n167gat, n906gat, n343gat, n55gat, n2914gat;
wire n2928gat, n2927gat, n944gat, n2896gat, n2922gat, n1228gat, n2894gat, n2921gat, n2895gat, n1050gat, n933gat;
wire n709gat, n728gat, n493gat, n504gat, I1277, I1278, n2913gat, n2920gat, n2905gat, n803gat, n586gat;
wire n2898gat, n686gat, n567gat, I1515, I1516, I1584, I1585, n2989gat, I1723, I1724, I1733;
wire I1734, n2918gat, n2952gat, n2919gat, n1184gat, n2910gat, n2907gat, n2970gat, n2911gat, n2912gat, n2909gat;
wire n1201gat, n1269gat, n2908gat, n2971gat, n2904gat, n2891gat, n2903gat, n2915gat, n779gat, n2901gat, n2890gat;
wire n2876gat, n2888gat, n2887gat, n2886gat, n221gat, n120gat, n3010gat, n3016gat, n2568gat, n2409gat, n2579gat;
wire n3014gat, n2880gat, n2646gat, n2601gat, n2545gat, n2613gat, n3013gat, n2930gat, n2957gat, n2975gat, n2974gat;
wire n2966gat, n2979gat, n2978gat, n2982gat, n2954gat, n2964gat, n2958gat, n2963gat, n2973gat, n2953gat, n2949gat;
wire n2934gat, n2959gat, n2977gat, I2720, I2721, I2735, I2736, I2812, I2813, I2831, I2832;
wire I2889, I2890, I2925, I2926, I2934, I2935, n2988gat, n2983gat, n2987gat, n2992gat, n2986gat;
wire n2991gat, I3148, I3149, I3178, I3179, n2981gat, n3000gat, n3004gat, n3003gat, n3001gat, n3006gat;
wire n3007gat, n2990gat, n2994gat, n2993gat, n2998gat, n2996gat, n3008gat, n3005gat, n2997gat, n3009gat, n3002gat;
wire n2995gat, n2999gat, n3011gat, n3015gat, n2874gat, n2917gat, n2878gat, n2892gat, n2885gat, n2900gat, n2883gat;
wire n2929gat, n2884gat, n2902gat, n2925gat, n2879gat, n2916gat, n2875gat, n2899gat, n2877gat, n2893gat, n2926gat;
wire n2882gat, n2924gat, n2881gat, n2923gat, n2710gat, n2704gat, n2684gat, n2830gat, I3999, I4000, n2695gat;
wire n2703gat, n2744gat, n2800gat, I4023, I4024, n2980gat, I4144, I4145, n2984gat, n2985gat, I4216;
wire I4217, n2931gat, n2943gat, n2941gat, n2946gat, n2960gat, n2950gat, n2969gat, n2933gat, n2935gat, n2942gat;
wire n2940gat, n2937gat, n2947gat, n2965gat, n2956gat, n2961gat, n2939gat, n2938gat, n2967gat, n2932gat, n2936gat;
wire n2948gat, n2968gat, n2955gat, n2944gat, n2945gat, n2962gat, n2951gat, n2764gat, n2762gat, n2761gat, n2757gat;
wire n2756gat, n2750gat, n2749gat, n2742gat, n2741gat, n2694gat, n2693gat, n2702gat, n2701gat, n2709gat, n2708gat;
wire n2799gat, n2798gat, n2812gat, n2822gat, n421gat, n648gat, n442gat, n1499gat, n1616gat, n1614gat, n1641gat;
wire n1642gat, n1556gat, n1557gat, n1639gat, n1605gat, n1555gat, n1558gat, n1256gat, n1117gat, n1618gat, n1114gat;
wire n1621gat, n1318gat, n1619gat, n1622gat, n1214gat, n1215gat, n1216gat, n1217gat, n745gat, n638gat, n423gat;
wire n362gat, n749gat, n750gat, n751gat, n752gat, n259gat, n260gat, n261gat, n262gat, n1014gat, n1015gat;
wire n1016gat, n1017gat, n476gat, n477gat, n478gat, n479gat, n44gat, n45gat, n46gat, n47gat, n1376gat;
wire n1617gat, n1377gat, n1624gat, n1113gat, n1501gat, n1623gat, n1620gat, n1827gat, n1817gat, n1935gat, n529gat;
wire n361gat, n168gat, n169gat, n170gat, n171gat, n907gat, n908gat, n909gat, n910gat, n344gat, n345gat;
wire n346gat, n347gat, n56gat, n57gat, n58gat, n59gat, n768gat, n655gat, n963gat, n868gat, n962gat;
wire n959gat, n945gat, n946gat, n947gat, n948gat, n647gat, n441gat, n967gat, n792gat, n1229gat, n1230gat;
wire n1231gat, n1232gat, n443gat, n439gat, n966gat, n790gat, n444gat, n440gat, n1051gat, n1052gat, n1053gat;
wire n1054gat, n934gat, n935gat, n936gat, n937gat, n746gat, n360gat, n710gat, n711gat, n712gat, n713gat;
wire n729gat, n730gat, n731gat, n732gat, n494gat, n495gat, n496gat, n497gat, n505gat, n506gat, n507gat;
wire n508gat, n564gat, n86gat, n78gat, n767gat, n286gat, n287gat, n288gat, n181gat, n182gat, n653gat;
wire n867gat, n771gat, n964gat, n961gat, n804gat, n805gat, n806gat, n807gat, n587gat, n588gat, n589gat;
wire n590gat, n447gat, n445gat, n687gat, n688gat, n689gat, n690gat, n568gat, n569gat, n570gat, n571gat;
wire n187gat, n197gat, n15gat, n22gat, n93gat, n769gat, n2534gat, n2430gat, n1606gat, n2239gat, n1934gat;
wire n1610gat, n1692gat, n2433gat, n2531gat, n2480gat, n2427gat, n2428gat, n1778gat, n1609gat, n1702gat, n1700gat;
wire n1604gat, n1076gat, n766gat, n1185gat, n1186gat, n1187gat, n1188gat, n645gat, n646gat, n1383gat, n1327gat;
wire n651gat, n652gat, n765gat, n1202gat, n1203gat, n1204gat, n1205gat, n1270gat, n1271gat, n1272gat, n1273gat;
wire n763gat, n1287gat, n1285gat, n853gat, n793gat, n854gat, n556gat, n795gat, n656gat, n794gat, n773gat;
wire n965gat, n960gat, n780gat, n781gat, n782gat, n783gat, n555gat, n450gat, n654gat, n557gat, n874gat;
wire n132gat, n649gat, n449gat, n791gat, n650gat, n774gat, n764gat, n222gat, n223gat, n224gat, n225gat;
wire n121gat, n122gat, n123gat, n124gat, n2460gat, n2423gat, n2594gat, n2569gat, n2570gat, n2571gat, n2572gat;
wire n2410gat, n2411gat, n2412gat, n2413gat, n2583gat, n2580gat, n2581gat, n2567gat, n2499gat, n299gat, n207gat;
wire n2650gat, n2647gat, n2648gat, n2602gat, n2603gat, n2604gat, n2605gat, n2546gat, n2547gat, n2548gat, n2549gat;
wire n2617gat, n2614gat, n2615gat, n2655gat, n2293gat, n2219gat, n1529gat, n1704gat, n2461gat, n2421gat, n1598gat;
wire n2218gat, n2358gat, n1415gat, n1153gat, n2292gat, n1416gat, n1151gat, n2306gat, n1481gat, n982gat, n2357gat;
wire n1347gat, n877gat, n1484gat, n1159gat, n2363gat, n1483gat, n1158gat, n2364gat, n1308gat, n1156gat, n2291gat;
wire n1349gat, n1155gat, n1154gat, n1703gat, n1608gat, n1411gat, n2223gat, n1438gat, n1625gat, n1626gat, n1831gat;
wire n1443gat, n1325gat, n1441gat, n1321gat, n1320gat, n1486gat, n1440gat, n1426gat, n1368gat, n1258gat, n1371gat;
wire n1365gat, n1373gat, n1372gat, n1367gat, n2220gat, n1423gat, n1498gat, n1504gat, n1607gat, n1494gat, n1502gat;
wire n1250gat, n1103gat, n1417gat, n1352gat, n1304gat, n1249gat, n1419gat, n1351gat, n1246gat, n1161gat, n1422gat;
wire n1303gat, n1291gat, n1245gat, n1485gat, n1302gat, n1163gat, n1102gat, n1354gat, n1360gat, n1435gat, n1101gat;
wire n996gat, n1359gat, n1421gat, n1104gat, n887gat, n1358gat, n1420gat, n1305gat, n1162gat, n1357gat, n1428gat;
wire n1794gat, n1796gat, n1792gat, n1865gat, n1861gat, n1793gat, n1406gat, n1780gat, n2016gat, n2664gat, n1666gat;
wire n1578gat, n1516gat, n1864gat, n1565gat, n1921gat, n1798gat, n1920gat, n1926gat, n1916gat, n1994gat, n1924gat;
wire n2078gat, n1690gat, n1660gat, n1576gat, n1733gat, n1582gat, n1577gat, n1581gat, n2129gat, n2079gat, n1695gat;
wire n2073gat, n1696gat, n1758gat, n1574gat, n1573gat, n1521gat, n1737gat, n1732gat, n1723gat, n1663gat, n1655gat;
wire n1647gat, n1667gat, n1570gat, n1646gat, n1575gat, n1728gat, n1650gat, n1801gat, n1731gat, n1649gat, n1571gat;
wire n1563gat, n1734gat, n1669gat, n1654gat, n1657gat, n1653gat, n1729gat, n1644gat, n1726gat, n1929gat, n2009gat;
wire n1413gat, n1636gat, n1401gat, n1408gat, n1476gat, n1407gat, n1412gat, n2663gat, n2662gat, n2238gat, n87gat;
wire n200gat, n184gat, n196gat, n204gat, n2163gat, n2258gat, n2255gat, n2015gat, n2017gat, n2018gat, n2014gat;
wire n2194gat, n2192gat, n2185gat, n2132gat, n2130gat, n2057gat, n2250gat, n2249gat, n2329gat, n1958gat, n1895gat;
wire n1710gat, n1630gat, n2195gat, n2556gat, n2539gat, n1894gat, n1847gat, n1846gat, n2436gat, n2055gat, n1967gat;
wire n2387gat, n1959gat, n1957gat, n2330gat, n2147gat, n2498gat, n2193gat, n2211gat, n2210gat, n2396gat, n2053gat;
wire n1964gat, n2198gat, n2215gat, n2350gat, n2282gat, n2197gat, n2213gat, n2150gat, n2149gat, n2196gat, n1882gat;
wire n1962gat, n1896gat, n1972gat, n1971gat, n2559gat, n2331gat, n2352gat, n2566gat, n2565gat, n2637gat, n84gat;
wire n89gat, n110gat, n1074gat, n141gat, n38gat, n37gat, n872gat, n234gat, n137gat, n378gat, n377gat;
wire n869gat, n212gat, n250gat, n249gat, n248gat, n453gat, n448gat, n974gat, n251gat, n244gat, n973gat;
wire n870gat, n975gat, n246gat, n245gat, n460gat, n459gat, n972gat, n969gat, n971gat, n247gat, n145gat;
wire n143gat, n970gat, n968gat, n772gat, n142gat, n40gat, n39gat, n451gat, n446gat, n139gat, n136gat;
wire n391gat, n390gat, n1083gat, n1077gat, n140gat, n242gat, n240gat, n871gat, n797gat, n324gat, n238gat;
wire n237gat, n1082gat, n796gat, n85gat, n180gat, n68gat, n186gat, n357gat, n82gat, n12gat, n1599gat;
wire n1613gat, n1756gat, n1586gat, n1755gat, n2538gat, n2483gat, n1391gat, n1471gat, n1469gat, n1472gat, n1927gat;
wire n1470gat, n1402gat, n1400gat, n1567gat, n1399gat, n1564gat, n1600gat, n1519gat, n1397gat, n1398gat, n2008gat;
wire n2005gat, n1818gat, n1759gat, n1686gat, n1533gat, n1863gat, n1860gat, n1915gat, n1510gat, n1800gat, n1459gat;
wire n1458gat, n1532gat, n1467gat, n1466gat, n1531gat, n1593gat, n1602gat, n1761gat, n1760gat, n1721gat, n520gat;
wire n519gat, n518gat, n418gat, n411gat, n522gat, n516gat, n410gat, n354gat, n355gat, n408gat, n526gat;
wire n531gat, n530gat, n525gat, n356gat, n415gat, n521gat, n532gat, n359gat, n420gat, n523gat, n634gat;
wire n414gat, n635gat, n1100gat, n630gat, n994gat, n629gat, n989gat, n632gat, n880gat, n636gat, n801gat;
wire n879gat, n1003gat, n1255gat, n1012gat, n905gat, n1009gat, n409gat, n292gat, n291gat, n419gat, n902gat;
wire n1099gat, n998gat, n995gat, n980gat, n1001gat, n1175gat, n1174gat, n1243gat, n1171gat, n999gat, n1244gat;
wire n1323gat, n1264gat, n1265gat, n892gat, n981gat, n890gat, n889gat, n886gat, n891gat, n904gat, n903gat;
wire n1254gat, n1008gat, n900gat, n1152gat, n1092gat, n997gat, n993gat, n895gat, n1094gat, n1093gat, n988gat;
wire n984gat, n1178gat, n1267gat, n1257gat, n1253gat, n1266gat, n1116gat, n1375gat, n1324gat, n1200gat, n1172gat;
wire n899gat, n1091gat, n1088gat, n992gat, n987gat, n896gat, n1262gat, n1260gat, n1251gat, n1259gat, n901gat;
wire n1098gat, n1090gat, n986gat, n885gat, n893gat, n1097gat, n1089gat, n1087gat, n991gat, n1177gat, n1212gat;
wire n1326gat, n1261gat, n1263gat, n1115gat, n977gat, n631gat, n1096gat, n1095gat, n990gat, n979gat, n978gat;
wire n1004gat, n1199gat, n1176gat, n1173gat, n1252gat, n1000gat, n1029gat, n1028gat, n1031gat, n1030gat, n1011gat;
wire n1181gat, n1010gat, n1005gat, n1182gat, n1757gat, n1745gat, n73gat, n70gat, n77gat, n13gat;
wire line1, line2, line3, line4, line5, line6, line7, line8, line9, line10, line11;
wire line12, line13, line14, line15, line16, line17, line18, line19, line20, line21, line22;
wire line23, line24, line25, line26, line27, line28, line29, line30, line31, line32, line33;
wire line34, line35, line36, line37, line38, line39, line40, line41, line42, line43, line44;
wire line45, line46, line47, line48, line49, line50, line51, line52, line53, line54, line55;
wire line56, line57, line58, line59, line60, line61, line62, line63, line64, line65, line66;
wire line67, line68, line69, line70, line71, line72, line73, line74, line75, line76, line77;
wire line78, line79, line80, line81, line82, line83, line84, line85, line86, line87, line88;
wire line89, line90, line91, line92, line93, line94, line95, line96, line97, line98, line99;
wire line100, line101, line102, line103, line104, line105, line106, line107, line108, line109, line110;
wire line111, line112, line113, line114, line115, line116, line117, line118, line119, line120, line121;
wire line122, line123, line124, line125, line126, line127, line128, line129, line130, line131, line132;
wire line133, line134, line135, line136, line137, line138, line139, line140, line141, line142, line143;
wire line144, line145, line146, line147, line148, line149, line150, line151, line152, line153, line154;
wire line155, line156, line157, line158, line159, line160, line161, line162, line163, line164, line165;
wire line166, line167, line168, line169, line170, line171, line172, line173, line174, line175, line176;
wire line177, line178, line179;
DFFX1 gate1(.Q (n673gat), .QB (line1), .D(n2897gat), .CK(clk));
DFFX1 gate2(.Q (n398gat), .QB (line2), .D(n2782gat), .CK(clk));
DFFX1 gate3(.Q (n402gat), .QB (line3), .D(n2790gat), .CK(clk));
DFFX1 gate4(.Q (n919gat), .QB (line4), .D(n2670gat), .CK(clk));
DFFX1 gate5(.Q (n846gat), .QB (line5), .D(n2793gat), .CK(clk));
DFFX1 gate6(.Q (n394gat), .QB (line6), .D(n2782gat), .CK(clk));
DFFX1 gate7(.Q (n703gat), .QB (line7), .D(n2790gat), .CK(clk));
DFFX1 gate8(.Q (n722gat), .QB (line8), .D(n2670gat), .CK(clk));
DFFX1 gate9(.Q (n726gat), .QB (line9), .D(n2793gat), .CK(clk));
DFFX1 gate10(.Q (n2510gat), .QB (line10), .D(n748gat), .CK(clk));
DFFX1 gate11(.Q (n271gat), .QB (line11), .D(n2732gat), .CK(clk));
DFFX1 gate12(.Q (n160gat), .QB (line12), .D(n2776gat), .CK(clk));
DFFX1 gate13(.Q (n337gat), .QB (line13), .D(n2735gat), .CK(clk));
DFFX1 gate14(.Q (n842gat), .QB (line14), .D(n2673gat), .CK(clk));
DFFX1 gate15(.Q (n341gat), .QB (line15), .D(n2779gat), .CK(clk));
DFFX1 gate16(.Q (n2522gat), .QB (line16), .D(n43gat), .CK(clk));
DFFX1 gate17(.Q (n2472gat), .QB (line17), .D(n1620gat), .CK(clk));
DFFX1 gate18(.Q (n2319gat), .QB (line18), .D(n2470gat), .CK(clk));
DFFX1 gate19(.Q (n1821gat), .QB (line19), .D(n1827gat), .CK(clk));
DFFX1 gate20(.Q (n1825gat), .QB (line20), .D(n1827gat), .CK(clk));
DFFX1 gate21(.Q (n2029gat), .QB (line21), .D(n1816gat), .CK(clk));
DFFX1 gate22(.Q (n1829gat), .QB (line22), .D(n2027gat), .CK(clk));
DFFX1 gate23(.Q (n283gat), .QB (line23), .D(n2732gat), .CK(clk));
DFFX1 gate24(.Q (n165gat), .QB (line24), .D(n2776gat), .CK(clk));
DFFX1 gate25(.Q (n279gat), .QB (line25), .D(n2735gat), .CK(clk));
DFFX1 gate26(.Q (n1026gat), .QB (line26), .D(n2673gat), .CK(clk));
DFFX1 gate27(.Q (n275gat), .QB (line27), .D(n2779gat), .CK(clk));
DFFX1 gate28(.Q (n2476gat), .QB (line28), .D(n55gat), .CK(clk));
DFFX1 gate29(.Q (n1068gat), .QB (line29), .D(n2914gat), .CK(clk));
DFFX1 gate30(.Q (n957gat), .QB (line30), .D(n2928gat), .CK(clk));
DFFX1 gate31(.Q (n861gat), .QB (line31), .D(n2927gat), .CK(clk));
DFFX1 gate32(.Q (n1294gat), .QB (line32), .D(n2896gat), .CK(clk));
DFFX1 gate33(.Q (n1241gat), .QB (line33), .D(n2922gat), .CK(clk));
DFFX1 gate34(.Q (n1298gat), .QB (line34), .D(n2897gat), .CK(clk));
DFFX1 gate35(.Q (n865gat), .QB (line35), .D(n2894gat), .CK(clk));
DFFX1 gate36(.Q (n1080gat), .QB (line36), .D(n2921gat), .CK(clk));
DFFX1 gate37(.Q (n1148gat), .QB (line37), .D(n2895gat), .CK(clk));
DFFX1 gate38(.Q (n2468gat), .QB (line38), .D(n933gat), .CK(clk));
DFFX1 gate39(.Q (n618gat), .QB (line39), .D(n2790gat), .CK(clk));
DFFX1 gate40(.Q (n491gat), .QB (line40), .D(n2782gat), .CK(clk));
DFFX1 gate41(.Q (n622gat), .QB (line41), .D(n2793gat), .CK(clk));
DFFX1 gate42(.Q (n626gat), .QB (line42), .D(n2670gat), .CK(clk));
DFFX1 gate43(.Q (n834gat), .QB (line43), .D(n3064gat), .CK(clk));
DFFX1 gate44(.Q (n707gat), .QB (line44), .D(n3055gat), .CK(clk));
DFFX1 gate45(.Q (n838gat), .QB (line45), .D(n3063gat), .CK(clk));
DFFX1 gate46(.Q (n830gat), .QB (line46), .D(n3062gat), .CK(clk));
DFFX1 gate47(.Q (n614gat), .QB (line47), .D(n3056gat), .CK(clk));
DFFX1 gate48(.Q (n2526gat), .QB (line48), .D(n504gat), .CK(clk));
DFFX1 gate49(.Q (n680gat), .QB (line49), .D(n2913gat), .CK(clk));
DFFX1 gate50(.Q (n816gat), .QB (line50), .D(n2920gat), .CK(clk));
DFFX1 gate51(.Q (n580gat), .QB (line51), .D(n2905gat), .CK(clk));
DFFX1 gate52(.Q (n824gat), .QB (line52), .D(n3057gat), .CK(clk));
DFFX1 gate53(.Q (n820gat), .QB (line53), .D(n3059gat), .CK(clk));
DFFX1 gate54(.Q (n883gat), .QB (line54), .D(n3058gat), .CK(clk));
DFFX1 gate55(.Q (n584gat), .QB (line55), .D(n2898gat), .CK(clk));
DFFX1 gate56(.Q (n684gat), .QB (line56), .D(n3060gat), .CK(clk));
DFFX1 gate57(.Q (n699gat), .QB (line57), .D(n3061gat), .CK(clk));
DFFX1 gate58(.Q (n2464gat), .QB (line58), .D(n567gat), .CK(clk));
DFFX1 gate59(.Q (n2399gat), .QB (line59), .D(n3048gat), .CK(clk));
DFFX1 gate60(.Q (n2343gat), .QB (line60), .D(n3049gat), .CK(clk));
DFFX1 gate61(.Q (n2203gat), .QB (line61), .D(n3051gat), .CK(clk));
DFFX1 gate62(.Q (n2562gat), .QB (line62), .D(n3047gat), .CK(clk));
DFFX1 gate63(.Q (n2207gat), .QB (line63), .D(n3050gat), .CK(clk));
DFFX1 gate64(.Q (n2626gat), .QB (line64), .D(n3040gat), .CK(clk));
DFFX1 gate65(.Q (n2490gat), .QB (line65), .D(n3044gat), .CK(clk));
DFFX1 gate66(.Q (n2622gat), .QB (line66), .D(n3042gat), .CK(clk));
DFFX1 gate67(.Q (n2630gat), .QB (line67), .D(n3037gat), .CK(clk));
DFFX1 gate68(.Q (n2543gat), .QB (line68), .D(n3041gat), .CK(clk));
DFFX1 gate69(.Q (n2102gat), .QB (line69), .D(n1606gat), .CK(clk));
DFFX1 gate70(.Q (n1880gat), .QB (line70), .D(n3052gat), .CK(clk));
DFFX1 gate71(.Q (n1763gat), .QB (line71), .D(n1610gat), .CK(clk));
DFFX1 gate72(.Q (n2155gat), .QB (line72), .D(n1858gat), .CK(clk));
DFFX1 gate73(.Q (n1035gat), .QB (line73), .D(n2918gat), .CK(clk));
DFFX1 gate74(.Q (n1121gat), .QB (line74), .D(n2952gat), .CK(clk));
DFFX1 gate75(.Q (n1072gat), .QB (line75), .D(n2919gat), .CK(clk));
DFFX1 gate76(.Q (n1282gat), .QB (line76), .D(n2910gat), .CK(clk));
DFFX1 gate77(.Q (n1226gat), .QB (line77), .D(n2907gat), .CK(clk));
DFFX1 gate78(.Q (n931gat), .QB (line78), .D(n2911gat), .CK(clk));
DFFX1 gate79(.Q (n1135gat), .QB (line79), .D(n2912gat), .CK(clk));
DFFX1 gate80(.Q (n1045gat), .QB (line80), .D(n2909gat), .CK(clk));
DFFX1 gate81(.Q (n1197gat), .QB (line81), .D(n2908gat), .CK(clk));
DFFX1 gate82(.Q (n2518gat), .QB (line82), .D(n2971gat), .CK(clk));
DFFX1 gate83(.Q (n667gat), .QB (line83), .D(n2904gat), .CK(clk));
DFFX1 gate84(.Q (n659gat), .QB (line84), .D(n2891gat), .CK(clk));
DFFX1 gate85(.Q (n553gat), .QB (line85), .D(n2903gat), .CK(clk));
DFFX1 gate86(.Q (n777gat), .QB (line86), .D(n2915gat), .CK(clk));
DFFX1 gate87(.Q (n561gat), .QB (line87), .D(n2901gat), .CK(clk));
DFFX1 gate88(.Q (n366gat), .QB (line88), .D(n2890gat), .CK(clk));
DFFX1 gate89(.Q (n322gat), .QB (line89), .D(n2888gat), .CK(clk));
DFFX1 gate90(.Q (n318gat), .QB (line90), .D(n2887gat), .CK(clk));
DFFX1 gate91(.Q (n314gat), .QB (line91), .D(n2886gat), .CK(clk));
DFFX1 gate92(.Q (n2599gat), .QB (line92), .D(n3010gat), .CK(clk));
DFFX1 gate93(.Q (n2588gat), .QB (line93), .D(n3016gat), .CK(clk));
DFFX1 gate94(.Q (n2640gat), .QB (line94), .D(n3054gat), .CK(clk));
DFFX1 gate95(.Q (n2658gat), .QB (line95), .D(n2579gat), .CK(clk));
DFFX1 gate96(.Q (n2495gat), .QB (line96), .D(n3036gat), .CK(clk));
DFFX1 gate97(.Q (n2390gat), .QB (line97), .D(n3034gat), .CK(clk));
DFFX1 gate98(.Q (n2270gat), .QB (line98), .D(n3031gat), .CK(clk));
DFFX1 gate99(.Q (n2339gat), .QB (line99), .D(n3035gat), .CK(clk));
DFFX1 gate100(.Q (n2502gat), .QB (line100), .D(n2646gat), .CK(clk));
DFFX1 gate101(.Q (n2634gat), .QB (line101), .D(n3053gat), .CK(clk));
DFFX1 gate102(.Q (n2506gat), .QB (line102), .D(n2613gat), .CK(clk));
DFFX1 gate103(.Q (n1834gat), .QB (line103), .D(n1625gat), .CK(clk));
DFFX1 gate104(.Q (n1767gat), .QB (line104), .D(n1626gat), .CK(clk));
DFFX1 gate105(.Q (n2084gat), .QB (line105), .D(n1603gat), .CK(clk));
DFFX1 gate106(.Q (n2143gat), .QB (line106), .D(n2541gat), .CK(clk));
DFFX1 gate107(.Q (n2061gat), .QB (line107), .D(n2557gat), .CK(clk));
DFFX1 gate108(.Q (n2139gat), .QB (line108), .D(n2487gat), .CK(clk));
DFFX1 gate109(.Q (n1899gat), .QB (line109), .D(n2532gat), .CK(clk));
DFFX1 gate110(.Q (n1850gat), .QB (line110), .D(n2628gat), .CK(clk));
DFFX1 gate111(.Q (n2403gat), .QB (line111), .D(n2397gat), .CK(clk));
DFFX1 gate112(.Q (n2394gat), .QB (line112), .D(n2341gat), .CK(clk));
DFFX1 gate113(.Q (n2440gat), .QB (line113), .D(n2560gat), .CK(clk));
DFFX1 gate114(.Q (n2407gat), .QB (line114), .D(n2205gat), .CK(clk));
DFFX1 gate115(.Q (n2347gat), .QB (line115), .D(n2201gat), .CK(clk));
DFFX1 gate116(.Q (n1389gat), .QB (line116), .D(n1793gat), .CK(clk));
DFFX1 gate117(.Q (n2021gat), .QB (line117), .D(n1781gat), .CK(clk));
DFFX1 gate118(.Q (n1394gat), .QB (line118), .D(n1516gat), .CK(clk));
DFFX1 gate119(.Q (n1496gat), .QB (line119), .D(n1392gat), .CK(clk));
DFFX1 gate120(.Q (n2091gat), .QB (line120), .D(n1685gat), .CK(clk));
DFFX1 gate121(.Q (n1332gat), .QB (line121), .D(n1565gat), .CK(clk));
DFFX1 gate122(.Q (n1740gat), .QB (line122), .D(n1330gat), .CK(clk));
DFFX1 gate123(.Q (n2179gat), .QB (line123), .D(n1945gat), .CK(clk));
DFFX1 gate124(.Q (n2190gat), .QB (line124), .D(n2268gat), .CK(clk));
DFFX1 gate125(.Q (n2135gat), .QB (line125), .D(n2337gat), .CK(clk));
DFFX1 gate126(.Q (n2262gat), .QB (line126), .D(n2388gat), .CK(clk));
DFFX1 gate127(.Q (n2182gat), .QB (line127), .D(n1836gat), .CK(clk));
DFFX1 gate128(.Q (n1433gat), .QB (line128), .D(n2983gat), .CK(clk));
DFFX1 gate129(.Q (n1316gat), .QB (line129), .D(n1431gat), .CK(clk));
DFFX1 gate130(.Q (n1363gat), .QB (line130), .D(n1314gat), .CK(clk));
DFFX1 gate131(.Q (n1312gat), .QB (line131), .D(n1361gat), .CK(clk));
DFFX1 gate132(.Q (n1775gat), .QB (line132), .D(n1696gat), .CK(clk));
DFFX1 gate133(.Q (n1871gat), .QB (line133), .D(n2009gat), .CK(clk));
DFFX1 gate134(.Q (n2592gat), .QB (line134), .D(n1773gat), .CK(clk));
DFFX1 gate135(.Q (n1508gat), .QB (line135), .D(n1636gat), .CK(clk));
DFFX1 gate136(.Q (n1678gat), .QB (line136), .D(n1712gat), .CK(clk));
DFFX1 gate137(.Q (n2309gat), .QB (line137), .D(n3000gat), .CK(clk));
DFFX1 gate138(.Q (n2450gat), .QB (line138), .D(n2307gat), .CK(clk));
DFFX1 gate139(.Q (n2446gat), .QB (line139), .D(n2661gat), .CK(clk));
DFFX1 gate140(.Q (n2095gat), .QB (line140), .D(n827gat), .CK(clk));
DFFX1 gate141(.Q (n2176gat), .QB (line141), .D(n2093gat), .CK(clk));
DFFX1 gate142(.Q (n2169gat), .QB (line142), .D(n2174gat), .CK(clk));
DFFX1 gate143(.Q (n2454gat), .QB (line143), .D(n2163gat), .CK(clk));
DFFX1 gate144(.Q (n2040gat), .QB (line144), .D(n1777gat), .CK(clk));
DFFX1 gate145(.Q (n2044gat), .QB (line145), .D(n2015gat), .CK(clk));
DFFX1 gate146(.Q (n2037gat), .QB (line146), .D(n2042gat), .CK(clk));
DFFX1 gate147(.Q (n2025gat), .QB (line147), .D(n2017gat), .CK(clk));
DFFX1 gate148(.Q (n2099gat), .QB (line148), .D(n2023gat), .CK(clk));
DFFX1 gate149(.Q (n2266gat), .QB (line149), .D(n2493gat), .CK(clk));
DFFX1 gate150(.Q (n2033gat), .QB (line150), .D(n2035gat), .CK(clk));
DFFX1 gate151(.Q (n2110gat), .QB (line151), .D(n2031gat), .CK(clk));
DFFX1 gate152(.Q (n2125gat), .QB (line152), .D(n2108gat), .CK(clk));
DFFX1 gate153(.Q (n2121gat), .QB (line153), .D(n2123gat), .CK(clk));
DFFX1 gate154(.Q (n2117gat), .QB (line154), .D(n2119gat), .CK(clk));
DFFX1 gate155(.Q (n1975gat), .QB (line155), .D(n2632gat), .CK(clk));
DFFX1 gate156(.Q (n2644gat), .QB (line156), .D(n2638gat), .CK(clk));
DFFX1 gate157(.Q (n156gat), .QB (line157), .D(n612gat), .CK(clk));
DFFX1 gate158(.Q (n152gat), .QB (line158), .D(n705gat), .CK(clk));
DFFX1 gate159(.Q (n331gat), .QB (line159), .D(n822gat), .CK(clk));
DFFX1 gate160(.Q (n388gat), .QB (line160), .D(n881gat), .CK(clk));
DFFX1 gate161(.Q (n463gat), .QB (line161), .D(n818gat), .CK(clk));
DFFX1 gate162(.Q (n327gat), .QB (line162), .D(n682gat), .CK(clk));
DFFX1 gate163(.Q (n384gat), .QB (line163), .D(n697gat), .CK(clk));
DFFX1 gate164(.Q (n256gat), .QB (line164), .D(n836gat), .CK(clk));
DFFX1 gate165(.Q (n470gat), .QB (line165), .D(n828gat), .CK(clk));
DFFX1 gate166(.Q (n148gat), .QB (line166), .D(n832gat), .CK(clk));
DFFX1 gate167(.Q (n2458gat), .QB (line167), .D(n2590gat), .CK(clk));
DFFX1 gate168(.Q (n2514gat), .QB (line168), .D(n2456gat), .CK(clk));
DFFX1 gate169(.Q (n1771gat), .QB (line169), .D(n1613gat), .CK(clk));
DFFX1 gate170(.Q (n1336gat), .QB (line170), .D(n1391gat), .CK(clk));
DFFX1 gate171(.Q (n1748gat), .QB (line171), .D(n1927gat), .CK(clk));
DFFX1 gate172(.Q (n1675gat), .QB (line172), .D(n1713gat), .CK(clk));
DFFX1 gate173(.Q (n1807gat), .QB (line173), .D(n1717gat), .CK(clk));
DFFX1 gate174(.Q (n1340gat), .QB (line174), .D(n1567gat), .CK(clk));
DFFX1 gate175(.Q (n1456gat), .QB (line175), .D(n1564gat), .CK(clk));
DFFX1 gate176(.Q (n1525gat), .QB (line176), .D(n1632gat), .CK(clk));
DFFX1 gate177(.Q (n1462gat), .QB (line177), .D(n1915gat), .CK(clk));
DFFX1 gate178(.Q (n1596gat), .QB (line178), .D(n1800gat), .CK(clk));
DFFX1 gate179(.Q (n1588gat), .QB (line179), .D(n1593gat), .CK(clk));
INVX1 gate180(.O (I1), .I (n3088gat));
INVX1 gate181(.O (n2717gat), .I (I1));
INVX1 gate182(.O (n2715gat), .I (n2717gat));
INVX1 gate183(.O (I5), .I (n3087gat));
INVX1 gate184(.O (n2725gat), .I (I5));
INVX1 gate185(.O (n2723gat), .I (n2725gat));
INVX1 gate186(.O (n296gat), .I (n421gat));
INVX1 gate187(.O (I11), .I (n3093gat));
INVX1 gate188(.O (n2768gat), .I (I11));
INVX1 gate189(.O (I14), .I (n2768gat));
INVX1 gate190(.O (n2767gat), .I (I14));
INVX1 gate191(.O (n373gat), .I (n2767gat));
INVX1 gate192(.O (I18), .I (n3072gat));
INVX1 gate193(.O (n2671gat), .I (I18));
INVX1 gate194(.O (n2669gat), .I (n2671gat));
INVX1 gate195(.O (I23), .I (n3081gat));
INVX1 gate196(.O (n2845gat), .I (I23));
INVX1 gate197(.O (n2844gat), .I (n2845gat));
INVX1 gate198(.O (I27), .I (n3095gat));
INVX1 gate199(.O (n2668gat), .I (I27));
INVX1 gate200(.O (I30), .I (n2668gat));
INVX1 gate201(.O (n2667gat), .I (I30));
INVX1 gate202(.O (n856gat), .I (n2667gat));
INVX1 gate203(.O (I44), .I (n673gat));
INVX1 gate204(.O (n672gat), .I (I44));
INVX1 gate205(.O (I47), .I (n3069gat));
INVX1 gate206(.O (n2783gat), .I (I47));
INVX1 gate207(.O (I50), .I (n2783gat));
INVX1 gate208(.O (n2782gat), .I (I50));
INVX1 gate209(.O (n396gat), .I (n398gat));
INVX1 gate210(.O (I62), .I (n3070gat));
INVX1 gate211(.O (n2791gat), .I (I62));
INVX1 gate212(.O (I65), .I (n2791gat));
INVX1 gate213(.O (n2790gat), .I (I65));
INVX1 gate214(.O (I76), .I (n402gat));
INVX1 gate215(.O (n401gat), .I (I76));
INVX1 gate216(.O (n1645gat), .I (n1499gat));
INVX1 gate217(.O (I81), .I (n2671gat));
INVX1 gate218(.O (n2670gat), .I (I81));
INVX1 gate219(.O (I92), .I (n919gat));
INVX1 gate220(.O (n918gat), .I (I92));
INVX1 gate221(.O (n1553gat), .I (n1616gat));
INVX1 gate222(.O (I97), .I (n3071gat));
INVX1 gate223(.O (n2794gat), .I (I97));
INVX1 gate224(.O (I100), .I (n2794gat));
INVX1 gate225(.O (n2793gat), .I (I100));
INVX1 gate226(.O (I111), .I (n846gat));
INVX1 gate227(.O (n845gat), .I (I111));
INVX1 gate228(.O (n1559gat), .I (n1614gat));
INVX1 gate229(.O (n1643gat), .I (n1641gat));
INVX1 gate230(.O (n1651gat), .I (n1642gat));
INVX1 gate231(.O (n1562gat), .I (n1556gat));
INVX1 gate232(.O (n1560gat), .I (n1557gat));
INVX1 gate233(.O (n1640gat), .I (n1639gat));
INVX1 gate234(.O (n1566gat), .I (n1605gat));
INVX1 gate235(.O (n1554gat), .I (n1555gat));
INVX1 gate236(.O (n1722gat), .I (n1558gat));
INVX1 gate237(.O (n392gat), .I (n394gat));
INVX1 gate238(.O (I149), .I (n703gat));
INVX1 gate239(.O (n702gat), .I (I149));
INVX1 gate240(.O (n1319gat), .I (n1256gat));
INVX1 gate241(.O (n720gat), .I (n722gat));
INVX1 gate242(.O (I171), .I (n726gat));
INVX1 gate243(.O (n725gat), .I (I171));
INVX1 gate244(.O (n1447gat), .I (n1117gat));
INVX1 gate245(.O (n1627gat), .I (n1618gat));
INVX1 gate246(.O (I178), .I (n722gat));
INVX1 gate247(.O (n721gat), .I (I178));
INVX1 gate248(.O (n1380gat), .I (n1114gat));
INVX1 gate249(.O (n1628gat), .I (n1621gat));
INVX1 gate250(.O (n701gat), .I (n703gat));
INVX1 gate251(.O (n1446gat), .I (n1318gat));
INVX1 gate252(.O (n1705gat), .I (n1619gat));
INVX1 gate253(.O (n1706gat), .I (n1622gat));
INVX1 gate254(.O (I192), .I (n3083gat));
INVX1 gate255(.O (n2856gat), .I (I192));
INVX1 gate256(.O (n2854gat), .I (n2856gat));
INVX1 gate257(.O (I196), .I (n2854gat));
INVX1 gate258(.O (n1218gat), .I (I196));
INVX1 gate259(.O (I199), .I (n3085gat));
INVX1 gate260(.O (n2861gat), .I (I199));
INVX1 gate261(.O (n2859gat), .I (n2861gat));
INVX1 gate262(.O (I203), .I (n2859gat));
INVX1 gate263(.O (n1219gat), .I (I203));
INVX1 gate264(.O (I206), .I (n3084gat));
INVX1 gate265(.O (n2864gat), .I (I206));
INVX1 gate266(.O (n2862gat), .I (n2864gat));
INVX1 gate267(.O (I210), .I (n2862gat));
INVX1 gate268(.O (n1220gat), .I (I210));
INVX1 gate269(.O (I214), .I (n2861gat));
INVX1 gate270(.O (n2860gat), .I (I214));
INVX1 gate271(.O (I217), .I (n2860gat));
INVX1 gate272(.O (n1221gat), .I (I217));
INVX1 gate273(.O (I220), .I (n2864gat));
INVX1 gate274(.O (n2863gat), .I (I220));
INVX1 gate275(.O (I223), .I (n2863gat));
INVX1 gate276(.O (n1222gat), .I (I223));
INVX1 gate277(.O (I227), .I (n2856gat));
INVX1 gate278(.O (n2855gat), .I (I227));
INVX1 gate279(.O (I230), .I (n2855gat));
INVX1 gate280(.O (n1223gat), .I (I230));
INVX1 gate281(.O (n640gat), .I (n1213gat));
INVX1 gate282(.O (I237), .I (n640gat));
INVX1 gate283(.O (n753gat), .I (I237));
INVX1 gate284(.O (I240), .I (n2717gat));
INVX1 gate285(.O (n2716gat), .I (I240));
INVX1 gate286(.O (I243), .I (n3089gat));
INVX1 gate287(.O (n2869gat), .I (I243));
INVX1 gate288(.O (n2867gat), .I (n2869gat));
INVX1 gate289(.O (I248), .I (n2869gat));
INVX1 gate290(.O (n2868gat), .I (I248));
INVX1 gate291(.O (I253), .I (n2906gat));
INVX1 gate292(.O (n754gat), .I (I253));
INVX1 gate293(.O (I256), .I (n2725gat));
INVX1 gate294(.O (n2724gat), .I (I256));
INVX1 gate295(.O (I259), .I (n3086gat));
INVX1 gate296(.O (n2728gat), .I (I259));
INVX1 gate297(.O (n2726gat), .I (n2728gat));
INVX1 gate298(.O (I264), .I (n2728gat));
INVX1 gate299(.O (n2727gat), .I (I264));
INVX1 gate300(.O (n422gat), .I (n2889gat));
INVX1 gate301(.O (I270), .I (n422gat));
INVX1 gate302(.O (n755gat), .I (I270));
INVX1 gate303(.O (n747gat), .I (n2906gat));
INVX1 gate304(.O (I275), .I (n747gat));
INVX1 gate305(.O (n756gat), .I (I275));
INVX1 gate306(.O (I278), .I (n2889gat));
INVX1 gate307(.O (n757gat), .I (I278));
INVX1 gate308(.O (I282), .I (n1213gat));
INVX1 gate309(.O (n758gat), .I (I282));
INVX1 gate310(.O (n2508gat), .I (n2510gat));
INVX1 gate311(.O (I297), .I (n3065gat));
INVX1 gate312(.O (n2733gat), .I (I297));
INVX1 gate313(.O (I300), .I (n2733gat));
INVX1 gate314(.O (n2732gat), .I (I300));
INVX1 gate315(.O (I311), .I (n271gat));
INVX1 gate316(.O (n270gat), .I (I311));
INVX1 gate317(.O (I314), .I (n270gat));
INVX1 gate318(.O (n263gat), .I (I314));
INVX1 gate319(.O (I317), .I (n3067gat));
INVX1 gate320(.O (n2777gat), .I (I317));
INVX1 gate321(.O (I320), .I (n2777gat));
INVX1 gate322(.O (n2776gat), .I (I320));
INVX1 gate323(.O (I331), .I (n160gat));
INVX1 gate324(.O (n159gat), .I (I331));
INVX1 gate325(.O (I334), .I (n159gat));
INVX1 gate326(.O (n264gat), .I (I334));
INVX1 gate327(.O (I337), .I (n3066gat));
INVX1 gate328(.O (n2736gat), .I (I337));
INVX1 gate329(.O (I340), .I (n2736gat));
INVX1 gate330(.O (n2735gat), .I (I340));
INVX1 gate331(.O (I351), .I (n337gat));
INVX1 gate332(.O (n336gat), .I (I351));
INVX1 gate333(.O (I354), .I (n336gat));
INVX1 gate334(.O (n265gat), .I (I354));
INVX1 gate335(.O (n158gat), .I (n160gat));
INVX1 gate336(.O (I359), .I (n158gat));
INVX1 gate337(.O (n266gat), .I (I359));
INVX1 gate338(.O (n335gat), .I (n337gat));
INVX1 gate339(.O (I363), .I (n335gat));
INVX1 gate340(.O (n267gat), .I (I363));
INVX1 gate341(.O (n269gat), .I (n271gat));
INVX1 gate342(.O (I368), .I (n269gat));
INVX1 gate343(.O (n268gat), .I (I368));
INVX1 gate344(.O (n41gat), .I (n258gat));
INVX1 gate345(.O (I375), .I (n41gat));
INVX1 gate346(.O (n48gat), .I (I375));
INVX1 gate347(.O (I378), .I (n725gat));
INVX1 gate348(.O (n1018gat), .I (I378));
INVX1 gate349(.O (I381), .I (n3073gat));
INVX1 gate350(.O (n2674gat), .I (I381));
INVX1 gate351(.O (I384), .I (n2674gat));
INVX1 gate352(.O (n2673gat), .I (I384));
INVX1 gate353(.O (I395), .I (n842gat));
INVX1 gate354(.O (n841gat), .I (I395));
INVX1 gate355(.O (I398), .I (n841gat));
INVX1 gate356(.O (n1019gat), .I (I398));
INVX1 gate357(.O (I401), .I (n721gat));
INVX1 gate358(.O (n1020gat), .I (I401));
INVX1 gate359(.O (n840gat), .I (n842gat));
INVX1 gate360(.O (I406), .I (n840gat));
INVX1 gate361(.O (n1021gat), .I (I406));
INVX1 gate362(.O (I409), .I (n720gat));
INVX1 gate363(.O (n1022gat), .I (I409));
INVX1 gate364(.O (n724gat), .I (n726gat));
INVX1 gate365(.O (I414), .I (n724gat));
INVX1 gate366(.O (n1023gat), .I (I414));
INVX1 gate367(.O (I420), .I (n1013gat));
INVX1 gate368(.O (n49gat), .I (I420));
INVX1 gate369(.O (I423), .I (n3068gat));
INVX1 gate370(.O (n2780gat), .I (I423));
INVX1 gate371(.O (I426), .I (n2780gat));
INVX1 gate372(.O (n2779gat), .I (I426));
INVX1 gate373(.O (I437), .I (n341gat));
INVX1 gate374(.O (n340gat), .I (I437));
INVX1 gate375(.O (I440), .I (n340gat));
INVX1 gate376(.O (n480gat), .I (I440));
INVX1 gate377(.O (I443), .I (n702gat));
INVX1 gate378(.O (n481gat), .I (I443));
INVX1 gate379(.O (I446), .I (n394gat));
INVX1 gate380(.O (n393gat), .I (I446));
INVX1 gate381(.O (I449), .I (n393gat));
INVX1 gate382(.O (n482gat), .I (I449));
INVX1 gate383(.O (I453), .I (n701gat));
INVX1 gate384(.O (n483gat), .I (I453));
INVX1 gate385(.O (I456), .I (n392gat));
INVX1 gate386(.O (n484gat), .I (I456));
INVX1 gate387(.O (n339gat), .I (n341gat));
INVX1 gate388(.O (I461), .I (n339gat));
INVX1 gate389(.O (n485gat), .I (I461));
INVX1 gate390(.O (n42gat), .I (n475gat));
INVX1 gate391(.O (I468), .I (n42gat));
INVX1 gate392(.O (n50gat), .I (I468));
INVX1 gate393(.O (n162gat), .I (n1013gat));
INVX1 gate394(.O (I473), .I (n162gat));
INVX1 gate395(.O (n51gat), .I (I473));
INVX1 gate396(.O (I476), .I (n475gat));
INVX1 gate397(.O (n52gat), .I (I476));
INVX1 gate398(.O (I480), .I (n258gat));
INVX1 gate399(.O (n53gat), .I (I480));
INVX1 gate400(.O (n2520gat), .I (n2522gat));
INVX1 gate401(.O (n1448gat), .I (n1376gat));
INVX1 gate402(.O (n1701gat), .I (n1617gat));
INVX1 gate403(.O (n1379gat), .I (n1377gat));
INVX1 gate404(.O (n1615gat), .I (n1624gat));
INVX1 gate405(.O (n1500gat), .I (n1113gat));
INVX1 gate406(.O (n1503gat), .I (n1501gat));
INVX1 gate407(.O (n1779gat), .I (n1623gat));
INVX1 gate408(.O (I509), .I (n3099gat));
INVX1 gate409(.O (n2730gat), .I (I509));
INVX1 gate410(.O (I512), .I (n2730gat));
INVX1 gate411(.O (n2729gat), .I (I512));
INVX1 gate412(.O (n2470gat), .I (n2472gat));
INVX1 gate413(.O (n2317gat), .I (n2319gat));
INVX1 gate414(.O (n1819gat), .I (n1821gat));
INVX1 gate415(.O (n1823gat), .I (n1825gat));
INVX1 gate416(.O (n1816gat), .I (n1817gat));
INVX1 gate417(.O (n2027gat), .I (n2029gat));
INVX1 gate418(.O (I572), .I (n1829gat));
INVX1 gate419(.O (n1828gat), .I (I572));
INVX1 gate420(.O (I576), .I (n3100gat));
INVX1 gate421(.O (n2851gat), .I (I576));
INVX1 gate422(.O (I579), .I (n2851gat));
INVX1 gate423(.O (n2850gat), .I (I579));
INVX1 gate424(.O (I583), .I (n2786gat));
INVX1 gate425(.O (n2785gat), .I (I583));
INVX1 gate426(.O (n92gat), .I (n2785gat));
INVX1 gate427(.O (n637gat), .I (n529gat));
INVX1 gate428(.O (n293gat), .I (n361gat));
INVX1 gate429(.O (I591), .I (n3094gat));
INVX1 gate430(.O (n2722gat), .I (I591));
INVX1 gate431(.O (I594), .I (n2722gat));
INVX1 gate432(.O (n2721gat), .I (I594));
INVX1 gate433(.O (n297gat), .I (n2721gat));
INVX1 gate434(.O (I606), .I (n283gat));
INVX1 gate435(.O (n282gat), .I (I606));
INVX1 gate436(.O (I609), .I (n282gat));
INVX1 gate437(.O (n172gat), .I (I609));
INVX1 gate438(.O (I620), .I (n165gat));
INVX1 gate439(.O (n164gat), .I (I620));
INVX1 gate440(.O (I623), .I (n164gat));
INVX1 gate441(.O (n173gat), .I (I623));
INVX1 gate442(.O (I634), .I (n279gat));
INVX1 gate443(.O (n278gat), .I (I634));
INVX1 gate444(.O (I637), .I (n278gat));
INVX1 gate445(.O (n174gat), .I (I637));
INVX1 gate446(.O (n163gat), .I (n165gat));
INVX1 gate447(.O (I642), .I (n163gat));
INVX1 gate448(.O (n175gat), .I (I642));
INVX1 gate449(.O (n277gat), .I (n279gat));
INVX1 gate450(.O (I646), .I (n277gat));
INVX1 gate451(.O (n176gat), .I (I646));
INVX1 gate452(.O (n281gat), .I (n283gat));
INVX1 gate453(.O (I651), .I (n281gat));
INVX1 gate454(.O (n177gat), .I (I651));
INVX1 gate455(.O (n54gat), .I (n167gat));
INVX1 gate456(.O (I658), .I (n54gat));
INVX1 gate457(.O (n60gat), .I (I658));
INVX1 gate458(.O (I661), .I (n845gat));
INVX1 gate459(.O (n911gat), .I (I661));
INVX1 gate460(.O (I672), .I (n1026gat));
INVX1 gate461(.O (n1025gat), .I (I672));
INVX1 gate462(.O (I675), .I (n1025gat));
INVX1 gate463(.O (n912gat), .I (I675));
INVX1 gate464(.O (I678), .I (n918gat));
INVX1 gate465(.O (n913gat), .I (I678));
INVX1 gate466(.O (n1024gat), .I (n1026gat));
INVX1 gate467(.O (I683), .I (n1024gat));
INVX1 gate468(.O (n914gat), .I (I683));
INVX1 gate469(.O (n917gat), .I (n919gat));
INVX1 gate470(.O (I687), .I (n917gat));
INVX1 gate471(.O (n915gat), .I (I687));
INVX1 gate472(.O (n844gat), .I (n846gat));
INVX1 gate473(.O (I692), .I (n844gat));
INVX1 gate474(.O (n916gat), .I (I692));
INVX1 gate475(.O (I698), .I (n906gat));
INVX1 gate476(.O (n61gat), .I (I698));
INVX1 gate477(.O (I709), .I (n275gat));
INVX1 gate478(.O (n274gat), .I (I709));
INVX1 gate479(.O (I712), .I (n274gat));
INVX1 gate480(.O (n348gat), .I (I712));
INVX1 gate481(.O (I715), .I (n401gat));
INVX1 gate482(.O (n349gat), .I (I715));
INVX1 gate483(.O (I718), .I (n398gat));
INVX1 gate484(.O (n397gat), .I (I718));
INVX1 gate485(.O (I721), .I (n397gat));
INVX1 gate486(.O (n350gat), .I (I721));
INVX1 gate487(.O (n400gat), .I (n402gat));
INVX1 gate488(.O (I726), .I (n400gat));
INVX1 gate489(.O (n351gat), .I (I726));
INVX1 gate490(.O (I729), .I (n396gat));
INVX1 gate491(.O (n352gat), .I (I729));
INVX1 gate492(.O (n273gat), .I (n275gat));
INVX1 gate493(.O (I734), .I (n273gat));
INVX1 gate494(.O (n353gat), .I (I734));
INVX1 gate495(.O (n178gat), .I (n343gat));
INVX1 gate496(.O (I741), .I (n178gat));
INVX1 gate497(.O (n62gat), .I (I741));
INVX1 gate498(.O (n66gat), .I (n906gat));
INVX1 gate499(.O (I746), .I (n66gat));
INVX1 gate500(.O (n63gat), .I (I746));
INVX1 gate501(.O (I749), .I (n343gat));
INVX1 gate502(.O (n64gat), .I (I749));
INVX1 gate503(.O (I753), .I (n167gat));
INVX1 gate504(.O (n65gat), .I (I753));
INVX1 gate505(.O (n2474gat), .I (n2476gat));
INVX1 gate506(.O (I768), .I (n3090gat));
INVX1 gate507(.O (n2832gat), .I (I768));
INVX1 gate508(.O (I771), .I (n2832gat));
INVX1 gate509(.O (n2831gat), .I (I771));
INVX1 gate510(.O (n2731gat), .I (n2733gat));
INVX1 gate511(.O (I776), .I (n3074gat));
INVX1 gate512(.O (n2719gat), .I (I776));
INVX1 gate513(.O (n2718gat), .I (n2719gat));
INVX1 gate514(.O (I790), .I (n1068gat));
INVX1 gate515(.O (n1067gat), .I (I790));
INVX1 gate516(.O (I793), .I (n1067gat));
INVX1 gate517(.O (n949gat), .I (I793));
INVX1 gate518(.O (I796), .I (n3076gat));
INVX1 gate519(.O (n2839gat), .I (I796));
INVX1 gate520(.O (n2838gat), .I (n2839gat));
INVX1 gate521(.O (n2775gat), .I (n2777gat));
INVX1 gate522(.O (I812), .I (n957gat));
INVX1 gate523(.O (n956gat), .I (I812));
INVX1 gate524(.O (I815), .I (n956gat));
INVX1 gate525(.O (n950gat), .I (I815));
INVX1 gate526(.O (I818), .I (n3075gat));
INVX1 gate527(.O (n2712gat), .I (I818));
INVX1 gate528(.O (n2711gat), .I (n2712gat));
INVX1 gate529(.O (n2734gat), .I (n2736gat));
INVX1 gate530(.O (I834), .I (n861gat));
INVX1 gate531(.O (n860gat), .I (I834));
INVX1 gate532(.O (I837), .I (n860gat));
INVX1 gate533(.O (n951gat), .I (I837));
INVX1 gate534(.O (n955gat), .I (n957gat));
INVX1 gate535(.O (I842), .I (n955gat));
INVX1 gate536(.O (n952gat), .I (I842));
INVX1 gate537(.O (n859gat), .I (n861gat));
INVX1 gate538(.O (I846), .I (n859gat));
INVX1 gate539(.O (n953gat), .I (I846));
INVX1 gate540(.O (n1066gat), .I (n1068gat));
INVX1 gate541(.O (I851), .I (n1066gat));
INVX1 gate542(.O (n954gat), .I (I851));
INVX1 gate543(.O (n857gat), .I (n944gat));
INVX1 gate544(.O (I858), .I (n857gat));
INVX1 gate545(.O (n938gat), .I (I858));
INVX1 gate546(.O (n2792gat), .I (n2794gat));
INVX1 gate547(.O (I863), .I (n3080gat));
INVX1 gate548(.O (n2847gat), .I (I863));
INVX1 gate549(.O (n2846gat), .I (n2847gat));
INVX1 gate550(.O (I877), .I (n1294gat));
INVX1 gate551(.O (n1293gat), .I (I877));
INVX1 gate552(.O (I880), .I (n1293gat));
INVX1 gate553(.O (n1233gat), .I (I880));
INVX1 gate554(.O (n2672gat), .I (n2674gat));
INVX1 gate555(.O (I885), .I (n3082gat));
INVX1 gate556(.O (n2853gat), .I (I885));
INVX1 gate557(.O (n2852gat), .I (n2853gat));
INVX1 gate558(.O (I899), .I (n1241gat));
INVX1 gate559(.O (n1240gat), .I (I899));
INVX1 gate560(.O (I902), .I (n1240gat));
INVX1 gate561(.O (n1234gat), .I (I902));
INVX1 gate562(.O (I913), .I (n1298gat));
INVX1 gate563(.O (n1297gat), .I (I913));
INVX1 gate564(.O (I916), .I (n1297gat));
INVX1 gate565(.O (n1235gat), .I (I916));
INVX1 gate566(.O (n1239gat), .I (n1241gat));
INVX1 gate567(.O (I921), .I (n1239gat));
INVX1 gate568(.O (n1236gat), .I (I921));
INVX1 gate569(.O (n1296gat), .I (n1298gat));
INVX1 gate570(.O (I925), .I (n1296gat));
INVX1 gate571(.O (n1237gat), .I (I925));
INVX1 gate572(.O (n1292gat), .I (n1294gat));
INVX1 gate573(.O (I930), .I (n1292gat));
INVX1 gate574(.O (n1238gat), .I (I930));
INVX1 gate575(.O (I936), .I (n1228gat));
INVX1 gate576(.O (n939gat), .I (I936));
INVX1 gate577(.O (n2778gat), .I (n2780gat));
INVX1 gate578(.O (I941), .I (n3077gat));
INVX1 gate579(.O (n2837gat), .I (I941));
INVX1 gate580(.O (n2836gat), .I (n2837gat));
INVX1 gate581(.O (I955), .I (n865gat));
INVX1 gate582(.O (n864gat), .I (I955));
INVX1 gate583(.O (I958), .I (n864gat));
INVX1 gate584(.O (n1055gat), .I (I958));
INVX1 gate585(.O (n2789gat), .I (n2791gat));
INVX1 gate586(.O (I963), .I (n3079gat));
INVX1 gate587(.O (n2841gat), .I (I963));
INVX1 gate588(.O (n2840gat), .I (n2841gat));
INVX1 gate589(.O (I977), .I (n1080gat));
INVX1 gate590(.O (n1079gat), .I (I977));
INVX1 gate591(.O (I980), .I (n1079gat));
INVX1 gate592(.O (n1056gat), .I (I980));
INVX1 gate593(.O (n2781gat), .I (n2783gat));
INVX1 gate594(.O (I985), .I (n3078gat));
INVX1 gate595(.O (n2843gat), .I (I985));
INVX1 gate596(.O (n2842gat), .I (n2843gat));
INVX1 gate597(.O (I999), .I (n1148gat));
INVX1 gate598(.O (n1147gat), .I (I999));
INVX1 gate599(.O (I1002), .I (n1147gat));
INVX1 gate600(.O (n1057gat), .I (I1002));
INVX1 gate601(.O (n1078gat), .I (n1080gat));
INVX1 gate602(.O (I1007), .I (n1078gat));
INVX1 gate603(.O (n1058gat), .I (I1007));
INVX1 gate604(.O (n1146gat), .I (n1148gat));
INVX1 gate605(.O (I1011), .I (n1146gat));
INVX1 gate606(.O (n1059gat), .I (I1011));
INVX1 gate607(.O (n863gat), .I (n865gat));
INVX1 gate608(.O (I1016), .I (n863gat));
INVX1 gate609(.O (n1060gat), .I (I1016));
INVX1 gate610(.O (n928gat), .I (n1050gat));
INVX1 gate611(.O (I1023), .I (n928gat));
INVX1 gate612(.O (n940gat), .I (I1023));
INVX1 gate613(.O (n858gat), .I (n1228gat));
INVX1 gate614(.O (I1028), .I (n858gat));
INVX1 gate615(.O (n941gat), .I (I1028));
INVX1 gate616(.O (I1031), .I (n1050gat));
INVX1 gate617(.O (n942gat), .I (I1031));
INVX1 gate618(.O (I1035), .I (n944gat));
INVX1 gate619(.O (n943gat), .I (I1035));
INVX1 gate620(.O (n2466gat), .I (n2468gat));
INVX1 gate621(.O (n2720gat), .I (n2722gat));
INVX1 gate622(.O (n740gat), .I (n2667gat));
INVX1 gate623(.O (n2784gat), .I (n2786gat));
INVX1 gate624(.O (n743gat), .I (n746gat));
INVX1 gate625(.O (n294gat), .I (n360gat));
INVX1 gate626(.O (n374gat), .I (n2767gat));
INVX1 gate627(.O (n616gat), .I (n618gat));
INVX1 gate628(.O (I1067), .I (n616gat));
INVX1 gate629(.O (n501gat), .I (I1067));
INVX1 gate630(.O (n489gat), .I (n491gat));
INVX1 gate631(.O (I1079), .I (n489gat));
INVX1 gate632(.O (n502gat), .I (I1079));
INVX1 gate633(.O (I1082), .I (n618gat));
INVX1 gate634(.O (n617gat), .I (I1082));
INVX1 gate635(.O (I1085), .I (n617gat));
INVX1 gate636(.O (n499gat), .I (I1085));
INVX1 gate637(.O (I1088), .I (n491gat));
INVX1 gate638(.O (n490gat), .I (I1088));
INVX1 gate639(.O (I1091), .I (n490gat));
INVX1 gate640(.O (n500gat), .I (I1091));
INVX1 gate641(.O (n620gat), .I (n622gat));
INVX1 gate642(.O (I1103), .I (n620gat));
INVX1 gate643(.O (n738gat), .I (I1103));
INVX1 gate644(.O (n624gat), .I (n626gat));
INVX1 gate645(.O (I1115), .I (n624gat));
INVX1 gate646(.O (n737gat), .I (I1115));
INVX1 gate647(.O (I1118), .I (n622gat));
INVX1 gate648(.O (n621gat), .I (I1118));
INVX1 gate649(.O (I1121), .I (n621gat));
INVX1 gate650(.O (n733gat), .I (I1121));
INVX1 gate651(.O (I1124), .I (n626gat));
INVX1 gate652(.O (n625gat), .I (I1124));
INVX1 gate653(.O (I1127), .I (n625gat));
INVX1 gate654(.O (n735gat), .I (I1127));
INVX1 gate655(.O (I1138), .I (n834gat));
INVX1 gate656(.O (n833gat), .I (I1138));
INVX1 gate657(.O (I1141), .I (n833gat));
INVX1 gate658(.O (n714gat), .I (I1141));
INVX1 gate659(.O (I1152), .I (n707gat));
INVX1 gate660(.O (n706gat), .I (I1152));
INVX1 gate661(.O (I1155), .I (n706gat));
INVX1 gate662(.O (n715gat), .I (I1155));
INVX1 gate663(.O (I1166), .I (n838gat));
INVX1 gate664(.O (n837gat), .I (I1166));
INVX1 gate665(.O (I1169), .I (n837gat));
INVX1 gate666(.O (n716gat), .I (I1169));
INVX1 gate667(.O (n705gat), .I (n707gat));
INVX1 gate668(.O (I1174), .I (n705gat));
INVX1 gate669(.O (n717gat), .I (I1174));
INVX1 gate670(.O (n836gat), .I (n838gat));
INVX1 gate671(.O (I1178), .I (n836gat));
INVX1 gate672(.O (n718gat), .I (I1178));
INVX1 gate673(.O (n832gat), .I (n834gat));
INVX1 gate674(.O (I1183), .I (n832gat));
INVX1 gate675(.O (n719gat), .I (I1183));
INVX1 gate676(.O (n515gat), .I (n709gat));
INVX1 gate677(.O (I1190), .I (n515gat));
INVX1 gate678(.O (n509gat), .I (I1190));
INVX1 gate679(.O (I1201), .I (n830gat));
INVX1 gate680(.O (n829gat), .I (I1201));
INVX1 gate681(.O (I1204), .I (n829gat));
INVX1 gate682(.O (n734gat), .I (I1204));
INVX1 gate683(.O (n828gat), .I (n830gat));
INVX1 gate684(.O (I1209), .I (n828gat));
INVX1 gate685(.O (n736gat), .I (I1209));
INVX1 gate686(.O (I1216), .I (n728gat));
INVX1 gate687(.O (n510gat), .I (I1216));
INVX1 gate688(.O (I1227), .I (n614gat));
INVX1 gate689(.O (n613gat), .I (I1227));
INVX1 gate690(.O (I1230), .I (n613gat));
INVX1 gate691(.O (n498gat), .I (I1230));
INVX1 gate692(.O (n612gat), .I (n614gat));
INVX1 gate693(.O (I1236), .I (n612gat));
INVX1 gate694(.O (n503gat), .I (I1236));
INVX1 gate695(.O (n404gat), .I (n493gat));
INVX1 gate696(.O (I1243), .I (n404gat));
INVX1 gate697(.O (n511gat), .I (I1243));
INVX1 gate698(.O (n405gat), .I (n728gat));
INVX1 gate699(.O (I1248), .I (n405gat));
INVX1 gate700(.O (n512gat), .I (I1248));
INVX1 gate701(.O (I1251), .I (n493gat));
INVX1 gate702(.O (n513gat), .I (I1251));
INVX1 gate703(.O (I1255), .I (n709gat));
INVX1 gate704(.O (n514gat), .I (I1255));
INVX1 gate705(.O (n2524gat), .I (n2526gat));
INVX1 gate706(.O (n17gat), .I (n564gat));
INVX1 gate707(.O (n79gat), .I (n86gat));
INVX1 gate708(.O (n219gat), .I (n78gat));
INVX1 gate709(.O (n563gat), .I (I1278));
INVX1 gate710(.O (n289gat), .I (n563gat));
INVX1 gate711(.O (n179gat), .I (n287gat));
INVX1 gate712(.O (n188gat), .I (n288gat));
INVX1 gate713(.O (n72gat), .I (n181gat));
INVX1 gate714(.O (n111gat), .I (n182gat));
INVX1 gate715(.O (I1302), .I (n680gat));
INVX1 gate716(.O (n679gat), .I (I1302));
INVX1 gate717(.O (I1305), .I (n679gat));
INVX1 gate718(.O (n808gat), .I (I1305));
INVX1 gate719(.O (I1319), .I (n816gat));
INVX1 gate720(.O (n815gat), .I (I1319));
INVX1 gate721(.O (I1322), .I (n815gat));
INVX1 gate722(.O (n809gat), .I (I1322));
INVX1 gate723(.O (I1336), .I (n580gat));
INVX1 gate724(.O (n579gat), .I (I1336));
INVX1 gate725(.O (I1339), .I (n579gat));
INVX1 gate726(.O (n810gat), .I (I1339));
INVX1 gate727(.O (n814gat), .I (n816gat));
INVX1 gate728(.O (I1344), .I (n814gat));
INVX1 gate729(.O (n811gat), .I (I1344));
INVX1 gate730(.O (n578gat), .I (n580gat));
INVX1 gate731(.O (I1348), .I (n578gat));
INVX1 gate732(.O (n812gat), .I (I1348));
INVX1 gate733(.O (n678gat), .I (n680gat));
INVX1 gate734(.O (I1353), .I (n678gat));
INVX1 gate735(.O (n813gat), .I (I1353));
INVX1 gate736(.O (n677gat), .I (n803gat));
INVX1 gate737(.O (I1360), .I (n677gat));
INVX1 gate738(.O (n572gat), .I (I1360));
INVX1 gate739(.O (I1371), .I (n824gat));
INVX1 gate740(.O (n823gat), .I (I1371));
INVX1 gate741(.O (I1374), .I (n823gat));
INVX1 gate742(.O (n591gat), .I (I1374));
INVX1 gate743(.O (I1385), .I (n820gat));
INVX1 gate744(.O (n819gat), .I (I1385));
INVX1 gate745(.O (I1388), .I (n819gat));
INVX1 gate746(.O (n592gat), .I (I1388));
INVX1 gate747(.O (I1399), .I (n883gat));
INVX1 gate748(.O (n882gat), .I (I1399));
INVX1 gate749(.O (I1402), .I (n882gat));
INVX1 gate750(.O (n593gat), .I (I1402));
INVX1 gate751(.O (n818gat), .I (n820gat));
INVX1 gate752(.O (I1407), .I (n818gat));
INVX1 gate753(.O (n594gat), .I (I1407));
INVX1 gate754(.O (n881gat), .I (n883gat));
INVX1 gate755(.O (I1411), .I (n881gat));
INVX1 gate756(.O (n595gat), .I (I1411));
INVX1 gate757(.O (n822gat), .I (n824gat));
INVX1 gate758(.O (I1416), .I (n822gat));
INVX1 gate759(.O (n596gat), .I (I1416));
INVX1 gate760(.O (I1422), .I (n586gat));
INVX1 gate761(.O (n573gat), .I (I1422));
INVX1 gate762(.O (I1436), .I (n584gat));
INVX1 gate763(.O (n583gat), .I (I1436));
INVX1 gate764(.O (I1439), .I (n583gat));
INVX1 gate765(.O (n691gat), .I (I1439));
INVX1 gate766(.O (I1450), .I (n684gat));
INVX1 gate767(.O (n683gat), .I (I1450));
INVX1 gate768(.O (I1453), .I (n683gat));
INVX1 gate769(.O (n692gat), .I (I1453));
INVX1 gate770(.O (I1464), .I (n699gat));
INVX1 gate771(.O (n698gat), .I (I1464));
INVX1 gate772(.O (I1467), .I (n698gat));
INVX1 gate773(.O (n693gat), .I (I1467));
INVX1 gate774(.O (n682gat), .I (n684gat));
INVX1 gate775(.O (I1472), .I (n682gat));
INVX1 gate776(.O (n694gat), .I (I1472));
INVX1 gate777(.O (n697gat), .I (n699gat));
INVX1 gate778(.O (I1476), .I (n697gat));
INVX1 gate779(.O (n695gat), .I (I1476));
INVX1 gate780(.O (n582gat), .I (n584gat));
INVX1 gate781(.O (I1481), .I (n582gat));
INVX1 gate782(.O (n696gat), .I (I1481));
INVX1 gate783(.O (n456gat), .I (n686gat));
INVX1 gate784(.O (I1488), .I (n456gat));
INVX1 gate785(.O (n574gat), .I (I1488));
INVX1 gate786(.O (n565gat), .I (n586gat));
INVX1 gate787(.O (I1493), .I (n565gat));
INVX1 gate788(.O (n575gat), .I (I1493));
INVX1 gate789(.O (I1496), .I (n686gat));
INVX1 gate790(.O (n576gat), .I (I1496));
INVX1 gate791(.O (I1500), .I (n803gat));
INVX1 gate792(.O (n577gat), .I (I1500));
INVX1 gate793(.O (n2462gat), .I (n2464gat));
INVX1 gate794(.O (n2665gat), .I (I1516));
INVX1 gate795(.O (n2596gat), .I (n2665gat));
INVX1 gate796(.O (n189gat), .I (n286gat));
INVX1 gate797(.O (n194gat), .I (n187gat));
INVX1 gate798(.O (n21gat), .I (n15gat));
INVX1 gate799(.O (I1538), .I (n2399gat));
INVX1 gate800(.O (n2398gat), .I (I1538));
INVX1 gate801(.O (n2353gat), .I (n2398gat));
INVX1 gate802(.O (I1550), .I (n2343gat));
INVX1 gate803(.O (n2342gat), .I (I1550));
INVX1 gate804(.O (n2284gat), .I (n2342gat));
INVX1 gate805(.O (n2201gat), .I (n2203gat));
INVX1 gate806(.O (n2354gat), .I (n2201gat));
INVX1 gate807(.O (n2560gat), .I (n2562gat));
INVX1 gate808(.O (n2356gat), .I (n2560gat));
INVX1 gate809(.O (n2205gat), .I (n2207gat));
INVX1 gate810(.O (n2214gat), .I (n2205gat));
INVX1 gate811(.O (n2286gat), .I (I1585));
INVX1 gate812(.O (n2624gat), .I (n2626gat));
INVX1 gate813(.O (I1606), .I (n2490gat));
INVX1 gate814(.O (n2489gat), .I (I1606));
INVX1 gate815(.O (I1617), .I (n2622gat));
INVX1 gate816(.O (n2621gat), .I (I1617));
INVX1 gate817(.O (n2533gat), .I (n2534gat));
INVX1 gate818(.O (I1630), .I (n2630gat));
INVX1 gate819(.O (n2629gat), .I (I1630));
INVX1 gate820(.O (n2486gat), .I (n2629gat));
INVX1 gate821(.O (n2541gat), .I (n2543gat));
INVX1 gate822(.O (n2429gat), .I (n2541gat));
INVX1 gate823(.O (n2432gat), .I (n2430gat));
INVX1 gate824(.O (I1655), .I (n2102gat));
INVX1 gate825(.O (n2101gat), .I (I1655));
INVX1 gate826(.O (n1693gat), .I (n2101gat));
INVX1 gate827(.O (I1667), .I (n1880gat));
INVX1 gate828(.O (n1879gat), .I (I1667));
INVX1 gate829(.O (n1698gat), .I (n1934gat));
INVX1 gate830(.O (n1543gat), .I (n1606gat));
INVX1 gate831(.O (I1683), .I (n1763gat));
INVX1 gate832(.O (n1762gat), .I (I1683));
INVX1 gate833(.O (n1673gat), .I (n2989gat));
INVX1 gate834(.O (n1858gat), .I (n1673gat));
INVX1 gate835(.O (I1698), .I (n2155gat));
INVX1 gate836(.O (n2154gat), .I (I1698));
INVX1 gate837(.O (n2488gat), .I (n2490gat));
INVX1 gate838(.O (I1703), .I (n2626gat));
INVX1 gate839(.O (n2625gat), .I (I1703));
INVX1 gate840(.O (n2530gat), .I (n2531gat));
INVX1 gate841(.O (I1708), .I (n2543gat));
INVX1 gate842(.O (n2542gat), .I (I1708));
INVX1 gate843(.O (n2482gat), .I (n2542gat));
INVX1 gate844(.O (n2426gat), .I (n2480gat));
INVX1 gate845(.O (n2153gat), .I (n2155gat));
INVX1 gate846(.O (n2341gat), .I (n2343gat));
INVX1 gate847(.O (n2355gat), .I (n2341gat));
INVX1 gate848(.O (I1719), .I (n2562gat));
INVX1 gate849(.O (n2561gat), .I (I1719));
INVX1 gate850(.O (n2443gat), .I (n2561gat));
INVX1 gate851(.O (n2289gat), .I (I1724));
INVX1 gate852(.O (n2148gat), .I (I1734));
INVX1 gate853(.O (n855gat), .I (n2148gat));
INVX1 gate854(.O (n759gat), .I (n855gat));
INVX1 gate855(.O (I1749), .I (n1035gat));
INVX1 gate856(.O (n1034gat), .I (I1749));
INVX1 gate857(.O (I1752), .I (n1034gat));
INVX1 gate858(.O (n1189gat), .I (I1752));
INVX1 gate859(.O (n1075gat), .I (n855gat));
INVX1 gate860(.O (I1766), .I (n1121gat));
INVX1 gate861(.O (n1120gat), .I (I1766));
INVX1 gate862(.O (I1769), .I (n1120gat));
INVX1 gate863(.O (n1190gat), .I (I1769));
INVX1 gate864(.O (n760gat), .I (n855gat));
INVX1 gate865(.O (I1783), .I (n1072gat));
INVX1 gate866(.O (n1071gat), .I (I1783));
INVX1 gate867(.O (I1786), .I (n1071gat));
INVX1 gate868(.O (n1191gat), .I (I1786));
INVX1 gate869(.O (n1119gat), .I (n1121gat));
INVX1 gate870(.O (I1791), .I (n1119gat));
INVX1 gate871(.O (n1192gat), .I (I1791));
INVX1 gate872(.O (n1070gat), .I (n1072gat));
INVX1 gate873(.O (I1795), .I (n1070gat));
INVX1 gate874(.O (n1193gat), .I (I1795));
INVX1 gate875(.O (n1033gat), .I (n1035gat));
INVX1 gate876(.O (I1800), .I (n1033gat));
INVX1 gate877(.O (n1194gat), .I (I1800));
INVX1 gate878(.O (n1183gat), .I (n1184gat));
INVX1 gate879(.O (I1807), .I (n1183gat));
INVX1 gate880(.O (n1274gat), .I (I1807));
INVX1 gate881(.O (n644gat), .I (n855gat));
INVX1 gate882(.O (n1280gat), .I (n1282gat));
INVX1 gate883(.O (n641gat), .I (n855gat));
INVX1 gate884(.O (I1833), .I (n1226gat));
INVX1 gate885(.O (n1225gat), .I (I1833));
INVX1 gate886(.O (I1837), .I (n1282gat));
INVX1 gate887(.O (n1281gat), .I (I1837));
INVX1 gate888(.O (n1224gat), .I (n1226gat));
INVX1 gate889(.O (I1843), .I (n2970gat));
INVX1 gate890(.O (n1275gat), .I (I1843));
INVX1 gate891(.O (n761gat), .I (n855gat));
INVX1 gate892(.O (I1857), .I (n931gat));
INVX1 gate893(.O (n930gat), .I (I1857));
INVX1 gate894(.O (I1860), .I (n930gat));
INVX1 gate895(.O (n1206gat), .I (I1860));
INVX1 gate896(.O (n762gat), .I (n855gat));
INVX1 gate897(.O (I1874), .I (n1135gat));
INVX1 gate898(.O (n1134gat), .I (I1874));
INVX1 gate899(.O (I1877), .I (n1134gat));
INVX1 gate900(.O (n1207gat), .I (I1877));
INVX1 gate901(.O (n643gat), .I (n855gat));
INVX1 gate902(.O (I1891), .I (n1045gat));
INVX1 gate903(.O (n1044gat), .I (I1891));
INVX1 gate904(.O (I1894), .I (n1044gat));
INVX1 gate905(.O (n1208gat), .I (I1894));
INVX1 gate906(.O (n1133gat), .I (n1135gat));
INVX1 gate907(.O (I1899), .I (n1133gat));
INVX1 gate908(.O (n1209gat), .I (I1899));
INVX1 gate909(.O (n1043gat), .I (n1045gat));
INVX1 gate910(.O (I1903), .I (n1043gat));
INVX1 gate911(.O (n1210gat), .I (I1903));
INVX1 gate912(.O (n929gat), .I (n931gat));
INVX1 gate913(.O (I1908), .I (n929gat));
INVX1 gate914(.O (n1211gat), .I (I1908));
INVX1 gate915(.O (n1268gat), .I (n1201gat));
INVX1 gate916(.O (I1915), .I (n1268gat));
INVX1 gate917(.O (n1276gat), .I (I1915));
INVX1 gate918(.O (n1329gat), .I (n2970gat));
INVX1 gate919(.O (I1920), .I (n1329gat));
INVX1 gate920(.O (n1277gat), .I (I1920));
INVX1 gate921(.O (I1923), .I (n1201gat));
INVX1 gate922(.O (n1278gat), .I (I1923));
INVX1 gate923(.O (I1927), .I (n1184gat));
INVX1 gate924(.O (n1279gat), .I (I1927));
INVX1 gate925(.O (n1284gat), .I (n1269gat));
INVX1 gate926(.O (n642gat), .I (n855gat));
INVX1 gate927(.O (n1195gat), .I (n1197gat));
INVX1 gate928(.O (I1947), .I (n1197gat));
INVX1 gate929(.O (n1196gat), .I (I1947));
INVX1 gate930(.O (n2516gat), .I (n2518gat));
INVX1 gate931(.O (I1961), .I (n2516gat));
INVX1 gate932(.O (n3017gat), .I (I1961));
INVX1 gate933(.O (n851gat), .I (n853gat));
INVX1 gate934(.O (n1725gat), .I (n2148gat));
INVX1 gate935(.O (n664gat), .I (n1725gat));
INVX1 gate936(.O (n852gat), .I (n854gat));
INVX1 gate937(.O (I1981), .I (n667gat));
INVX1 gate938(.O (n666gat), .I (I1981));
INVX1 gate939(.O (n368gat), .I (n1725gat));
INVX1 gate940(.O (I1996), .I (n659gat));
INVX1 gate941(.O (n658gat), .I (I1996));
INVX1 gate942(.O (I1999), .I (n658gat));
INVX1 gate943(.O (n784gat), .I (I1999));
INVX1 gate944(.O (n662gat), .I (n1725gat));
INVX1 gate945(.O (I2014), .I (n553gat));
INVX1 gate946(.O (n552gat), .I (I2014));
INVX1 gate947(.O (I2017), .I (n552gat));
INVX1 gate948(.O (n785gat), .I (I2017));
INVX1 gate949(.O (n661gat), .I (n1725gat));
INVX1 gate950(.O (I2032), .I (n777gat));
INVX1 gate951(.O (n776gat), .I (I2032));
INVX1 gate952(.O (I2035), .I (n776gat));
INVX1 gate953(.O (n786gat), .I (I2035));
INVX1 gate954(.O (n551gat), .I (n553gat));
INVX1 gate955(.O (I2040), .I (n551gat));
INVX1 gate956(.O (n787gat), .I (I2040));
INVX1 gate957(.O (n775gat), .I (n777gat));
INVX1 gate958(.O (I2044), .I (n775gat));
INVX1 gate959(.O (n788gat), .I (I2044));
INVX1 gate960(.O (n657gat), .I (n659gat));
INVX1 gate961(.O (I2049), .I (n657gat));
INVX1 gate962(.O (n789gat), .I (I2049));
INVX1 gate963(.O (n35gat), .I (n779gat));
INVX1 gate964(.O (I2056), .I (n35gat));
INVX1 gate965(.O (n125gat), .I (I2056));
INVX1 gate966(.O (n558gat), .I (n1725gat));
INVX1 gate967(.O (n559gat), .I (n561gat));
INVX1 gate968(.O (n371gat), .I (n1725gat));
INVX1 gate969(.O (I2084), .I (n366gat));
INVX1 gate970(.O (n365gat), .I (I2084));
INVX1 gate971(.O (I2088), .I (n561gat));
INVX1 gate972(.O (n560gat), .I (I2088));
INVX1 gate973(.O (n364gat), .I (n366gat));
INVX1 gate974(.O (I2094), .I (n2876gat));
INVX1 gate975(.O (n126gat), .I (I2094));
INVX1 gate976(.O (n663gat), .I (n1725gat));
INVX1 gate977(.O (I2109), .I (n322gat));
INVX1 gate978(.O (n321gat), .I (I2109));
INVX1 gate979(.O (I2112), .I (n321gat));
INVX1 gate980(.O (n226gat), .I (I2112));
INVX1 gate981(.O (n370gat), .I (n1725gat));
INVX1 gate982(.O (I2127), .I (n318gat));
INVX1 gate983(.O (n317gat), .I (I2127));
INVX1 gate984(.O (I2130), .I (n317gat));
INVX1 gate985(.O (n227gat), .I (I2130));
INVX1 gate986(.O (n369gat), .I (n1725gat));
INVX1 gate987(.O (I2145), .I (n314gat));
INVX1 gate988(.O (n313gat), .I (I2145));
INVX1 gate989(.O (I2148), .I (n313gat));
INVX1 gate990(.O (n228gat), .I (I2148));
INVX1 gate991(.O (n316gat), .I (n318gat));
INVX1 gate992(.O (I2153), .I (n316gat));
INVX1 gate993(.O (n229gat), .I (I2153));
INVX1 gate994(.O (n312gat), .I (n314gat));
INVX1 gate995(.O (I2157), .I (n312gat));
INVX1 gate996(.O (n230gat), .I (I2157));
INVX1 gate997(.O (n320gat), .I (n322gat));
INVX1 gate998(.O (I2162), .I (n320gat));
INVX1 gate999(.O (n231gat), .I (I2162));
INVX1 gate1000(.O (n34gat), .I (n221gat));
INVX1 gate1001(.O (I2169), .I (n34gat));
INVX1 gate1002(.O (n127gat), .I (I2169));
INVX1 gate1003(.O (n133gat), .I (n2876gat));
INVX1 gate1004(.O (I2174), .I (n133gat));
INVX1 gate1005(.O (n128gat), .I (I2174));
INVX1 gate1006(.O (I2177), .I (n221gat));
INVX1 gate1007(.O (n129gat), .I (I2177));
INVX1 gate1008(.O (I2181), .I (n779gat));
INVX1 gate1009(.O (n130gat), .I (I2181));
INVX1 gate1010(.O (n665gat), .I (n667gat));
INVX1 gate1011(.O (n1601gat), .I (n120gat));
INVX1 gate1012(.O (n2597gat), .I (n2599gat));
INVX1 gate1013(.O (n2595gat), .I (n2594gat));
INVX1 gate1014(.O (n2586gat), .I (n2588gat));
INVX1 gate1015(.O (I2213), .I (n2342gat));
INVX1 gate1016(.O (n2573gat), .I (I2213));
INVX1 gate1017(.O (n2638gat), .I (n2640gat));
INVX1 gate1018(.O (I2225), .I (n2638gat));
INVX1 gate1019(.O (n2574gat), .I (I2225));
INVX1 gate1020(.O (I2228), .I (n2561gat));
INVX1 gate1021(.O (n2575gat), .I (I2228));
INVX1 gate1022(.O (I2232), .I (n2640gat));
INVX1 gate1023(.O (n2639gat), .I (I2232));
INVX1 gate1024(.O (I2235), .I (n2639gat));
INVX1 gate1025(.O (n2576gat), .I (I2235));
INVX1 gate1026(.O (I2238), .I (n2560gat));
INVX1 gate1027(.O (n2577gat), .I (I2238));
INVX1 gate1028(.O (I2242), .I (n2341gat));
INVX1 gate1029(.O (n2578gat), .I (I2242));
INVX1 gate1030(.O (I2248), .I (n2568gat));
INVX1 gate1031(.O (n2582gat), .I (I2248));
INVX1 gate1032(.O (I2251), .I (n2207gat));
INVX1 gate1033(.O (n2206gat), .I (I2251));
INVX1 gate1034(.O (I2254), .I (n2206gat));
INVX1 gate1035(.O (n2414gat), .I (I2254));
INVX1 gate1036(.O (I2257), .I (n2398gat));
INVX1 gate1037(.O (n2415gat), .I (I2257));
INVX1 gate1038(.O (I2260), .I (n2203gat));
INVX1 gate1039(.O (n2202gat), .I (I2260));
INVX1 gate1040(.O (I2263), .I (n2202gat));
INVX1 gate1041(.O (n2416gat), .I (I2263));
INVX1 gate1042(.O (n2397gat), .I (n2399gat));
INVX1 gate1043(.O (I2268), .I (n2397gat));
INVX1 gate1044(.O (n2417gat), .I (I2268));
INVX1 gate1045(.O (I2271), .I (n2201gat));
INVX1 gate1046(.O (n2418gat), .I (I2271));
INVX1 gate1047(.O (I2275), .I (n2205gat));
INVX1 gate1048(.O (n2419gat), .I (I2275));
INVX1 gate1049(.O (I2281), .I (n2409gat));
INVX1 gate1050(.O (n2585gat), .I (I2281));
INVX1 gate1051(.O (n2656gat), .I (n2658gat));
INVX1 gate1052(.O (n2493gat), .I (n2495gat));
INVX1 gate1053(.O (n2388gat), .I (n2390gat));
INVX1 gate1054(.O (I2316), .I (n2390gat));
INVX1 gate1055(.O (n2389gat), .I (I2316));
INVX1 gate1056(.O (I2319), .I (n2495gat));
INVX1 gate1057(.O (n2494gat), .I (I2319));
INVX1 gate1058(.O (I2324), .I (n3014gat));
INVX1 gate1059(.O (n2649gat), .I (I2324));
INVX1 gate1060(.O (n2268gat), .I (n2270gat));
INVX1 gate1061(.O (I2344), .I (n2339gat));
INVX1 gate1062(.O (n2338gat), .I (I2344));
INVX1 gate1063(.O (n2337gat), .I (n2339gat));
INVX1 gate1064(.O (I2349), .I (n2270gat));
INVX1 gate1065(.O (n2269gat), .I (I2349));
INVX1 gate1066(.O (I2354), .I (n2880gat));
INVX1 gate1067(.O (n2652gat), .I (I2354));
INVX1 gate1068(.O (n2500gat), .I (n2502gat));
INVX1 gate1069(.O (n2620gat), .I (n2622gat));
INVX1 gate1070(.O (n2612gat), .I (n2620gat));
INVX1 gate1071(.O (I2372), .I (n2612gat));
INVX1 gate1072(.O (n2606gat), .I (I2372));
INVX1 gate1073(.O (n2532gat), .I (n2625gat));
INVX1 gate1074(.O (I2376), .I (n2532gat));
INVX1 gate1075(.O (n2607gat), .I (I2376));
INVX1 gate1076(.O (n2540gat), .I (n2488gat));
INVX1 gate1077(.O (I2380), .I (n2540gat));
INVX1 gate1078(.O (n2608gat), .I (I2380));
INVX1 gate1079(.O (n2536gat), .I (n2624gat));
INVX1 gate1080(.O (I2385), .I (n2536gat));
INVX1 gate1081(.O (n2609gat), .I (I2385));
INVX1 gate1082(.O (n2487gat), .I (n2489gat));
INVX1 gate1083(.O (I2389), .I (n2487gat));
INVX1 gate1084(.O (n2610gat), .I (I2389));
INVX1 gate1085(.O (n2557gat), .I (n2621gat));
INVX1 gate1086(.O (I2394), .I (n2557gat));
INVX1 gate1087(.O (n2611gat), .I (I2394));
INVX1 gate1088(.O (I2400), .I (n2601gat));
INVX1 gate1089(.O (n2616gat), .I (I2400));
INVX1 gate1090(.O (I2403), .I (n2629gat));
INVX1 gate1091(.O (n2550gat), .I (I2403));
INVX1 gate1092(.O (I2414), .I (n2634gat));
INVX1 gate1093(.O (n2633gat), .I (I2414));
INVX1 gate1094(.O (I2417), .I (n2633gat));
INVX1 gate1095(.O (n2551gat), .I (I2417));
INVX1 gate1096(.O (I2420), .I (n2542gat));
INVX1 gate1097(.O (n2552gat), .I (I2420));
INVX1 gate1098(.O (n2632gat), .I (n2634gat));
INVX1 gate1099(.O (I2425), .I (n2632gat));
INVX1 gate1100(.O (n2553gat), .I (I2425));
INVX1 gate1101(.O (I2428), .I (n2541gat));
INVX1 gate1102(.O (n2554gat), .I (I2428));
INVX1 gate1103(.O (n2628gat), .I (n2630gat));
INVX1 gate1104(.O (I2433), .I (n2628gat));
INVX1 gate1105(.O (n2555gat), .I (I2433));
INVX1 gate1106(.O (I2439), .I (n2545gat));
INVX1 gate1107(.O (n2619gat), .I (I2439));
INVX1 gate1108(.O (n2504gat), .I (n2506gat));
INVX1 gate1109(.O (n2660gat), .I (n2655gat));
INVX1 gate1110(.O (n1528gat), .I (n2293gat));
INVX1 gate1111(.O (n1523gat), .I (n2219gat));
INVX1 gate1112(.O (n1592gat), .I (n1529gat));
INVX1 gate1113(.O (n2666gat), .I (n1704gat));
INVX1 gate1114(.O (n2422gat), .I (n3013gat));
INVX1 gate1115(.O (n2290gat), .I (n2202gat));
INVX1 gate1116(.O (n2081gat), .I (n2218gat));
INVX1 gate1117(.O (n2285gat), .I (n2397gat));
INVX1 gate1118(.O (n2359gat), .I (n2358gat));
INVX1 gate1119(.O (n1414gat), .I (n1415gat));
INVX1 gate1120(.O (n566gat), .I (n364gat));
INVX1 gate1121(.O (n1480gat), .I (n2292gat));
INVX1 gate1122(.O (n1301gat), .I (n1416gat));
INVX1 gate1123(.O (n1150gat), .I (n312gat));
INVX1 gate1124(.O (n873gat), .I (n316gat));
INVX1 gate1125(.O (n2011gat), .I (n2306gat));
INVX1 gate1126(.O (n1478gat), .I (n1481gat));
INVX1 gate1127(.O (n875gat), .I (n559gat));
INVX1 gate1128(.O (n1410gat), .I (n2357gat));
INVX1 gate1129(.O (n876gat), .I (n1347gat));
INVX1 gate1130(.O (n1160gat), .I (n1484gat));
INVX1 gate1131(.O (n1084gat), .I (n657gat));
INVX1 gate1132(.O (n983gat), .I (n320gat));
INVX1 gate1133(.O (n1482gat), .I (n2363gat));
INVX1 gate1134(.O (n1157gat), .I (n1483gat));
INVX1 gate1135(.O (n985gat), .I (n775gat));
INVX1 gate1136(.O (n1530gat), .I (n2364gat));
INVX1 gate1137(.O (n1307gat), .I (n1308gat));
INVX1 gate1138(.O (n1085gat), .I (n551gat));
INVX1 gate1139(.O (n1479gat), .I (n2291gat));
INVX1 gate1140(.O (n1348gat), .I (n1349gat));
INVX1 gate1141(.O (n2217gat), .I (n2206gat));
INVX1 gate1142(.O (n1591gat), .I (n2223gat));
INVX1 gate1143(.O (n1437gat), .I (n1438gat));
INVX1 gate1144(.O (n1832gat), .I (n1834gat));
INVX1 gate1145(.O (n1765gat), .I (n1767gat));
INVX1 gate1146(.O (n1878gat), .I (n1880gat));
INVX1 gate1147(.O (n1442gat), .I (n1831gat));
INVX1 gate1148(.O (n1444gat), .I (n1442gat));
INVX1 gate1149(.O (n1378gat), .I (n2975gat));
INVX1 gate1150(.O (n1322gat), .I (n2974gat));
INVX1 gate1151(.O (n1439gat), .I (n1486gat));
INVX1 gate1152(.O (n1370gat), .I (n1426gat));
INVX1 gate1153(.O (n1369gat), .I (n2966gat));
INVX1 gate1154(.O (n1366gat), .I (n1365gat));
INVX1 gate1155(.O (n1374gat), .I (n2979gat));
INVX1 gate1156(.O (n2162gat), .I (n2220gat));
INVX1 gate1157(.O (n1450gat), .I (n1423gat));
INVX1 gate1158(.O (n1427gat), .I (n1608gat));
INVX1 gate1159(.O (n1603gat), .I (n1831gat));
INVX1 gate1160(.O (n2082gat), .I (n2084gat));
INVX1 gate1161(.O (n1449gat), .I (n1494gat));
INVX1 gate1162(.O (n1590gat), .I (n1603gat));
INVX1 gate1163(.O (n1248gat), .I (n2954gat));
INVX1 gate1164(.O (n1418gat), .I (n1417gat));
INVX1 gate1165(.O (n1306gat), .I (n2964gat));
INVX1 gate1166(.O (n1353gat), .I (n1419gat));
INVX1 gate1167(.O (n1247gat), .I (n2958gat));
INVX1 gate1168(.O (n1355gat), .I (n1422gat));
INVX1 gate1169(.O (n1300gat), .I (n2963gat));
INVX1 gate1170(.O (n1487gat), .I (n1485gat));
INVX1 gate1171(.O (n1164gat), .I (n2953gat));
INVX1 gate1172(.O (n1356gat), .I (n1354gat));
INVX1 gate1173(.O (n1436gat), .I (n1435gat));
INVX1 gate1174(.O (n1106gat), .I (n2949gat));
INVX1 gate1175(.O (n1425gat), .I (n1421gat));
INVX1 gate1176(.O (n1105gat), .I (n2934gat));
INVX1 gate1177(.O (n1424gat), .I (n1420gat));
INVX1 gate1178(.O (n1309gat), .I (n2959gat));
INVX1 gate1179(.O (I2672), .I (n2143gat));
INVX1 gate1180(.O (n2142gat), .I (I2672));
INVX1 gate1181(.O (n1788gat), .I (n2142gat));
INVX1 gate1182(.O (I2684), .I (n2061gat));
INVX1 gate1183(.O (n2060gat), .I (I2684));
INVX1 gate1184(.O (n1786gat), .I (n2060gat));
INVX1 gate1185(.O (I2696), .I (n2139gat));
INVX1 gate1186(.O (n2138gat), .I (I2696));
INVX1 gate1187(.O (n1839gat), .I (n2138gat));
INVX1 gate1188(.O (n1897gat), .I (n1899gat));
INVX1 gate1189(.O (n1884gat), .I (n1897gat));
INVX1 gate1190(.O (n1848gat), .I (n1850gat));
INVX1 gate1191(.O (n1783gat), .I (n1848gat));
INVX1 gate1192(.O (n1548gat), .I (I2721));
INVX1 gate1193(.O (n1719gat), .I (n1548gat));
INVX1 gate1194(.O (n2137gat), .I (n2139gat));
INVX1 gate1195(.O (n1633gat), .I (n2137gat));
INVX1 gate1196(.O (n2059gat), .I (n2061gat));
INVX1 gate1197(.O (n1785gat), .I (n2059gat));
INVX1 gate1198(.O (I2731), .I (n1850gat));
INVX1 gate1199(.O (n1849gat), .I (I2731));
INVX1 gate1200(.O (n1784gat), .I (n1849gat));
INVX1 gate1201(.O (n1716gat), .I (I2736));
INVX1 gate1202(.O (n1635gat), .I (n1716gat));
INVX1 gate1203(.O (n2401gat), .I (n2403gat));
INVX1 gate1204(.O (n1989gat), .I (n2401gat));
INVX1 gate1205(.O (n2392gat), .I (n2394gat));
INVX1 gate1206(.O (n1918gat), .I (n2392gat));
INVX1 gate1207(.O (I2771), .I (n2440gat));
INVX1 gate1208(.O (n2439gat), .I (I2771));
INVX1 gate1209(.O (n1986gat), .I (n2439gat));
INVX1 gate1210(.O (n1866gat), .I (n1865gat));
INVX1 gate1211(.O (I2785), .I (n2407gat));
INVX1 gate1212(.O (n2406gat), .I (I2785));
INVX1 gate1213(.O (n2216gat), .I (n2406gat));
INVX1 gate1214(.O (n2345gat), .I (n2347gat));
INVX1 gate1215(.O (n1988gat), .I (n2345gat));
INVX1 gate1216(.O (n1735gat), .I (n1861gat));
INVX1 gate1217(.O (n1387gat), .I (n1389gat));
INVX1 gate1218(.O (n1694gat), .I (I2813));
INVX1 gate1219(.O (n1777gat), .I (n1694gat));
INVX1 gate1220(.O (n1781gat), .I (n1780gat));
INVX1 gate1221(.O (n2019gat), .I (n2021gat));
INVX1 gate1222(.O (n1549gat), .I (I2832));
INVX1 gate1223(.O (n1551gat), .I (n1549gat));
INVX1 gate1224(.O (I2837), .I (n2347gat));
INVX1 gate1225(.O (n2346gat), .I (I2837));
INVX1 gate1226(.O (n2152gat), .I (n2346gat));
INVX1 gate1227(.O (n2405gat), .I (n2407gat));
INVX1 gate1228(.O (n2351gat), .I (n2405gat));
INVX1 gate1229(.O (I2843), .I (n2403gat));
INVX1 gate1230(.O (n2402gat), .I (I2843));
INVX1 gate1231(.O (n2212gat), .I (n2402gat));
INVX1 gate1232(.O (I2847), .I (n2394gat));
INVX1 gate1233(.O (n2393gat), .I (I2847));
INVX1 gate1234(.O (n1991gat), .I (n2393gat));
INVX1 gate1235(.O (n1665gat), .I (n1666gat));
INVX1 gate1236(.O (n1517gat), .I (n1578gat));
INVX1 gate1237(.O (n1392gat), .I (n1394gat));
INVX1 gate1238(.O (I2873), .I (n1496gat));
INVX1 gate1239(.O (n1495gat), .I (I2873));
INVX1 gate1240(.O (n1685gat), .I (n1604gat));
INVX1 gate1241(.O (I2885), .I (n2091gat));
INVX1 gate1242(.O (n2090gat), .I (I2885));
INVX1 gate1243(.O (n1550gat), .I (I2890));
INVX1 gate1244(.O (n1552gat), .I (n1550gat));
INVX1 gate1245(.O (n1330gat), .I (n1332gat));
INVX1 gate1246(.O (n1738gat), .I (n1740gat));
INVX1 gate1247(.O (I2915), .I (n1740gat));
INVX1 gate1248(.O (n1739gat), .I (I2915));
INVX1 gate1249(.O (n1925gat), .I (n1920gat));
INVX1 gate1250(.O (n1917gat), .I (n1921gat));
INVX1 gate1251(.O (n2141gat), .I (n2143gat));
INVX1 gate1252(.O (n1787gat), .I (n2141gat));
INVX1 gate1253(.O (n1717gat), .I (I2926));
INVX1 gate1254(.O (n1859gat), .I (n1717gat));
INVX1 gate1255(.O (n1922gat), .I (n1798gat));
INVX1 gate1256(.O (n1713gat), .I (I2935));
INVX1 gate1257(.O (n1743gat), .I (n1713gat));
INVX1 gate1258(.O (n1923gat), .I (n1864gat));
INVX1 gate1259(.O (n1945gat), .I (n1690gat));
INVX1 gate1260(.O (I2953), .I (n2179gat));
INVX1 gate1261(.O (n2178gat), .I (I2953));
INVX1 gate1262(.O (n1661gat), .I (n1660gat));
INVX1 gate1263(.O (n1572gat), .I (n1576gat));
INVX1 gate1264(.O (n2438gat), .I (n2440gat));
INVX1 gate1265(.O (n2283gat), .I (n2438gat));
INVX1 gate1266(.O (n1520gat), .I (n1582gat));
INVX1 gate1267(.O (n1580gat), .I (n1577gat));
INVX1 gate1268(.O (n1990gat), .I (n2988gat));
INVX1 gate1269(.O (I2978), .I (n2190gat));
INVX1 gate1270(.O (n2189gat), .I (I2978));
INVX1 gate1271(.O (I2989), .I (n2135gat));
INVX1 gate1272(.O (n2134gat), .I (I2989));
INVX1 gate1273(.O (I3000), .I (n2262gat));
INVX1 gate1274(.O (n2261gat), .I (I3000));
INVX1 gate1275(.O (n2128gat), .I (n2129gat));
INVX1 gate1276(.O (n1836gat), .I (n1695gat));
INVX1 gate1277(.O (I3016), .I (n2182gat));
INVX1 gate1278(.O (n2181gat), .I (I3016));
INVX1 gate1279(.O (n1431gat), .I (n1433gat));
INVX1 gate1280(.O (n1314gat), .I (n1316gat));
INVX1 gate1281(.O (n1361gat), .I (n1363gat));
INVX1 gate1282(.O (I3056), .I (n1312gat));
INVX1 gate1283(.O (n1311gat), .I (I3056));
INVX1 gate1284(.O (n1707gat), .I (n1626gat));
INVX1 gate1285(.O (n1773gat), .I (n1775gat));
INVX1 gate1286(.O (n1659gat), .I (n2987gat));
INVX1 gate1287(.O (n1515gat), .I (n1521gat));
INVX1 gate1288(.O (n1736gat), .I (n1737gat));
INVX1 gate1289(.O (n1658gat), .I (n2216gat));
INVX1 gate1290(.O (n1724gat), .I (n1732gat));
INVX1 gate1291(.O (n1662gat), .I (n1663gat));
INVX1 gate1292(.O (n1656gat), .I (n1655gat));
INVX1 gate1293(.O (n1670gat), .I (n1667gat));
INVX1 gate1294(.O (n1569gat), .I (n1570gat));
INVX1 gate1295(.O (n1568gat), .I (n1575gat));
INVX1 gate1296(.O (n1727gat), .I (n1728gat));
INVX1 gate1297(.O (n1797gat), .I (n1801gat));
INVX1 gate1298(.O (n1730gat), .I (n1731gat));
INVX1 gate1299(.O (n1561gat), .I (n1571gat));
INVX1 gate1300(.O (n1668gat), .I (n1734gat));
INVX1 gate1301(.O (n1742gat), .I (n2216gat));
INVX1 gate1302(.O (n1671gat), .I (n1669gat));
INVX1 gate1303(.O (n1652gat), .I (n1657gat));
INVX1 gate1304(.O (n1648gat), .I (n1729gat));
INVX1 gate1305(.O (n1790gat), .I (n1726gat));
INVX1 gate1306(.O (n2004gat), .I (n1929gat));
INVX1 gate1307(.O (n1869gat), .I (n1871gat));
INVX1 gate1308(.O (I3143), .I (n2592gat));
INVX1 gate1309(.O (n2591gat), .I (I3143));
INVX1 gate1310(.O (n1584gat), .I (n2989gat));
INVX1 gate1311(.O (n1714gat), .I (I3149));
INVX1 gate1312(.O (n1718gat), .I (n1714gat));
INVX1 gate1313(.O (I3163), .I (n1508gat));
INVX1 gate1314(.O (n1507gat), .I (I3163));
INVX1 gate1315(.O (n1396gat), .I (n1401gat));
INVX1 gate1316(.O (I3168), .I (n1394gat));
INVX1 gate1317(.O (n1393gat), .I (I3168));
INVX1 gate1318(.O (n1409gat), .I (n1476gat));
INVX1 gate1319(.O (I3174), .I (n1899gat));
INVX1 gate1320(.O (n1898gat), .I (I3174));
INVX1 gate1321(.O (n1838gat), .I (n1898gat));
INVX1 gate1322(.O (n1712gat), .I (I3179));
INVX1 gate1323(.O (I3191), .I (n1678gat));
INVX1 gate1324(.O (n1677gat), .I (I3191));
INVX1 gate1325(.O (n2000gat), .I (n1412gat));
INVX1 gate1326(.O (n2001gat), .I (n1412gat));
INVX1 gate1327(.O (n1999gat), .I (n2001gat));
INVX1 gate1328(.O (n2307gat), .I (n2309gat));
INVX1 gate1329(.O (I3211), .I (n2663gat));
INVX1 gate1330(.O (n3018gat), .I (I3211));
INVX1 gate1331(.O (n2448gat), .I (n2450gat));
INVX1 gate1332(.O (n2661gat), .I (n2662gat));
INVX1 gate1333(.O (n2444gat), .I (n2446gat));
INVX1 gate1334(.O (I3235), .I (n2238gat));
INVX1 gate1335(.O (n3019gat), .I (I3235));
INVX1 gate1336(.O (n1310gat), .I (n1312gat));
INVX1 gate1337(.O (n199gat), .I (n87gat));
INVX1 gate1338(.O (n195gat), .I (n184gat));
INVX1 gate1339(.O (n827gat), .I (n204gat));
INVX1 gate1340(.O (n2093gat), .I (n2095gat));
INVX1 gate1341(.O (n2174gat), .I (n2176gat));
INVX1 gate1342(.O (I3273), .I (n2169gat));
INVX1 gate1343(.O (n2168gat), .I (I3273));
INVX1 gate1344(.O (n2452gat), .I (n2454gat));
INVX1 gate1345(.O (n1691gat), .I (n2452gat));
INVX1 gate1346(.O (I3287), .I (n1691gat));
INVX1 gate1347(.O (n3020gat), .I (I3287));
INVX1 gate1348(.O (I3290), .I (n1691gat));
INVX1 gate1349(.O (n3021gat), .I (I3290));
INVX1 gate1350(.O (I3293), .I (n1691gat));
INVX1 gate1351(.O (n3022gat), .I (I3293));
INVX1 gate1352(.O (n1699gat), .I (n2452gat));
INVX1 gate1353(.O (I3297), .I (n1699gat));
INVX1 gate1354(.O (n3023gat), .I (I3297));
INVX1 gate1355(.O (I3300), .I (n1699gat));
INVX1 gate1356(.O (n3024gat), .I (I3300));
INVX1 gate1357(.O (I3303), .I (n1691gat));
INVX1 gate1358(.O (n3025gat), .I (I3303));
INVX1 gate1359(.O (I3306), .I (n1699gat));
INVX1 gate1360(.O (n3026gat), .I (I3306));
INVX1 gate1361(.O (I3309), .I (n1699gat));
INVX1 gate1362(.O (n3027gat), .I (I3309));
INVX1 gate1363(.O (I3312), .I (n1699gat));
INVX1 gate1364(.O (n3028gat), .I (I3312));
INVX1 gate1365(.O (I3315), .I (n1869gat));
INVX1 gate1366(.O (n3029gat), .I (I3315));
INVX1 gate1367(.O (I3318), .I (n1869gat));
INVX1 gate1368(.O (n3030gat), .I (I3318));
INVX1 gate1369(.O (n2260gat), .I (n2262gat));
INVX1 gate1370(.O (n2257gat), .I (n2189gat));
INVX1 gate1371(.O (n2188gat), .I (n2190gat));
INVX1 gate1372(.O (n2187gat), .I (n3004gat));
INVX1 gate1373(.O (I3336), .I (n2040gat));
INVX1 gate1374(.O (n2039gat), .I (I3336));
INVX1 gate1375(.O (I3339), .I (n1775gat));
INVX1 gate1376(.O (n1774gat), .I (I3339));
INVX1 gate1377(.O (I3342), .I (n1316gat));
INVX1 gate1378(.O (n1315gat), .I (I3342));
INVX1 gate1379(.O (n2042gat), .I (n2044gat));
INVX1 gate1380(.O (n2035gat), .I (n2037gat));
INVX1 gate1381(.O (n2023gat), .I (n2025gat));
INVX1 gate1382(.O (n2097gat), .I (n2099gat));
INVX1 gate1383(.O (n1855gat), .I (n2014gat));
INVX1 gate1384(.O (I3387), .I (n2194gat));
INVX1 gate1385(.O (n3031gat), .I (I3387));
INVX1 gate1386(.O (I3390), .I (n2261gat));
INVX1 gate1387(.O (n3032gat), .I (I3390));
INVX1 gate1388(.O (n2256gat), .I (n3032gat));
INVX1 gate1389(.O (I3394), .I (n2260gat));
INVX1 gate1390(.O (n3033gat), .I (I3394));
INVX1 gate1391(.O (n2251gat), .I (n3033gat));
INVX1 gate1392(.O (n2184gat), .I (n3003gat));
INVX1 gate1393(.O (I3401), .I (n2192gat));
INVX1 gate1394(.O (n3034gat), .I (I3401));
INVX1 gate1395(.O (n2133gat), .I (n2135gat));
INVX1 gate1396(.O (n2131gat), .I (n2185gat));
INVX1 gate1397(.O (n2049gat), .I (n3001gat));
INVX1 gate1398(.O (I3412), .I (n2057gat));
INVX1 gate1399(.O (n3035gat), .I (I3412));
INVX1 gate1400(.O (n2253gat), .I (n2189gat));
INVX1 gate1401(.O (n2252gat), .I (n2260gat));
INVX1 gate1402(.O (n2248gat), .I (n3006gat));
INVX1 gate1403(.O (n2264gat), .I (n2266gat));
INVX1 gate1404(.O (I3429), .I (n2266gat));
INVX1 gate1405(.O (n2265gat), .I (I3429));
INVX1 gate1406(.O (n2492gat), .I (n2329gat));
INVX1 gate1407(.O (I3436), .I (n2492gat));
INVX1 gate1408(.O (n3036gat), .I (I3436));
INVX1 gate1409(.O (n1709gat), .I (n1849gat));
INVX1 gate1410(.O (n1845gat), .I (n2141gat));
INVX1 gate1411(.O (n1891gat), .I (n2059gat));
INVX1 gate1412(.O (n1963gat), .I (n2137gat));
INVX1 gate1413(.O (n1886gat), .I (n1897gat));
INVX1 gate1414(.O (n1968gat), .I (n1958gat));
INVX1 gate1415(.O (n1629gat), .I (n1895gat));
INVX1 gate1416(.O (n1631gat), .I (n1848gat));
INVX1 gate1417(.O (n1711gat), .I (n2990gat));
INVX1 gate1418(.O (n2200gat), .I (n2078gat));
INVX1 gate1419(.O (n2437gat), .I (n2195gat));
INVX1 gate1420(.O (I3457), .I (n2556gat));
INVX1 gate1421(.O (n3037gat), .I (I3457));
INVX1 gate1422(.O (n1956gat), .I (n1898gat));
INVX1 gate1423(.O (I3461), .I (n1956gat));
INVX1 gate1424(.O (n3038gat), .I (I3461));
INVX1 gate1425(.O (n1954gat), .I (n3038gat));
INVX1 gate1426(.O (I3465), .I (n1886gat));
INVX1 gate1427(.O (n3039gat), .I (I3465));
INVX1 gate1428(.O (n1888gat), .I (n3039gat));
INVX1 gate1429(.O (n2048gat), .I (n2994gat));
INVX1 gate1430(.O (I3472), .I (n2539gat));
INVX1 gate1431(.O (n3040gat), .I (I3472));
INVX1 gate1432(.O (n1969gat), .I (n2142gat));
INVX1 gate1433(.O (n1893gat), .I (n2060gat));
INVX1 gate1434(.O (n1892gat), .I (n2993gat));
INVX1 gate1435(.O (I3483), .I (n2436gat));
INVX1 gate1436(.O (n3041gat), .I (I3483));
INVX1 gate1437(.O (n2056gat), .I (n2998gat));
INVX1 gate1438(.O (I3491), .I (n2387gat));
INVX1 gate1439(.O (n3042gat), .I (I3491));
INVX1 gate1440(.O (I3494), .I (n1963gat));
INVX1 gate1441(.O (n3043gat), .I (I3494));
INVX1 gate1442(.O (n1960gat), .I (n3043gat));
INVX1 gate1443(.O (n1887gat), .I (n2138gat));
INVX1 gate1444(.O (n1961gat), .I (n2996gat));
INVX1 gate1445(.O (I3504), .I (n2330gat));
INVX1 gate1446(.O (n3044gat), .I (I3504));
INVX1 gate1447(.O (n2199gat), .I (n2147gat));
INVX1 gate1448(.O (I3509), .I (n2438gat));
INVX1 gate1449(.O (n3045gat), .I (I3509));
INVX1 gate1450(.O (n2332gat), .I (n3045gat));
INVX1 gate1451(.O (I3513), .I (n2439gat));
INVX1 gate1452(.O (n3046gat), .I (I3513));
INVX1 gate1453(.O (n2259gat), .I (n3046gat));
INVX1 gate1454(.O (n2328gat), .I (n3008gat));
INVX1 gate1455(.O (I3520), .I (n2498gat));
INVX1 gate1456(.O (n3047gat), .I (I3520));
INVX1 gate1457(.O (n2151gat), .I (n2193gat));
INVX1 gate1458(.O (n2209gat), .I (n3005gat));
INVX1 gate1459(.O (I3530), .I (n2396gat));
INVX1 gate1460(.O (n3048gat), .I (I3530));
INVX1 gate1461(.O (n2052gat), .I (n2393gat));
INVX1 gate1462(.O (n2058gat), .I (n2997gat));
INVX1 gate1463(.O (I3539), .I (n2198gat));
INVX1 gate1464(.O (n3049gat), .I (I3539));
INVX1 gate1465(.O (n2349gat), .I (n2215gat));
INVX1 gate1466(.O (n2281gat), .I (n3009gat));
INVX1 gate1467(.O (I3549), .I (n2197gat));
INVX1 gate1468(.O (n3050gat), .I (I3549));
INVX1 gate1469(.O (n2146gat), .I (n3002gat));
INVX1 gate1470(.O (I3558), .I (n2196gat));
INVX1 gate1471(.O (n3051gat), .I (I3558));
INVX1 gate1472(.O (n2031gat), .I (n2033gat));
INVX1 gate1473(.O (n2108gat), .I (n2110gat));
INVX1 gate1474(.O (I3587), .I (n2125gat));
INVX1 gate1475(.O (n2124gat), .I (I3587));
INVX1 gate1476(.O (n2123gat), .I (n2125gat));
INVX1 gate1477(.O (n2119gat), .I (n2121gat));
INVX1 gate1478(.O (n2115gat), .I (n2117gat));
INVX1 gate1479(.O (I3610), .I (n1882gat));
INVX1 gate1480(.O (n3052gat), .I (I3610));
INVX1 gate1481(.O (I3621), .I (n1975gat));
INVX1 gate1482(.O (n1974gat), .I (I3621));
INVX1 gate1483(.O (n1955gat), .I (n1956gat));
INVX1 gate1484(.O (n1970gat), .I (n1896gat));
INVX1 gate1485(.O (n1973gat), .I (n1975gat));
INVX1 gate1486(.O (n2558gat), .I (n2559gat));
INVX1 gate1487(.O (I3635), .I (n2558gat));
INVX1 gate1488(.O (n3053gat), .I (I3635));
INVX1 gate1489(.O (I3646), .I (n2644gat));
INVX1 gate1490(.O (n2643gat), .I (I3646));
INVX1 gate1491(.O (n2333gat), .I (n2438gat));
INVX1 gate1492(.O (n2564gat), .I (n2352gat));
INVX1 gate1493(.O (n2642gat), .I (n2644gat));
INVX1 gate1494(.O (n2636gat), .I (n2637gat));
INVX1 gate1495(.O (I3660), .I (n2636gat));
INVX1 gate1496(.O (n3054gat), .I (I3660));
INVX1 gate1497(.O (n88gat), .I (n84gat));
INVX1 gate1498(.O (n375gat), .I (n110gat));
INVX1 gate1499(.O (I3677), .I (n156gat));
INVX1 gate1500(.O (n155gat), .I (I3677));
INVX1 gate1501(.O (n253gat), .I (n1702gat));
INVX1 gate1502(.O (n150gat), .I (n152gat));
INVX1 gate1503(.O (I3691), .I (n152gat));
INVX1 gate1504(.O (n151gat), .I (I3691));
INVX1 gate1505(.O (n243gat), .I (n1702gat));
INVX1 gate1506(.O (n233gat), .I (n243gat));
INVX1 gate1507(.O (n154gat), .I (n156gat));
INVX1 gate1508(.O (n800gat), .I (n2874gat));
INVX1 gate1509(.O (I3703), .I (n2917gat));
INVX1 gate1510(.O (n3055gat), .I (I3703));
INVX1 gate1511(.O (n235gat), .I (n2878gat));
INVX1 gate1512(.O (I3713), .I (n2892gat));
INVX1 gate1513(.O (n3056gat), .I (I3713));
INVX1 gate1514(.O (n372gat), .I (n212gat));
INVX1 gate1515(.O (n329gat), .I (n331gat));
INVX1 gate1516(.O (I3736), .I (n388gat));
INVX1 gate1517(.O (n387gat), .I (I3736));
INVX1 gate1518(.O (n334gat), .I (n1700gat));
INVX1 gate1519(.O (n386gat), .I (n388gat));
INVX1 gate1520(.O (I3742), .I (n331gat));
INVX1 gate1521(.O (n330gat), .I (I3742));
INVX1 gate1522(.O (n1430gat), .I (n1700gat));
INVX1 gate1523(.O (n1490gat), .I (n1430gat));
INVX1 gate1524(.O (n452gat), .I (n2885gat));
INVX1 gate1525(.O (I3754), .I (n2900gat));
INVX1 gate1526(.O (n3057gat), .I (I3754));
INVX1 gate1527(.O (n333gat), .I (n2883gat));
INVX1 gate1528(.O (I3765), .I (n2929gat));
INVX1 gate1529(.O (n3058gat), .I (I3765));
INVX1 gate1530(.O (I3777), .I (n463gat));
INVX1 gate1531(.O (n462gat), .I (I3777));
INVX1 gate1532(.O (n325gat), .I (n327gat));
INVX1 gate1533(.O (n457gat), .I (n2884gat));
INVX1 gate1534(.O (n461gat), .I (n463gat));
INVX1 gate1535(.O (n458gat), .I (n2902gat));
INVX1 gate1536(.O (I3801), .I (n2925gat));
INVX1 gate1537(.O (n3059gat), .I (I3801));
INVX1 gate1538(.O (n144gat), .I (n247gat));
INVX1 gate1539(.O (I3808), .I (n327gat));
INVX1 gate1540(.O (n326gat), .I (I3808));
INVX1 gate1541(.O (n878gat), .I (n2879gat));
INVX1 gate1542(.O (I3817), .I (n2916gat));
INVX1 gate1543(.O (n3060gat), .I (I3817));
INVX1 gate1544(.O (n382gat), .I (n384gat));
INVX1 gate1545(.O (I3831), .I (n384gat));
INVX1 gate1546(.O (n383gat), .I (I3831));
INVX1 gate1547(.O (n134gat), .I (n2875gat));
INVX1 gate1548(.O (I3841), .I (n2899gat));
INVX1 gate1549(.O (n3061gat), .I (I3841));
INVX1 gate1550(.O (n254gat), .I (n256gat));
INVX1 gate1551(.O (n252gat), .I (n2877gat));
INVX1 gate1552(.O (n468gat), .I (n470gat));
INVX1 gate1553(.O (I3867), .I (n470gat));
INVX1 gate1554(.O (n469gat), .I (I3867));
INVX1 gate1555(.O (n381gat), .I (n2893gat));
INVX1 gate1556(.O (I3876), .I (n2926gat));
INVX1 gate1557(.O (n3062gat), .I (I3876));
INVX1 gate1558(.O (n241gat), .I (n140gat));
INVX1 gate1559(.O (I3882), .I (n256gat));
INVX1 gate1560(.O (n255gat), .I (I3882));
INVX1 gate1561(.O (n802gat), .I (n2882gat));
INVX1 gate1562(.O (I3891), .I (n2924gat));
INVX1 gate1563(.O (n3063gat), .I (I3891));
INVX1 gate1564(.O (n146gat), .I (n148gat));
INVX1 gate1565(.O (I3904), .I (n148gat));
INVX1 gate1566(.O (n147gat), .I (I3904));
INVX1 gate1567(.O (n380gat), .I (n2881gat));
INVX1 gate1568(.O (I3914), .I (n2923gat));
INVX1 gate1569(.O (n3064gat), .I (I3914));
INVX1 gate1570(.O (n69gat), .I (n68gat));
INVX1 gate1571(.O (n1885gat), .I (n2048gat));
INVX1 gate1572(.O (I3923), .I (n2710gat));
INVX1 gate1573(.O (n2707gat), .I (I3923));
INVX1 gate1574(.O (n16gat), .I (n564gat));
INVX1 gate1575(.O (n295gat), .I (n357gat));
INVX1 gate1576(.O (n11gat), .I (n12gat));
INVX1 gate1577(.O (n1889gat), .I (n1961gat));
INVX1 gate1578(.O (I3935), .I (n2704gat));
INVX1 gate1579(.O (n2700gat), .I (I3935));
INVX1 gate1580(.O (n2051gat), .I (n2056gat));
INVX1 gate1581(.O (I3941), .I (n2684gat));
INVX1 gate1582(.O (n2680gat), .I (I3941));
INVX1 gate1583(.O (n1350gat), .I (n1831gat));
INVX1 gate1584(.O (I3945), .I (n1350gat));
INVX1 gate1585(.O (n2696gat), .I (I3945));
INVX1 gate1586(.O (I3948), .I (n2696gat));
INVX1 gate1587(.O (n2692gat), .I (I3948));
INVX1 gate1588(.O (I3951), .I (n2448gat));
INVX1 gate1589(.O (n2683gat), .I (I3951));
INVX1 gate1590(.O (I3954), .I (n2683gat));
INVX1 gate1591(.O (n2679gat), .I (I3954));
INVX1 gate1592(.O (I3957), .I (n2450gat));
INVX1 gate1593(.O (n2449gat), .I (I3957));
INVX1 gate1594(.O (n1754gat), .I (n2449gat));
INVX1 gate1595(.O (I3962), .I (n2830gat));
INVX1 gate1596(.O (n2827gat), .I (I3962));
INVX1 gate1597(.O (n2590gat), .I (n2592gat));
INVX1 gate1598(.O (n2456gat), .I (n2458gat));
INVX1 gate1599(.O (n2512gat), .I (n2514gat));
INVX1 gate1600(.O (n1544gat), .I (n1625gat));
INVX1 gate1601(.O (n1769gat), .I (n1771gat));
INVX1 gate1602(.O (n1683gat), .I (n1756gat));
INVX1 gate1603(.O (n2167gat), .I (n2169gat));
INVX1 gate1604(.O (n2013gat), .I (I4000));
INVX1 gate1605(.O (n1791gat), .I (n2013gat));
INVX1 gate1606(.O (n2691gat), .I (n2695gat));
INVX1 gate1607(.O (n1518gat), .I (n1694gat));
INVX1 gate1608(.O (n2699gat), .I (n2703gat));
INVX1 gate1609(.O (n2159gat), .I (n1412gat));
INVX1 gate1610(.O (n2478gat), .I (n2579gat));
INVX1 gate1611(.O (I4014), .I (n2744gat));
INVX1 gate1612(.O (n2740gat), .I (I4014));
INVX1 gate1613(.O (n2158gat), .I (n1412gat));
INVX1 gate1614(.O (n2186gat), .I (n2613gat));
INVX1 gate1615(.O (I4020), .I (n2800gat));
INVX1 gate1616(.O (n2797gat), .I (I4020));
INVX1 gate1617(.O (n2288gat), .I (I4024));
INVX1 gate1618(.O (n1513gat), .I (n2288gat));
INVX1 gate1619(.O (n2537gat), .I (n2538gat));
INVX1 gate1620(.O (n2442gat), .I (n2483gat));
INVX1 gate1621(.O (n1334gat), .I (n1336gat));
INVX1 gate1622(.O (I4055), .I (n1748gat));
INVX1 gate1623(.O (n1747gat), .I (I4055));
INVX1 gate1624(.O (I4067), .I (n1675gat));
INVX1 gate1625(.O (n1674gat), .I (I4067));
INVX1 gate1626(.O (n1403gat), .I (n1402gat));
INVX1 gate1627(.O (I4081), .I (n1807gat));
INVX1 gate1628(.O (n1806gat), .I (I4081));
INVX1 gate1629(.O (n1634gat), .I (n1712gat));
INVX1 gate1630(.O (n1338gat), .I (n1340gat));
INVX1 gate1631(.O (I4105), .I (n1456gat));
INVX1 gate1632(.O (n1455gat), .I (I4105));
INVX1 gate1633(.O (I4108), .I (n1340gat));
INVX1 gate1634(.O (n1339gat), .I (I4108));
INVX1 gate1635(.O (n1505gat), .I (n2980gat));
INVX1 gate1636(.O (I4117), .I (n1505gat));
INVX1 gate1637(.O (n2758gat), .I (I4117));
INVX1 gate1638(.O (n2755gat), .I (n2758gat));
INVX1 gate1639(.O (n1546gat), .I (n2980gat));
INVX1 gate1640(.O (I4122), .I (n1546gat));
INVX1 gate1641(.O (n2752gat), .I (I4122));
INVX1 gate1642(.O (n2748gat), .I (n2752gat));
INVX1 gate1643(.O (n2012gat), .I (n2016gat));
INVX1 gate1644(.O (n2002gat), .I (n2008gat));
INVX1 gate1645(.O (I4129), .I (n3097gat));
INVX1 gate1646(.O (n2858gat), .I (I4129));
INVX1 gate1647(.O (n2857gat), .I (n2858gat));
INVX1 gate1648(.O (I4135), .I (n3098gat));
INVX1 gate1649(.O (n2766gat), .I (I4135));
INVX1 gate1650(.O (I4138), .I (n2766gat));
INVX1 gate1651(.O (n2765gat), .I (I4138));
INVX1 gate1652(.O (n1684gat), .I (n1759gat));
INVX1 gate1653(.O (n1632gat), .I (I4145));
INVX1 gate1654(.O (I4157), .I (n1525gat));
INVX1 gate1655(.O (n1524gat), .I (I4157));
INVX1 gate1656(.O (n1862gat), .I (n1863gat));
INVX1 gate1657(.O (n1919gat), .I (n1860gat));
INVX1 gate1658(.O (n1460gat), .I (n1462gat));
INVX1 gate1659(.O (I4185), .I (n1596gat));
INVX1 gate1660(.O (n1595gat), .I (I4185));
INVX1 gate1661(.O (n1454gat), .I (n1469gat));
INVX1 gate1662(.O (n1468gat), .I (n1519gat));
INVX1 gate1663(.O (I4194), .I (n1462gat));
INVX1 gate1664(.O (n1461gat), .I (I4194));
INVX1 gate1665(.O (n1477gat), .I (n2984gat));
INVX1 gate1666(.O (n1594gat), .I (n1596gat));
INVX1 gate1667(.O (I4212), .I (n1588gat));
INVX1 gate1668(.O (n1587gat), .I (I4212));
INVX1 gate1669(.O (n1681gat), .I (I4217));
INVX1 gate1670(.O (I4222), .I (n1761gat));
INVX1 gate1671(.O (n2751gat), .I (I4222));
INVX1 gate1672(.O (n2747gat), .I (n2751gat));
INVX1 gate1673(.O (I4227), .I (n1760gat));
INVX1 gate1674(.O (n2743gat), .I (I4227));
INVX1 gate1675(.O (n2739gat), .I (n2743gat));
INVX1 gate1676(.O (n1978gat), .I (n2286gat));
INVX1 gate1677(.O (I4233), .I (n1721gat));
INVX1 gate1678(.O (n2808gat), .I (I4233));
INVX1 gate1679(.O (I4236), .I (n2808gat));
INVX1 gate1680(.O (n2804gat), .I (I4236));
INVX1 gate1681(.O (n517gat), .I (n518gat));
INVX1 gate1682(.O (n417gat), .I (n418gat));
INVX1 gate1683(.O (n413gat), .I (n411gat));
INVX1 gate1684(.O (n412gat), .I (n522gat));
INVX1 gate1685(.O (n406gat), .I (n516gat));
INVX1 gate1686(.O (n407gat), .I (n355gat));
INVX1 gate1687(.O (n290gat), .I (n525gat));
INVX1 gate1688(.O (n527gat), .I (n356gat));
INVX1 gate1689(.O (n416gat), .I (n415gat));
INVX1 gate1690(.O (n528gat), .I (n521gat));
INVX1 gate1691(.O (n358gat), .I (n532gat));
INVX1 gate1692(.O (n639gat), .I (n523gat));
INVX1 gate1693(.O (n1111gat), .I (n635gat));
INVX1 gate1694(.O (n524gat), .I (n414gat));
INVX1 gate1695(.O (n1112gat), .I (n630gat));
INVX1 gate1696(.O (n741gat), .I (n629gat));
INVX1 gate1697(.O (n633gat), .I (n634gat));
INVX1 gate1698(.O (n926gat), .I (n632gat));
INVX1 gate1699(.O (n670gat), .I (n636gat));
INVX1 gate1700(.O (n1123gat), .I (n632gat));
INVX1 gate1701(.O (n1007gat), .I (n635gat));
INVX1 gate1702(.O (n1006gat), .I (n630gat));
INVX1 gate1703(.O (I4309), .I (n2941gat));
INVX1 gate1704(.O (n2814gat), .I (I4309));
INVX1 gate1705(.O (I4312), .I (n2814gat));
INVX1 gate1706(.O (n2811gat), .I (I4312));
INVX1 gate1707(.O (n1002gat), .I (n2946gat));
INVX1 gate1708(.O (I4329), .I (n2950gat));
INVX1 gate1709(.O (n2813gat), .I (I4329));
INVX1 gate1710(.O (I4332), .I (n2813gat));
INVX1 gate1711(.O (n2810gat), .I (I4332));
INVX1 gate1712(.O (n888gat), .I (n2933gat));
INVX1 gate1713(.O (I4349), .I (n2935gat));
INVX1 gate1714(.O (n2818gat), .I (I4349));
INVX1 gate1715(.O (I4352), .I (n2818gat));
INVX1 gate1716(.O (n2816gat), .I (I4352));
INVX1 gate1717(.O (n898gat), .I (n2940gat));
INVX1 gate1718(.O (I4369), .I (n2937gat));
INVX1 gate1719(.O (n2817gat), .I (I4369));
INVX1 gate1720(.O (I4372), .I (n2817gat));
INVX1 gate1721(.O (n2815gat), .I (I4372));
INVX1 gate1722(.O (n1179gat), .I (n2947gat));
INVX1 gate1723(.O (I4389), .I (n2956gat));
INVX1 gate1724(.O (n2824gat), .I (I4389));
INVX1 gate1725(.O (I4392), .I (n2824gat));
INVX1 gate1726(.O (n2821gat), .I (I4392));
INVX1 gate1727(.O (n897gat), .I (n2939gat));
INVX1 gate1728(.O (I4409), .I (n2938gat));
INVX1 gate1729(.O (n2823gat), .I (I4409));
INVX1 gate1730(.O (I4412), .I (n2823gat));
INVX1 gate1731(.O (n2820gat), .I (I4412));
INVX1 gate1732(.O (n894gat), .I (n2932gat));
INVX1 gate1733(.O (I4429), .I (n2936gat));
INVX1 gate1734(.O (n2829gat), .I (I4429));
INVX1 gate1735(.O (I4432), .I (n2829gat));
INVX1 gate1736(.O (n2826gat), .I (I4432));
INVX1 gate1737(.O (n1180gat), .I (n2948gat));
INVX1 gate1738(.O (I4449), .I (n2955gat));
INVX1 gate1739(.O (n2828gat), .I (I4449));
INVX1 gate1740(.O (I4452), .I (n2828gat));
INVX1 gate1741(.O (n2825gat), .I (I4452));
INVX1 gate1742(.O (n671gat), .I (n673gat));
INVX1 gate1743(.O (n628gat), .I (n631gat));
INVX1 gate1744(.O (n976gat), .I (n628gat));
INVX1 gate1745(.O (I4475), .I (n2951gat));
INVX1 gate1746(.O (n2807gat), .I (I4475));
INVX1 gate1747(.O (I4478), .I (n2807gat));
INVX1 gate1748(.O (n2803gat), .I (I4478));
INVX1 gate1749(.O (n2127gat), .I (n2389gat));
INVX1 gate1750(.O (I4482), .I (n2127gat));
INVX1 gate1751(.O (n2682gat), .I (I4482));
INVX1 gate1752(.O (I4485), .I (n2682gat));
INVX1 gate1753(.O (n2678gat), .I (I4485));
INVX1 gate1754(.O (n2046gat), .I (n2269gat));
INVX1 gate1755(.O (I4489), .I (n2046gat));
INVX1 gate1756(.O (n2681gat), .I (I4489));
INVX1 gate1757(.O (I4492), .I (n2681gat));
INVX1 gate1758(.O (n2677gat), .I (I4492));
INVX1 gate1759(.O (n1708gat), .I (n2338gat));
INVX1 gate1760(.O (I4496), .I (n1708gat));
INVX1 gate1761(.O (n2688gat), .I (I4496));
INVX1 gate1762(.O (I4499), .I (n2688gat));
INVX1 gate1763(.O (n2686gat), .I (I4499));
INVX1 gate1764(.O (n455gat), .I (n291gat));
INVX1 gate1765(.O (n2237gat), .I (n2646gat));
INVX1 gate1766(.O (I4506), .I (n2764gat));
INVX1 gate1767(.O (n2763gat), .I (I4506));
INVX1 gate1768(.O (n1782gat), .I (n2971gat));
INVX1 gate1769(.O (I4512), .I (n2762gat));
INVX1 gate1770(.O (n2760gat), .I (I4512));
INVX1 gate1771(.O (n2325gat), .I (n3010gat));
INVX1 gate1772(.O (I4518), .I (n2761gat));
INVX1 gate1773(.O (n2759gat), .I (I4518));
INVX1 gate1774(.O (n2245gat), .I (n504gat));
INVX1 gate1775(.O (I4524), .I (n2757gat));
INVX1 gate1776(.O (n2754gat), .I (I4524));
INVX1 gate1777(.O (n2244gat), .I (n567gat));
INVX1 gate1778(.O (I4530), .I (n2756gat));
INVX1 gate1779(.O (n2753gat), .I (I4530));
INVX1 gate1780(.O (n2243gat), .I (n55gat));
INVX1 gate1781(.O (I4536), .I (n2750gat));
INVX1 gate1782(.O (n2746gat), .I (I4536));
INVX1 gate1783(.O (n2246gat), .I (n933gat));
INVX1 gate1784(.O (I4542), .I (n2749gat));
INVX1 gate1785(.O (n2745gat), .I (I4542));
INVX1 gate1786(.O (n2384gat), .I (n43gat));
INVX1 gate1787(.O (I4548), .I (n2742gat));
INVX1 gate1788(.O (n2738gat), .I (I4548));
INVX1 gate1789(.O (n2385gat), .I (n748gat));
INVX1 gate1790(.O (I4554), .I (n2741gat));
INVX1 gate1791(.O (n2737gat), .I (I4554));
INVX1 gate1792(.O (n1286gat), .I (n1269gat));
INVX1 gate1793(.O (I4558), .I (n1286gat));
INVX1 gate1794(.O (n2687gat), .I (I4558));
INVX1 gate1795(.O (n2685gat), .I (n2687gat));
INVX1 gate1796(.O (n1328gat), .I (n1224gat));
INVX1 gate1797(.O (n1381gat), .I (n1328gat));
INVX1 gate1798(.O (n1384gat), .I (n2184gat));
INVX1 gate1799(.O (I4566), .I (n2694gat));
INVX1 gate1800(.O (n2690gat), .I (I4566));
INVX1 gate1801(.O (n1382gat), .I (n1280gat));
INVX1 gate1802(.O (n1451gat), .I (n1382gat));
INVX1 gate1803(.O (n1453gat), .I (n2187gat));
INVX1 gate1804(.O (I4573), .I (n2693gat));
INVX1 gate1805(.O (n2689gat), .I (I4573));
INVX1 gate1806(.O (n927gat), .I (n1133gat));
INVX1 gate1807(.O (n925gat), .I (n927gat));
INVX1 gate1808(.O (n1452gat), .I (n2049gat));
INVX1 gate1809(.O (I4580), .I (n2702gat));
INVX1 gate1810(.O (n2698gat), .I (I4580));
INVX1 gate1811(.O (n923gat), .I (n1043gat));
INVX1 gate1812(.O (n921gat), .I (n923gat));
INVX1 gate1813(.O (n1890gat), .I (n2328gat));
INVX1 gate1814(.O (I4587), .I (n2701gat));
INVX1 gate1815(.O (n2697gat), .I (I4587));
INVX1 gate1816(.O (n850gat), .I (n929gat));
INVX1 gate1817(.O (n739gat), .I (n850gat));
INVX1 gate1818(.O (n1841gat), .I (n2058gat));
INVX1 gate1819(.O (I4594), .I (n2709gat));
INVX1 gate1820(.O (n2706gat), .I (I4594));
INVX1 gate1821(.O (n922gat), .I (n1119gat));
INVX1 gate1822(.O (n848gat), .I (n922gat));
INVX1 gate1823(.O (n2047gat), .I (n2209gat));
INVX1 gate1824(.O (I4601), .I (n2708gat));
INVX1 gate1825(.O (n2705gat), .I (I4601));
INVX1 gate1826(.O (n924gat), .I (n1070gat));
INVX1 gate1827(.O (n849gat), .I (n924gat));
INVX1 gate1828(.O (n2050gat), .I (n2146gat));
INVX1 gate1829(.O (I4608), .I (n2799gat));
INVX1 gate1830(.O (n2796gat), .I (I4608));
INVX1 gate1831(.O (n1118gat), .I (n1033gat));
INVX1 gate1832(.O (n1032gat), .I (n1118gat));
INVX1 gate1833(.O (n2054gat), .I (n2281gat));
INVX1 gate1834(.O (I4615), .I (n2798gat));
INVX1 gate1835(.O (n2795gat), .I (I4615));
INVX1 gate1836(.O (I4620), .I (n1745gat));
INVX1 gate1837(.O (n2806gat), .I (I4620));
INVX1 gate1838(.O (I4623), .I (n2806gat));
INVX1 gate1839(.O (n2802gat), .I (I4623));
INVX1 gate1840(.O (I4626), .I (n1871gat));
INVX1 gate1841(.O (n1870gat), .I (I4626));
INVX1 gate1842(.O (n1086gat), .I (n1870gat));
INVX1 gate1843(.O (I4630), .I (n1086gat));
INVX1 gate1844(.O (n2805gat), .I (I4630));
INVX1 gate1845(.O (I4633), .I (n2805gat));
INVX1 gate1846(.O (n2801gat), .I (I4633));
INVX1 gate1847(.O (n67gat), .I (n85gat));
INVX1 gate1848(.O (n71gat), .I (n180gat));
INVX1 gate1849(.O (n1840gat), .I (n1892gat));
INVX1 gate1850(.O (I4642), .I (n2812gat));
INVX1 gate1851(.O (n2809gat), .I (I4642));
INVX1 gate1852(.O (n76gat), .I (n82gat));
INVX1 gate1853(.O (n14gat), .I (n186gat));
INVX1 gate1854(.O (n1842gat), .I (n1711gat));
INVX1 gate1855(.O (I4651), .I (n2822gat));
INVX1 gate1856(.O (n2819gat), .I (I4651));
INVX1 gate1857(.O (I4654), .I (n2819gat));
INVX1 gate1858(.O (n3104gat), .I (I4654));
INVX1 gate1859(.O (I4657), .I (n2809gat));
INVX1 gate1860(.O (n3105gat), .I (I4657));
INVX1 gate1861(.O (I4660), .I (n2801gat));
INVX1 gate1862(.O (n3106gat), .I (I4660));
INVX1 gate1863(.O (I4663), .I (n2802gat));
INVX1 gate1864(.O (n3107gat), .I (I4663));
INVX1 gate1865(.O (I4666), .I (n2795gat));
INVX1 gate1866(.O (n3108gat), .I (I4666));
INVX1 gate1867(.O (I4669), .I (n2796gat));
INVX1 gate1868(.O (n3109gat), .I (I4669));
INVX1 gate1869(.O (I4672), .I (n2705gat));
INVX1 gate1870(.O (n3110gat), .I (I4672));
INVX1 gate1871(.O (I4675), .I (n2706gat));
INVX1 gate1872(.O (n3111gat), .I (I4675));
INVX1 gate1873(.O (I4678), .I (n2697gat));
INVX1 gate1874(.O (n3112gat), .I (I4678));
INVX1 gate1875(.O (I4681), .I (n2698gat));
INVX1 gate1876(.O (n3113gat), .I (I4681));
INVX1 gate1877(.O (I4684), .I (n2689gat));
INVX1 gate1878(.O (n3114gat), .I (I4684));
INVX1 gate1879(.O (I4687), .I (n2690gat));
INVX1 gate1880(.O (n3115gat), .I (I4687));
INVX1 gate1881(.O (I4690), .I (n2685gat));
INVX1 gate1882(.O (n3116gat), .I (I4690));
INVX1 gate1883(.O (I4693), .I (n2737gat));
INVX1 gate1884(.O (n3117gat), .I (I4693));
INVX1 gate1885(.O (I4696), .I (n2738gat));
INVX1 gate1886(.O (n3118gat), .I (I4696));
INVX1 gate1887(.O (I4699), .I (n2745gat));
INVX1 gate1888(.O (n3119gat), .I (I4699));
INVX1 gate1889(.O (I4702), .I (n2746gat));
INVX1 gate1890(.O (n3120gat), .I (I4702));
INVX1 gate1891(.O (I4705), .I (n2753gat));
INVX1 gate1892(.O (n3121gat), .I (I4705));
INVX1 gate1893(.O (I4708), .I (n2754gat));
INVX1 gate1894(.O (n3122gat), .I (I4708));
INVX1 gate1895(.O (I4711), .I (n2759gat));
INVX1 gate1896(.O (n3123gat), .I (I4711));
INVX1 gate1897(.O (I4714), .I (n2760gat));
INVX1 gate1898(.O (n3124gat), .I (I4714));
INVX1 gate1899(.O (I4717), .I (n2763gat));
INVX1 gate1900(.O (n3125gat), .I (I4717));
INVX1 gate1901(.O (I4720), .I (n2686gat));
INVX1 gate1902(.O (n3126gat), .I (I4720));
INVX1 gate1903(.O (I4723), .I (n2677gat));
INVX1 gate1904(.O (n3127gat), .I (I4723));
INVX1 gate1905(.O (I4726), .I (n2678gat));
INVX1 gate1906(.O (n3128gat), .I (I4726));
INVX1 gate1907(.O (I4729), .I (n2803gat));
INVX1 gate1908(.O (n3129gat), .I (I4729));
INVX1 gate1909(.O (I4732), .I (n2825gat));
INVX1 gate1910(.O (n3130gat), .I (I4732));
INVX1 gate1911(.O (I4735), .I (n2826gat));
INVX1 gate1912(.O (n3131gat), .I (I4735));
INVX1 gate1913(.O (I4738), .I (n2820gat));
INVX1 gate1914(.O (n3132gat), .I (I4738));
INVX1 gate1915(.O (I4741), .I (n2821gat));
INVX1 gate1916(.O (n3133gat), .I (I4741));
INVX1 gate1917(.O (I4744), .I (n2815gat));
INVX1 gate1918(.O (n3134gat), .I (I4744));
INVX1 gate1919(.O (I4747), .I (n2816gat));
INVX1 gate1920(.O (n3135gat), .I (I4747));
INVX1 gate1921(.O (I4750), .I (n2810gat));
INVX1 gate1922(.O (n3136gat), .I (I4750));
INVX1 gate1923(.O (I4753), .I (n2811gat));
INVX1 gate1924(.O (n3137gat), .I (I4753));
INVX1 gate1925(.O (I4756), .I (n2804gat));
INVX1 gate1926(.O (n3138gat), .I (I4756));
INVX1 gate1927(.O (I4759), .I (n2739gat));
INVX1 gate1928(.O (n3139gat), .I (I4759));
INVX1 gate1929(.O (I4762), .I (n2747gat));
INVX1 gate1930(.O (n3140gat), .I (I4762));
INVX1 gate1931(.O (I4765), .I (n2748gat));
INVX1 gate1932(.O (n3141gat), .I (I4765));
INVX1 gate1933(.O (I4768), .I (n2755gat));
INVX1 gate1934(.O (n3142gat), .I (I4768));
INVX1 gate1935(.O (I4771), .I (n2797gat));
INVX1 gate1936(.O (n3143gat), .I (I4771));
INVX1 gate1937(.O (I4774), .I (n2740gat));
INVX1 gate1938(.O (n3144gat), .I (I4774));
INVX1 gate1939(.O (I4777), .I (n2699gat));
INVX1 gate1940(.O (n3145gat), .I (I4777));
INVX1 gate1941(.O (I4780), .I (n2691gat));
INVX1 gate1942(.O (n3146gat), .I (I4780));
INVX1 gate1943(.O (I4783), .I (n2827gat));
INVX1 gate1944(.O (n3147gat), .I (I4783));
INVX1 gate1945(.O (I4786), .I (n2679gat));
INVX1 gate1946(.O (n3148gat), .I (I4786));
INVX1 gate1947(.O (I4789), .I (n2692gat));
INVX1 gate1948(.O (n3149gat), .I (I4789));
INVX1 gate1949(.O (I4792), .I (n2680gat));
INVX1 gate1950(.O (n3150gat), .I (I4792));
INVX1 gate1951(.O (I4795), .I (n2700gat));
INVX1 gate1952(.O (n3151gat), .I (I4795));
INVX1 gate1953(.O (I4798), .I (n2707gat));
INVX1 gate1954(.O (n3152gat), .I (I4798));
OR2X1 gate1955(.O (n2897gat), .I1 (n648gat), .I2 (n442gat));
OR4X1 gate1956(.O (n1213gat), .I1 (n1214gat), .I2 (n1215gat), .I3 (n1216gat), .I4 (n1217gat));
OR2X1 gate1957(.O (n2906gat), .I1 (n745gat), .I2 (n638gat));
OR2X1 gate1958(.O (n2889gat), .I1 (n423gat), .I2 (n362gat));
OR4X1 gate1959(.O (n748gat), .I1 (n749gat), .I2 (n750gat), .I3 (n751gat), .I4 (n752gat));
OR4X1 gate1960(.O (n258gat), .I1 (n259gat), .I2 (n260gat), .I3 (n261gat), .I4 (n262gat));
OR4X1 gate1961(.O (n1013gat), .I1 (n1014gat), .I2 (n1015gat), .I3 (n1016gat), .I4 (n1017gat));
OR4X1 gate1962(.O (n475gat), .I1 (n476gat), .I2 (n477gat), .I3 (n478gat), .I4 (n479gat));
OR4X1 gate1963(.O (n43gat), .I1 (n44gat), .I2 (n45gat), .I3 (n46gat), .I4 (n47gat));
OR2X1 gate1964(.O (n2786gat), .I1 (n3091gat), .I2 (n3092gat));
OR4X1 gate1965(.O (n167gat), .I1 (n168gat), .I2 (n169gat), .I3 (n170gat), .I4 (n171gat));
OR4X1 gate1966(.O (n906gat), .I1 (n907gat), .I2 (n908gat), .I3 (n909gat), .I4 (n910gat));
OR4X1 gate1967(.O (n343gat), .I1 (n344gat), .I2 (n345gat), .I3 (n346gat), .I4 (n347gat));
OR4X1 gate1968(.O (n55gat), .I1 (n56gat), .I2 (n57gat), .I3 (n58gat), .I4 (n59gat));
OR2X1 gate1969(.O (n2914gat), .I1 (n768gat), .I2 (n655gat));
OR2X1 gate1970(.O (n2928gat), .I1 (n963gat), .I2 (n868gat));
OR2X1 gate1971(.O (n2927gat), .I1 (n962gat), .I2 (n959gat));
OR4X1 gate1972(.O (n944gat), .I1 (n945gat), .I2 (n946gat), .I3 (n947gat), .I4 (n948gat));
OR2X1 gate1973(.O (n2896gat), .I1 (n647gat), .I2 (n441gat));
OR2X1 gate1974(.O (n2922gat), .I1 (n967gat), .I2 (n792gat));
OR4X1 gate1975(.O (n1228gat), .I1 (n1229gat), .I2 (n1230gat), .I3 (n1231gat), .I4 (n1232gat));
OR2X1 gate1976(.O (n2894gat), .I1 (n443gat), .I2 (n439gat));
OR2X1 gate1977(.O (n2921gat), .I1 (n966gat), .I2 (n790gat));
OR2X1 gate1978(.O (n2895gat), .I1 (n444gat), .I2 (n440gat));
OR4X1 gate1979(.O (n1050gat), .I1 (n1051gat), .I2 (n1052gat), .I3 (n1053gat), .I4 (n1054gat));
OR4X1 gate1980(.O (n933gat), .I1 (n934gat), .I2 (n935gat), .I3 (n936gat), .I4 (n937gat));
OR4X1 gate1981(.O (n709gat), .I1 (n710gat), .I2 (n711gat), .I3 (n712gat), .I4 (n713gat));
OR4X1 gate1982(.O (n728gat), .I1 (n729gat), .I2 (n730gat), .I3 (n731gat), .I4 (n732gat));
OR4X1 gate1983(.O (n493gat), .I1 (n494gat), .I2 (n495gat), .I3 (n496gat), .I4 (n497gat));
OR4X1 gate1984(.O (n504gat), .I1 (n505gat), .I2 (n506gat), .I3 (n507gat), .I4 (n508gat));
OR3X1 gate1985(.O (I1277), .I1 (n2860gat), .I2 (n2855gat), .I3 (n2863gat));
OR3X1 gate1986(.O (I1278), .I1 (n740gat), .I2 (n3030gat), .I3 (I1277));
OR2X1 gate1987(.O (n2913gat), .I1 (n767gat), .I2 (n653gat));
OR2X1 gate1988(.O (n2920gat), .I1 (n867gat), .I2 (n771gat));
OR2X1 gate1989(.O (n2905gat), .I1 (n964gat), .I2 (n961gat));
OR4X1 gate1990(.O (n803gat), .I1 (n804gat), .I2 (n805gat), .I3 (n806gat), .I4 (n807gat));
OR4X1 gate1991(.O (n586gat), .I1 (n587gat), .I2 (n588gat), .I3 (n589gat), .I4 (n590gat));
OR2X1 gate1992(.O (n2898gat), .I1 (n447gat), .I2 (n445gat));
OR4X1 gate1993(.O (n686gat), .I1 (n687gat), .I2 (n688gat), .I3 (n689gat), .I4 (n690gat));
OR4X1 gate1994(.O (n567gat), .I1 (n568gat), .I2 (n569gat), .I3 (n570gat), .I4 (n571gat));
OR3X1 gate1995(.O (I1515), .I1 (n2474gat), .I2 (n2524gat), .I3 (n2831gat));
OR3X1 gate1996(.O (I1516), .I1 (n2466gat), .I2 (n2462gat), .I3 (I1515));
OR3X1 gate1997(.O (I1584), .I1 (n2353gat), .I2 (n2284gat), .I3 (n2354gat));
OR3X1 gate1998(.O (I1585), .I1 (n2356gat), .I2 (n2214gat), .I3 (I1584));
OR2X1 gate1999(.O (n2989gat), .I1 (n1693gat), .I2 (n1692gat));
OR3X1 gate2000(.O (I1723), .I1 (n2354gat), .I2 (n2353gat), .I3 (n2214gat));
OR3X1 gate2001(.O (I1724), .I1 (n2355gat), .I2 (n2443gat), .I3 (I1723));
OR3X1 gate2002(.O (I1733), .I1 (n2286gat), .I2 (n2428gat), .I3 (n2289gat));
OR3X1 gate2003(.O (I1734), .I1 (n1604gat), .I2 (n2214gat), .I3 (I1733));
OR2X1 gate2004(.O (n2918gat), .I1 (n769gat), .I2 (n759gat));
OR2X1 gate2005(.O (n2952gat), .I1 (n1076gat), .I2 (n1075gat));
OR2X1 gate2006(.O (n2919gat), .I1 (n766gat), .I2 (n760gat));
OR4X1 gate2007(.O (n1184gat), .I1 (n1185gat), .I2 (n1186gat), .I3 (n1187gat), .I4 (n1188gat));
OR2X1 gate2008(.O (n2910gat), .I1 (n645gat), .I2 (n644gat));
OR2X1 gate2009(.O (n2907gat), .I1 (n646gat), .I2 (n641gat));
OR2X1 gate2010(.O (n2970gat), .I1 (n1383gat), .I2 (n1327gat));
OR2X1 gate2011(.O (n2911gat), .I1 (n761gat), .I2 (n651gat));
OR2X1 gate2012(.O (n2912gat), .I1 (n762gat), .I2 (n652gat));
OR2X1 gate2013(.O (n2909gat), .I1 (n765gat), .I2 (n643gat));
OR4X1 gate2014(.O (n1201gat), .I1 (n1202gat), .I2 (n1203gat), .I3 (n1204gat), .I4 (n1205gat));
OR4X1 gate2015(.O (n1269gat), .I1 (n1270gat), .I2 (n1271gat), .I3 (n1272gat), .I4 (n1273gat));
OR2X1 gate2016(.O (n2908gat), .I1 (n763gat), .I2 (n642gat));
OR2X1 gate2017(.O (n2971gat), .I1 (n1287gat), .I2 (n1285gat));
OR3X1 gate2018(.O (n2904gat), .I1 (n793gat), .I2 (n664gat), .I3 (n556gat));
OR3X1 gate2019(.O (n2891gat), .I1 (n795gat), .I2 (n656gat), .I3 (n368gat));
OR3X1 gate2020(.O (n2903gat), .I1 (n794gat), .I2 (n773gat), .I3 (n662gat));
OR3X1 gate2021(.O (n2915gat), .I1 (n965gat), .I2 (n960gat), .I3 (n661gat));
OR4X1 gate2022(.O (n779gat), .I1 (n780gat), .I2 (n781gat), .I3 (n782gat), .I4 (n783gat));
OR3X1 gate2023(.O (n2901gat), .I1 (n558gat), .I2 (n555gat), .I3 (n450gat));
OR3X1 gate2024(.O (n2890gat), .I1 (n654gat), .I2 (n557gat), .I3 (n371gat));
OR2X1 gate2025(.O (n2876gat), .I1 (n874gat), .I2 (n132gat));
OR3X1 gate2026(.O (n2888gat), .I1 (n663gat), .I2 (n649gat), .I3 (n449gat));
OR3X1 gate2027(.O (n2887gat), .I1 (n791gat), .I2 (n650gat), .I3 (n370gat));
OR3X1 gate2028(.O (n2886gat), .I1 (n774gat), .I2 (n764gat), .I3 (n369gat));
OR4X1 gate2029(.O (n221gat), .I1 (n222gat), .I2 (n223gat), .I3 (n224gat), .I4 (n225gat));
OR4X1 gate2030(.O (n120gat), .I1 (n121gat), .I2 (n122gat), .I3 (n123gat), .I4 (n124gat));
OR2X1 gate2031(.O (n3010gat), .I1 (n2460gat), .I2 (n2423gat));
OR2X1 gate2032(.O (n3016gat), .I1 (n2596gat), .I2 (n2595gat));
OR4X1 gate2033(.O (n2568gat), .I1 (n2569gat), .I2 (n2570gat), .I3 (n2571gat), .I4 (n2572gat));
OR4X1 gate2034(.O (n2409gat), .I1 (n2410gat), .I2 (n2411gat), .I3 (n2412gat), .I4 (n2413gat));
OR2X1 gate2035(.O (n2579gat), .I1 (n2580gat), .I2 (n2581gat));
OR2X1 gate2036(.O (n3014gat), .I1 (n2567gat), .I2 (n2499gat));
OR2X1 gate2037(.O (n2880gat), .I1 (n299gat), .I2 (n207gat));
OR2X1 gate2038(.O (n2646gat), .I1 (n2647gat), .I2 (n2648gat));
OR4X1 gate2039(.O (n2601gat), .I1 (n2602gat), .I2 (n2603gat), .I3 (n2604gat), .I4 (n2605gat));
OR4X1 gate2040(.O (n2545gat), .I1 (n2546gat), .I2 (n2547gat), .I3 (n2548gat), .I4 (n2549gat));
OR2X1 gate2041(.O (n2613gat), .I1 (n2614gat), .I2 (n2615gat));
OR2X1 gate2042(.O (n3013gat), .I1 (n2461gat), .I2 (n2421gat));
OR4X1 gate2043(.O (n2930gat), .I1 (n1153gat), .I2 (n1151gat), .I3 (n982gat), .I4 (n877gat));
OR4X1 gate2044(.O (n2957gat), .I1 (n1159gat), .I2 (n1158gat), .I3 (n1156gat), .I4 (n1155gat));
OR2X1 gate2045(.O (n2975gat), .I1 (n1443gat), .I2 (n1325gat));
OR2X1 gate2046(.O (n2974gat), .I1 (n1321gat), .I2 (n1320gat));
OR2X1 gate2047(.O (n2966gat), .I1 (n1368gat), .I2 (n1258gat));
OR2X1 gate2048(.O (n2979gat), .I1 (n1373gat), .I2 (n1372gat));
OR4X1 gate2049(.O (n2978gat), .I1 (n1441gat), .I2 (n1440gat), .I3 (n1371gat), .I4 (n1367gat));
OR2X1 gate2050(.O (n2982gat), .I1 (n1504gat), .I2 (n1502gat));
OR2X1 gate2051(.O (n2954gat), .I1 (n1250gat), .I2 (n1103gat));
OR2X1 gate2052(.O (n2964gat), .I1 (n1304gat), .I2 (n1249gat));
OR2X1 gate2053(.O (n2958gat), .I1 (n1246gat), .I2 (n1161gat));
OR2X1 gate2054(.O (n2963gat), .I1 (n1291gat), .I2 (n1245gat));
OR4X1 gate2055(.O (n2973gat), .I1 (n1352gat), .I2 (n1351gat), .I3 (n1303gat), .I4 (n1302gat));
OR2X1 gate2056(.O (n2953gat), .I1 (n1163gat), .I2 (n1102gat));
OR2X1 gate2057(.O (n2949gat), .I1 (n1101gat), .I2 (n996gat));
OR2X1 gate2058(.O (n2934gat), .I1 (n1104gat), .I2 (n887gat));
OR2X1 gate2059(.O (n2959gat), .I1 (n1305gat), .I2 (n1162gat));
OR4X1 gate2060(.O (n2977gat), .I1 (n1360gat), .I2 (n1359gat), .I3 (n1358gat), .I4 (n1357gat));
OR3X1 gate2061(.O (I2720), .I1 (n1788gat), .I2 (n1786gat), .I3 (n1839gat));
OR3X1 gate2062(.O (I2721), .I1 (n1884gat), .I2 (n1783gat), .I3 (I2720));
OR3X1 gate2063(.O (I2735), .I1 (n1788gat), .I2 (n1884gat), .I3 (n1633gat));
OR3X1 gate2064(.O (I2736), .I1 (n1785gat), .I2 (n1784gat), .I3 (I2735));
OR3X1 gate2065(.O (I2812), .I1 (n1703gat), .I2 (n1704gat), .I3 (n1778gat));
OR4X1 gate2066(.O (I2813), .I1 (n1609gat), .I2 (n1702gat), .I3 (n1700gat), .I4 (I2812));
OR3X1 gate2067(.O (I2831), .I1 (n1839gat), .I2 (n1786gat), .I3 (n1788gat));
OR3X1 gate2068(.O (I2832), .I1 (n1884gat), .I2 (n1784gat), .I3 (I2831));
OR3X1 gate2069(.O (I2889), .I1 (n1784gat), .I2 (n1633gat), .I3 (n1884gat));
OR3X1 gate2070(.O (I2890), .I1 (n1788gat), .I2 (n1786gat), .I3 (I2889));
OR3X1 gate2071(.O (I2925), .I1 (n1784gat), .I2 (n1785gat), .I3 (n1633gat));
OR3X1 gate2072(.O (I2926), .I1 (n1884gat), .I2 (n1787gat), .I3 (I2925));
OR3X1 gate2073(.O (I2934), .I1 (n1784gat), .I2 (n1839gat), .I3 (n1788gat));
OR3X1 gate2074(.O (I2935), .I1 (n1785gat), .I2 (n1884gat), .I3 (I2934));
OR2X1 gate2075(.O (n2988gat), .I1 (n1733gat), .I2 (n1581gat));
OR2X1 gate2076(.O (n2983gat), .I1 (n2079gat), .I2 (n2073gat));
OR2X1 gate2077(.O (n2987gat), .I1 (n1574gat), .I2 (n1573gat));
OR3X1 gate2078(.O (n2992gat), .I1 (n1723gat), .I2 (n1647gat), .I3 (n1646gat));
OR3X1 gate2079(.O (n2986gat), .I1 (n1650gat), .I2 (n1649gat), .I3 (n1563gat));
OR3X1 gate2080(.O (n2991gat), .I1 (n1654gat), .I2 (n1653gat), .I3 (n1644gat));
OR3X1 gate2081(.O (I3148), .I1 (n1839gat), .I2 (n1884gat), .I3 (n1784gat));
OR3X1 gate2082(.O (I3149), .I1 (n1786gat), .I2 (n1787gat), .I3 (I3148));
OR3X1 gate2083(.O (I3178), .I1 (n1838gat), .I2 (n1785gat), .I3 (n1788gat));
OR3X1 gate2084(.O (I3179), .I1 (n1839gat), .I2 (n1784gat), .I3 (I3178));
OR3X1 gate2085(.O (n2981gat), .I1 (n1413gat), .I2 (n1408gat), .I3 (n1407gat));
OR2X1 gate2086(.O (n3000gat), .I1 (n2000gat), .I2 (n1999gat));
OR3X1 gate2087(.O (n3004gat), .I1 (n2258gat), .I2 (n2257gat), .I3 (n2255gat));
OR2X1 gate2088(.O (n3003gat), .I1 (n2256gat), .I2 (n2251gat));
OR2X1 gate2089(.O (n3001gat), .I1 (n2132gat), .I2 (n2130gat));
OR2X1 gate2090(.O (n3006gat), .I1 (n2253gat), .I2 (n2252gat));
OR2X1 gate2091(.O (n3007gat), .I1 (n2250gat), .I2 (n2249gat));
OR2X1 gate2092(.O (n2990gat), .I1 (n1710gat), .I2 (n1630gat));
OR2X1 gate2093(.O (n2994gat), .I1 (n1954gat), .I2 (n1888gat));
OR3X1 gate2094(.O (n2993gat), .I1 (n1894gat), .I2 (n1847gat), .I3 (n1846gat));
OR2X1 gate2095(.O (n2998gat), .I1 (n2055gat), .I2 (n1967gat));
OR3X1 gate2096(.O (n2996gat), .I1 (n1960gat), .I2 (n1959gat), .I3 (n1957gat));
OR2X1 gate2097(.O (n3008gat), .I1 (n2332gat), .I2 (n2259gat));
OR2X1 gate2098(.O (n3005gat), .I1 (n2211gat), .I2 (n2210gat));
OR3X1 gate2099(.O (n2997gat), .I1 (n2053gat), .I2 (n2052gat), .I3 (n1964gat));
OR2X1 gate2100(.O (n3009gat), .I1 (n2350gat), .I2 (n2282gat));
OR3X1 gate2101(.O (n3002gat), .I1 (n2213gat), .I2 (n2150gat), .I3 (n2149gat));
OR2X1 gate2102(.O (n2995gat), .I1 (n1962gat), .I2 (n1955gat));
OR2X1 gate2103(.O (n2999gat), .I1 (n1972gat), .I2 (n1971gat));
OR2X1 gate2104(.O (n3011gat), .I1 (n2333gat), .I2 (n2331gat));
OR2X1 gate2105(.O (n3015gat), .I1 (n2566gat), .I2 (n2565gat));
OR3X1 gate2106(.O (n2874gat), .I1 (n141gat), .I2 (n38gat), .I3 (n37gat));
OR2X1 gate2107(.O (n2917gat), .I1 (n1074gat), .I2 (n872gat));
OR2X1 gate2108(.O (n2878gat), .I1 (n234gat), .I2 (n137gat));
OR2X1 gate2109(.O (n2892gat), .I1 (n378gat), .I2 (n377gat));
OR3X1 gate2110(.O (n2885gat), .I1 (n250gat), .I2 (n249gat), .I3 (n248gat));
OR3X1 gate2111(.O (n2900gat), .I1 (n869gat), .I2 (n453gat), .I3 (n448gat));
OR2X1 gate2112(.O (n2883gat), .I1 (n251gat), .I2 (n244gat));
OR3X1 gate2113(.O (n2929gat), .I1 (n974gat), .I2 (n973gat), .I3 (n870gat));
OR2X1 gate2114(.O (n2884gat), .I1 (n246gat), .I2 (n245gat));
OR2X1 gate2115(.O (n2902gat), .I1 (n460gat), .I2 (n459gat));
OR3X1 gate2116(.O (n2925gat), .I1 (n975gat), .I2 (n972gat), .I3 (n969gat));
OR2X1 gate2117(.O (n2879gat), .I1 (n145gat), .I2 (n143gat));
OR3X1 gate2118(.O (n2916gat), .I1 (n971gat), .I2 (n970gat), .I3 (n968gat));
OR3X1 gate2119(.O (n2875gat), .I1 (n142gat), .I2 (n40gat), .I3 (n39gat));
OR3X1 gate2120(.O (n2899gat), .I1 (n772gat), .I2 (n451gat), .I3 (n446gat));
OR2X1 gate2121(.O (n2877gat), .I1 (n139gat), .I2 (n136gat));
OR2X1 gate2122(.O (n2893gat), .I1 (n391gat), .I2 (n390gat));
OR2X1 gate2123(.O (n2926gat), .I1 (n1083gat), .I2 (n1077gat));
OR2X1 gate2124(.O (n2882gat), .I1 (n242gat), .I2 (n240gat));
OR2X1 gate2125(.O (n2924gat), .I1 (n871gat), .I2 (n797gat));
OR3X1 gate2126(.O (n2881gat), .I1 (n324gat), .I2 (n238gat), .I3 (n237gat));
OR2X1 gate2127(.O (n2923gat), .I1 (n1082gat), .I2 (n796gat));
OR2X1 gate2128(.O (n2710gat), .I1 (n69gat), .I2 (n1885gat));
OR2X1 gate2129(.O (n2704gat), .I1 (n11gat), .I2 (n1889gat));
OR2X1 gate2130(.O (n2684gat), .I1 (n1599gat), .I2 (n2051gat));
OR2X1 gate2131(.O (n2830gat), .I1 (n2444gat), .I2 (n1754gat));
OR3X1 gate2132(.O (I3999), .I1 (n2167gat), .I2 (n2031gat), .I3 (n2174gat));
OR4X1 gate2133(.O (I4000), .I1 (n2108gat), .I2 (n2093gat), .I3 (n2035gat), .I4 (I3999));
OR2X1 gate2134(.O (n2695gat), .I1 (n1586gat), .I2 (n1791gat));
OR2X1 gate2135(.O (n2703gat), .I1 (n1755gat), .I2 (n1518gat));
OR2X1 gate2136(.O (n2744gat), .I1 (n2159gat), .I2 (n2478gat));
OR2X1 gate2137(.O (n2800gat), .I1 (n2158gat), .I2 (n2186gat));
OR3X1 gate2138(.O (I4023), .I1 (n2443gat), .I2 (n2290gat), .I3 (n2214gat));
OR3X1 gate2139(.O (I4024), .I1 (n2353gat), .I2 (n2284gat), .I3 (I4023));
OR4X1 gate2140(.O (n2980gat), .I1 (n1470gat), .I2 (n1400gat), .I3 (n1399gat), .I4 (n1398gat));
OR3X1 gate2141(.O (I4144), .I1 (n1633gat), .I2 (n1838gat), .I3 (n1786gat));
OR3X1 gate2142(.O (I4145), .I1 (n1788gat), .I2 (n1784gat), .I3 (I4144));
OR2X1 gate2143(.O (n2984gat), .I1 (n1467gat), .I2 (n1466gat));
OR4X1 gate2144(.O (n2985gat), .I1 (n1686gat), .I2 (n1533gat), .I3 (n1532gat), .I4 (n1531gat));
OR3X1 gate2145(.O (I4216), .I1 (n1427gat), .I2 (n1595gat), .I3 (n1677gat));
OR3X1 gate2146(.O (I4217), .I1 (n1392gat), .I2 (n2989gat), .I3 (I4216));
OR4X1 gate2147(.O (n2931gat), .I1 (n1100gat), .I2 (n994gat), .I3 (n989gat), .I4 (n880gat));
OR2X1 gate2148(.O (n2943gat), .I1 (n1012gat), .I2 (n905gat));
OR2X1 gate2149(.O (n2941gat), .I1 (n1003gat), .I2 (n902gat));
OR4X1 gate2150(.O (n2946gat), .I1 (n1099gat), .I2 (n998gat), .I3 (n995gat), .I4 (n980gat));
OR2X1 gate2151(.O (n2960gat), .I1 (n1175gat), .I2 (n1174gat));
OR2X1 gate2152(.O (n2950gat), .I1 (n1001gat), .I2 (n999gat));
OR2X1 gate2153(.O (n2969gat), .I1 (n1323gat), .I2 (n1264gat));
OR4X1 gate2154(.O (n2933gat), .I1 (n981gat), .I2 (n890gat), .I3 (n889gat), .I4 (n886gat));
OR2X1 gate2155(.O (n2935gat), .I1 (n892gat), .I2 (n891gat));
OR2X1 gate2156(.O (n2942gat), .I1 (n904gat), .I2 (n903gat));
OR4X1 gate2157(.O (n2940gat), .I1 (n1152gat), .I2 (n1092gat), .I3 (n997gat), .I4 (n993gat));
OR2X1 gate2158(.O (n2937gat), .I1 (n900gat), .I2 (n895gat));
OR4X1 gate2159(.O (n2947gat), .I1 (n1094gat), .I2 (n1093gat), .I3 (n988gat), .I4 (n984gat));
OR2X1 gate2160(.O (n2965gat), .I1 (n1267gat), .I2 (n1257gat));
OR2X1 gate2161(.O (n2956gat), .I1 (n1178gat), .I2 (n1116gat));
OR2X1 gate2162(.O (n2961gat), .I1 (n1375gat), .I2 (n1324gat));
OR4X1 gate2163(.O (n2939gat), .I1 (n1091gat), .I2 (n1088gat), .I3 (n992gat), .I4 (n987gat));
OR2X1 gate2164(.O (n2938gat), .I1 (n899gat), .I2 (n896gat));
OR2X1 gate2165(.O (n2967gat), .I1 (n1262gat), .I2 (n1260gat));
OR4X1 gate2166(.O (n2932gat), .I1 (n1098gat), .I2 (n1090gat), .I3 (n986gat), .I4 (n885gat));
OR2X1 gate2167(.O (n2936gat), .I1 (n901gat), .I2 (n893gat));
OR4X1 gate2168(.O (n2948gat), .I1 (n1097gat), .I2 (n1089gat), .I3 (n1087gat), .I4 (n991gat));
OR2X1 gate2169(.O (n2968gat), .I1 (n1326gat), .I2 (n1261gat));
OR2X1 gate2170(.O (n2955gat), .I1 (n1177gat), .I2 (n1115gat));
OR2X1 gate2171(.O (n2944gat), .I1 (n977gat), .I2 (n976gat));
OR4X1 gate2172(.O (n2945gat), .I1 (n1096gat), .I2 (n1095gat), .I3 (n990gat), .I4 (n979gat));
OR2X1 gate2173(.O (n2962gat), .I1 (n1176gat), .I2 (n1173gat));
OR2X1 gate2174(.O (n2951gat), .I1 (n1004gat), .I2 (n1000gat));
OR2X1 gate2175(.O (n2764gat), .I1 (n1029gat), .I2 (n2237gat));
OR2X1 gate2176(.O (n2762gat), .I1 (n1028gat), .I2 (n1782gat));
OR2X1 gate2177(.O (n2761gat), .I1 (n1031gat), .I2 (n2325gat));
OR2X1 gate2178(.O (n2757gat), .I1 (n1030gat), .I2 (n2245gat));
OR2X1 gate2179(.O (n2756gat), .I1 (n1011gat), .I2 (n2244gat));
OR2X1 gate2180(.O (n2750gat), .I1 (n1181gat), .I2 (n2243gat));
OR2X1 gate2181(.O (n2749gat), .I1 (n1010gat), .I2 (n2246gat));
OR2X1 gate2182(.O (n2742gat), .I1 (n1005gat), .I2 (n2384gat));
OR2X1 gate2183(.O (n2741gat), .I1 (n1182gat), .I2 (n2385gat));
OR2X1 gate2184(.O (n2694gat), .I1 (n1381gat), .I2 (n1384gat));
OR2X1 gate2185(.O (n2693gat), .I1 (n1451gat), .I2 (n1453gat));
OR2X1 gate2186(.O (n2702gat), .I1 (n925gat), .I2 (n1452gat));
OR2X1 gate2187(.O (n2701gat), .I1 (n921gat), .I2 (n1890gat));
OR2X1 gate2188(.O (n2709gat), .I1 (n739gat), .I2 (n1841gat));
OR2X1 gate2189(.O (n2708gat), .I1 (n848gat), .I2 (n2047gat));
OR2X1 gate2190(.O (n2799gat), .I1 (n849gat), .I2 (n2050gat));
OR2X1 gate2191(.O (n2798gat), .I1 (n1032gat), .I2 (n2054gat));
OR3X1 gate2192(.O (n2812gat), .I1 (n73gat), .I2 (n70gat), .I3 (n1840gat));
OR3X1 gate2193(.O (n2822gat), .I1 (n77gat), .I2 (n13gat), .I3 (n1842gat));
NR2X1 gate2194(.O (n421gat), .I1 (n2715gat), .I2 (n2723gat));
NR2X1 gate2195(.O (n648gat), .I1 (n373gat), .I2 (n2669gat));
NR2X1 gate2196(.O (n442gat), .I1 (n2844gat), .I2 (n856gat));
NR2X1 gate2197(.O (n1499gat), .I1 (n396gat), .I2 (n401gat));
NR2X1 gate2198(.O (n1616gat), .I1 (n918gat), .I2 (n396gat));
NR2X1 gate2199(.O (n1614gat), .I1 (n396gat), .I2 (n845gat));
NR3X1 gate2200(.O (n1641gat), .I1 (n1645gat), .I2 (n1553gat), .I3 (n1559gat));
NR3X1 gate2201(.O (n1642gat), .I1 (n1559gat), .I2 (n1616gat), .I3 (n1645gat));
NR3X1 gate2202(.O (n1556gat), .I1 (n1614gat), .I2 (n1645gat), .I3 (n1616gat));
NR3X1 gate2203(.O (n1557gat), .I1 (n1553gat), .I2 (n1645gat), .I3 (n1614gat));
NR3X1 gate2204(.O (n1639gat), .I1 (n1499gat), .I2 (n1559gat), .I3 (n1553gat));
NR4X1 gate2205(.O (n1605gat), .I1 (n1614gat), .I2 (n1616gat), .I3 (n1499gat), .I4 (n396gat));
NR3X1 gate2206(.O (n1555gat), .I1 (n1616gat), .I2 (n1559gat), .I3 (n1499gat));
NR3X1 gate2207(.O (n1558gat), .I1 (n1614gat), .I2 (n1553gat), .I3 (n1499gat));
NR2X1 gate2208(.O (n1256gat), .I1 (n392gat), .I2 (n702gat));
NR2X1 gate2209(.O (n1117gat), .I1 (n720gat), .I2 (n725gat));
NR2X1 gate2210(.O (n1618gat), .I1 (n1319gat), .I2 (n1447gat));
NR2X1 gate2211(.O (n1114gat), .I1 (n725gat), .I2 (n721gat));
NR2X1 gate2212(.O (n1621gat), .I1 (n1319gat), .I2 (n1380gat));
NR2X1 gate2213(.O (n1318gat), .I1 (n392gat), .I2 (n701gat));
NR2X1 gate2214(.O (n1619gat), .I1 (n1447gat), .I2 (n1446gat));
NR2X1 gate2215(.O (n1622gat), .I1 (n1380gat), .I2 (n1446gat));
NR3X1 gate2216(.O (n1214gat), .I1 (n1218gat), .I2 (n1219gat), .I3 (n1220gat));
NR3X1 gate2217(.O (n1215gat), .I1 (n1218gat), .I2 (n1221gat), .I3 (n1222gat));
NR3X1 gate2218(.O (n1216gat), .I1 (n1223gat), .I2 (n1219gat), .I3 (n1222gat));
NR3X1 gate2219(.O (n1217gat), .I1 (n1223gat), .I2 (n1221gat), .I3 (n1220gat));
NR2X1 gate2220(.O (n745gat), .I1 (n2716gat), .I2 (n2867gat));
NR2X1 gate2221(.O (n638gat), .I1 (n2715gat), .I2 (n2868gat));
NR2X1 gate2222(.O (n423gat), .I1 (n2724gat), .I2 (n2726gat));
NR2X1 gate2223(.O (n362gat), .I1 (n2723gat), .I2 (n2727gat));
NR3X1 gate2224(.O (n749gat), .I1 (n753gat), .I2 (n754gat), .I3 (n755gat));
NR3X1 gate2225(.O (n750gat), .I1 (n753gat), .I2 (n756gat), .I3 (n757gat));
NR3X1 gate2226(.O (n751gat), .I1 (n758gat), .I2 (n754gat), .I3 (n757gat));
NR3X1 gate2227(.O (n752gat), .I1 (n758gat), .I2 (n756gat), .I3 (n755gat));
NR3X1 gate2228(.O (n259gat), .I1 (n263gat), .I2 (n264gat), .I3 (n265gat));
NR3X1 gate2229(.O (n260gat), .I1 (n263gat), .I2 (n266gat), .I3 (n267gat));
NR3X1 gate2230(.O (n261gat), .I1 (n268gat), .I2 (n264gat), .I3 (n267gat));
NR3X1 gate2231(.O (n262gat), .I1 (n268gat), .I2 (n266gat), .I3 (n265gat));
NR3X1 gate2232(.O (n1014gat), .I1 (n1018gat), .I2 (n1019gat), .I3 (n1020gat));
NR3X1 gate2233(.O (n1015gat), .I1 (n1018gat), .I2 (n1021gat), .I3 (n1022gat));
NR3X1 gate2234(.O (n1016gat), .I1 (n1023gat), .I2 (n1019gat), .I3 (n1022gat));
NR3X1 gate2235(.O (n1017gat), .I1 (n1023gat), .I2 (n1021gat), .I3 (n1020gat));
NR3X1 gate2236(.O (n476gat), .I1 (n480gat), .I2 (n481gat), .I3 (n482gat));
NR3X1 gate2237(.O (n477gat), .I1 (n480gat), .I2 (n483gat), .I3 (n484gat));
NR3X1 gate2238(.O (n478gat), .I1 (n485gat), .I2 (n481gat), .I3 (n484gat));
NR3X1 gate2239(.O (n479gat), .I1 (n485gat), .I2 (n483gat), .I3 (n482gat));
NR3X1 gate2240(.O (n44gat), .I1 (n48gat), .I2 (n49gat), .I3 (n50gat));
NR3X1 gate2241(.O (n45gat), .I1 (n48gat), .I2 (n51gat), .I3 (n52gat));
NR3X1 gate2242(.O (n46gat), .I1 (n53gat), .I2 (n49gat), .I3 (n52gat));
NR3X1 gate2243(.O (n47gat), .I1 (n53gat), .I2 (n51gat), .I3 (n50gat));
NR2X1 gate2244(.O (n1376gat), .I1 (n724gat), .I2 (n720gat));
NR2X1 gate2245(.O (n1617gat), .I1 (n1319gat), .I2 (n1448gat));
NR2X1 gate2246(.O (n1377gat), .I1 (n724gat), .I2 (n721gat));
NR2X1 gate2247(.O (n1624gat), .I1 (n1319gat), .I2 (n1379gat));
NR2X1 gate2248(.O (n1113gat), .I1 (n393gat), .I2 (n701gat));
NR2X1 gate2249(.O (n1501gat), .I1 (n1448gat), .I2 (n1500gat));
NR2X1 gate2250(.O (n1623gat), .I1 (n1379gat), .I2 (n1446gat));
NR2X1 gate2251(.O (n1620gat), .I1 (n1448gat), .I2 (n1446gat));
NR2X1 gate2252(.O (n1827gat), .I1 (n2729gat), .I2 (n2317gat));
NR2X1 gate2253(.O (n1817gat), .I1 (n1819gat), .I2 (n1823gat));
NR2X1 gate2254(.O (n1935gat), .I1 (n1816gat), .I2 (n1828gat));
NR2X1 gate2255(.O (n529gat), .I1 (n2724gat), .I2 (n2715gat));
NR2X1 gate2256(.O (n361gat), .I1 (n2859gat), .I2 (n2726gat));
NR3X1 gate2257(.O (n168gat), .I1 (n172gat), .I2 (n173gat), .I3 (n174gat));
NR3X1 gate2258(.O (n169gat), .I1 (n172gat), .I2 (n175gat), .I3 (n176gat));
NR3X1 gate2259(.O (n170gat), .I1 (n177gat), .I2 (n173gat), .I3 (n176gat));
NR3X1 gate2260(.O (n171gat), .I1 (n177gat), .I2 (n175gat), .I3 (n174gat));
NR3X1 gate2261(.O (n907gat), .I1 (n911gat), .I2 (n912gat), .I3 (n913gat));
NR3X1 gate2262(.O (n908gat), .I1 (n911gat), .I2 (n914gat), .I3 (n915gat));
NR3X1 gate2263(.O (n909gat), .I1 (n916gat), .I2 (n912gat), .I3 (n915gat));
NR3X1 gate2264(.O (n910gat), .I1 (n916gat), .I2 (n914gat), .I3 (n913gat));
NR3X1 gate2265(.O (n344gat), .I1 (n348gat), .I2 (n349gat), .I3 (n350gat));
NR3X1 gate2266(.O (n345gat), .I1 (n348gat), .I2 (n351gat), .I3 (n352gat));
NR3X1 gate2267(.O (n346gat), .I1 (n353gat), .I2 (n349gat), .I3 (n352gat));
NR3X1 gate2268(.O (n347gat), .I1 (n353gat), .I2 (n351gat), .I3 (n350gat));
NR3X1 gate2269(.O (n56gat), .I1 (n60gat), .I2 (n61gat), .I3 (n62gat));
NR3X1 gate2270(.O (n57gat), .I1 (n60gat), .I2 (n63gat), .I3 (n64gat));
NR3X1 gate2271(.O (n58gat), .I1 (n65gat), .I2 (n61gat), .I3 (n64gat));
NR3X1 gate2272(.O (n59gat), .I1 (n65gat), .I2 (n63gat), .I3 (n62gat));
NR2X1 gate2273(.O (n768gat), .I1 (n373gat), .I2 (n2731gat));
NR2X1 gate2274(.O (n655gat), .I1 (n856gat), .I2 (n2718gat));
NR2X1 gate2275(.O (n963gat), .I1 (n856gat), .I2 (n2838gat));
NR2X1 gate2276(.O (n868gat), .I1 (n2775gat), .I2 (n373gat));
NR2X1 gate2277(.O (n962gat), .I1 (n856gat), .I2 (n2711gat));
NR2X1 gate2278(.O (n959gat), .I1 (n373gat), .I2 (n2734gat));
NR3X1 gate2279(.O (n945gat), .I1 (n949gat), .I2 (n950gat), .I3 (n951gat));
NR3X1 gate2280(.O (n946gat), .I1 (n949gat), .I2 (n952gat), .I3 (n953gat));
NR3X1 gate2281(.O (n947gat), .I1 (n954gat), .I2 (n950gat), .I3 (n953gat));
NR3X1 gate2282(.O (n948gat), .I1 (n954gat), .I2 (n952gat), .I3 (n951gat));
NR2X1 gate2283(.O (n647gat), .I1 (n2792gat), .I2 (n373gat));
NR2X1 gate2284(.O (n441gat), .I1 (n856gat), .I2 (n2846gat));
NR2X1 gate2285(.O (n967gat), .I1 (n373gat), .I2 (n2672gat));
NR2X1 gate2286(.O (n792gat), .I1 (n2852gat), .I2 (n856gat));
NR3X1 gate2287(.O (n1229gat), .I1 (n1233gat), .I2 (n1234gat), .I3 (n1235gat));
NR3X1 gate2288(.O (n1230gat), .I1 (n1233gat), .I2 (n1236gat), .I3 (n1237gat));
NR3X1 gate2289(.O (n1231gat), .I1 (n1238gat), .I2 (n1234gat), .I3 (n1237gat));
NR3X1 gate2290(.O (n1232gat), .I1 (n1238gat), .I2 (n1236gat), .I3 (n1235gat));
NR2X1 gate2291(.O (n443gat), .I1 (n2778gat), .I2 (n373gat));
NR2X1 gate2292(.O (n439gat), .I1 (n856gat), .I2 (n2836gat));
NR2X1 gate2293(.O (n966gat), .I1 (n2789gat), .I2 (n373gat));
NR2X1 gate2294(.O (n790gat), .I1 (n856gat), .I2 (n2840gat));
NR2X1 gate2295(.O (n444gat), .I1 (n373gat), .I2 (n2781gat));
NR2X1 gate2296(.O (n440gat), .I1 (n856gat), .I2 (n2842gat));
NR3X1 gate2297(.O (n1051gat), .I1 (n1055gat), .I2 (n1056gat), .I3 (n1057gat));
NR3X1 gate2298(.O (n1052gat), .I1 (n1055gat), .I2 (n1058gat), .I3 (n1059gat));
NR3X1 gate2299(.O (n1053gat), .I1 (n1060gat), .I2 (n1056gat), .I3 (n1059gat));
NR3X1 gate2300(.O (n1054gat), .I1 (n1060gat), .I2 (n1058gat), .I3 (n1057gat));
NR3X1 gate2301(.O (n934gat), .I1 (n938gat), .I2 (n939gat), .I3 (n940gat));
NR3X1 gate2302(.O (n935gat), .I1 (n938gat), .I2 (n941gat), .I3 (n942gat));
NR3X1 gate2303(.O (n936gat), .I1 (n943gat), .I2 (n939gat), .I3 (n942gat));
NR3X1 gate2304(.O (n937gat), .I1 (n943gat), .I2 (n941gat), .I3 (n940gat));
NR2X1 gate2305(.O (n746gat), .I1 (n2716gat), .I2 (n2723gat));
NR2X1 gate2306(.O (n360gat), .I1 (n2859gat), .I2 (n2727gat));
NR3X1 gate2307(.O (n710gat), .I1 (n714gat), .I2 (n715gat), .I3 (n716gat));
NR3X1 gate2308(.O (n711gat), .I1 (n714gat), .I2 (n717gat), .I3 (n718gat));
NR3X1 gate2309(.O (n712gat), .I1 (n719gat), .I2 (n715gat), .I3 (n718gat));
NR3X1 gate2310(.O (n713gat), .I1 (n719gat), .I2 (n717gat), .I3 (n716gat));
NR3X1 gate2311(.O (n729gat), .I1 (n733gat), .I2 (n734gat), .I3 (n735gat));
NR3X1 gate2312(.O (n730gat), .I1 (n733gat), .I2 (n736gat), .I3 (n737gat));
NR3X1 gate2313(.O (n731gat), .I1 (n738gat), .I2 (n734gat), .I3 (n737gat));
NR3X1 gate2314(.O (n732gat), .I1 (n738gat), .I2 (n736gat), .I3 (n735gat));
NR3X1 gate2315(.O (n494gat), .I1 (n498gat), .I2 (n499gat), .I3 (n500gat));
NR3X1 gate2316(.O (n495gat), .I1 (n498gat), .I2 (n501gat), .I3 (n502gat));
NR3X1 gate2317(.O (n496gat), .I1 (n503gat), .I2 (n499gat), .I3 (n502gat));
NR3X1 gate2318(.O (n497gat), .I1 (n503gat), .I2 (n501gat), .I3 (n500gat));
NR3X1 gate2319(.O (n505gat), .I1 (n509gat), .I2 (n510gat), .I3 (n511gat));
NR3X1 gate2320(.O (n506gat), .I1 (n509gat), .I2 (n512gat), .I3 (n513gat));
NR3X1 gate2321(.O (n507gat), .I1 (n514gat), .I2 (n510gat), .I3 (n513gat));
NR3X1 gate2322(.O (n508gat), .I1 (n514gat), .I2 (n512gat), .I3 (n511gat));
NR4X1 gate2323(.O (n564gat), .I1 (n3029gat), .I2 (n2863gat), .I3 (n2855gat), .I4 (n374gat));
NR3X1 gate2324(.O (n86gat), .I1 (n743gat), .I2 (n294gat), .I3 (n17gat));
NR2X1 gate2325(.O (n78gat), .I1 (n2784gat), .I2 (n79gat));
NR2X1 gate2326(.O (n767gat), .I1 (n219gat), .I2 (n2731gat));
NR2X1 gate2327(.O (n286gat), .I1 (n289gat), .I2 (n2723gat));
NR2X1 gate2328(.O (n287gat), .I1 (n289gat), .I2 (n2715gat));
NR2X1 gate2329(.O (n288gat), .I1 (n289gat), .I2 (n2726gat));
NR3X1 gate2330(.O (n181gat), .I1 (n286gat), .I2 (n179gat), .I3 (n188gat));
NR2X1 gate2331(.O (n182gat), .I1 (n72gat), .I2 (n2720gat));
NR2X1 gate2332(.O (n653gat), .I1 (n2718gat), .I2 (n111gat));
NR2X1 gate2333(.O (n867gat), .I1 (n219gat), .I2 (n2775gat));
NR2X1 gate2334(.O (n771gat), .I1 (n2838gat), .I2 (n111gat));
NR2X1 gate2335(.O (n964gat), .I1 (n111gat), .I2 (n2711gat));
NR2X1 gate2336(.O (n961gat), .I1 (n219gat), .I2 (n2734gat));
NR3X1 gate2337(.O (n804gat), .I1 (n808gat), .I2 (n809gat), .I3 (n810gat));
NR3X1 gate2338(.O (n805gat), .I1 (n808gat), .I2 (n811gat), .I3 (n812gat));
NR3X1 gate2339(.O (n806gat), .I1 (n813gat), .I2 (n809gat), .I3 (n812gat));
NR3X1 gate2340(.O (n807gat), .I1 (n813gat), .I2 (n811gat), .I3 (n810gat));
NR3X1 gate2341(.O (n587gat), .I1 (n591gat), .I2 (n592gat), .I3 (n593gat));
NR3X1 gate2342(.O (n588gat), .I1 (n591gat), .I2 (n594gat), .I3 (n595gat));
NR3X1 gate2343(.O (n589gat), .I1 (n596gat), .I2 (n592gat), .I3 (n595gat));
NR3X1 gate2344(.O (n590gat), .I1 (n596gat), .I2 (n594gat), .I3 (n593gat));
NR2X1 gate2345(.O (n447gat), .I1 (n2836gat), .I2 (n111gat));
NR2X1 gate2346(.O (n445gat), .I1 (n2778gat), .I2 (n219gat));
NR3X1 gate2347(.O (n687gat), .I1 (n691gat), .I2 (n692gat), .I3 (n693gat));
NR3X1 gate2348(.O (n688gat), .I1 (n691gat), .I2 (n694gat), .I3 (n695gat));
NR3X1 gate2349(.O (n689gat), .I1 (n696gat), .I2 (n692gat), .I3 (n695gat));
NR3X1 gate2350(.O (n690gat), .I1 (n696gat), .I2 (n694gat), .I3 (n693gat));
NR3X1 gate2351(.O (n568gat), .I1 (n572gat), .I2 (n573gat), .I3 (n574gat));
NR3X1 gate2352(.O (n569gat), .I1 (n572gat), .I2 (n575gat), .I3 (n576gat));
NR3X1 gate2353(.O (n570gat), .I1 (n577gat), .I2 (n573gat), .I3 (n576gat));
NR3X1 gate2354(.O (n571gat), .I1 (n577gat), .I2 (n575gat), .I3 (n574gat));
NR3X1 gate2355(.O (n187gat), .I1 (n189gat), .I2 (n287gat), .I3 (n188gat));
NR2X1 gate2356(.O (n197gat), .I1 (n194gat), .I2 (n297gat));
NR3X1 gate2357(.O (n15gat), .I1 (n637gat), .I2 (n17gat), .I3 (n293gat));
NR2X1 gate2358(.O (n22gat), .I1 (n92gat), .I2 (n21gat));
NR2X1 gate2359(.O (n93gat), .I1 (n197gat), .I2 (n22gat));
NR2X1 gate2360(.O (n769gat), .I1 (n93gat), .I2 (n2731gat));
NR3X1 gate2361(.O (n2534gat), .I1 (n2624gat), .I2 (n2489gat), .I3 (n2621gat));
NR3X1 gate2362(.O (n2430gat), .I1 (n2533gat), .I2 (n2486gat), .I3 (n2429gat));
NR2X1 gate2363(.O (n1606gat), .I1 (n3020gat), .I2 (n270gat));
NR2X1 gate2364(.O (n2239gat), .I1 (n2850gat), .I2 (n3019gat));
NR3X1 gate2365(.O (n1934gat), .I1 (n2470gat), .I2 (n1935gat), .I3 (n2239gat));
NR2X1 gate2366(.O (n1610gat), .I1 (n1698gat), .I2 (n1543gat));
NR2X1 gate2367(.O (n1692gat), .I1 (n1879gat), .I2 (n1762gat));
NR2X1 gate2368(.O (n2433gat), .I1 (n2432gat), .I2 (n2154gat));
NR3X1 gate2369(.O (n2531gat), .I1 (n2488gat), .I2 (n2625gat), .I3 (n2621gat));
NR3X1 gate2370(.O (n2480gat), .I1 (n2530gat), .I2 (n2482gat), .I3 (n2486gat));
NR2X1 gate2371(.O (n2427gat), .I1 (n2426gat), .I2 (n2153gat));
NR2X1 gate2372(.O (n2428gat), .I1 (n2433gat), .I2 (n2427gat));
NR2X1 gate2373(.O (n1778gat), .I1 (n3026gat), .I2 (n1779gat));
NR2X1 gate2374(.O (n1609gat), .I1 (n1503gat), .I2 (n3025gat));
NR2X1 gate2375(.O (n1702gat), .I1 (n3024gat), .I2 (n1615gat));
NR2X1 gate2376(.O (n1700gat), .I1 (n1701gat), .I2 (n3023gat));
NR4X1 gate2377(.O (n1604gat), .I1 (n1778gat), .I2 (n1609gat), .I3 (n1702gat), .I4 (n1700gat));
NR2X1 gate2378(.O (n1076gat), .I1 (n93gat), .I2 (n2775gat));
NR2X1 gate2379(.O (n766gat), .I1 (n93gat), .I2 (n2734gat));
NR3X1 gate2380(.O (n1185gat), .I1 (n1189gat), .I2 (n1190gat), .I3 (n1191gat));
NR3X1 gate2381(.O (n1186gat), .I1 (n1189gat), .I2 (n1192gat), .I3 (n1193gat));
NR3X1 gate2382(.O (n1187gat), .I1 (n1194gat), .I2 (n1190gat), .I3 (n1193gat));
NR3X1 gate2383(.O (n1188gat), .I1 (n1194gat), .I2 (n1192gat), .I3 (n1191gat));
NR2X1 gate2384(.O (n645gat), .I1 (n2792gat), .I2 (n93gat));
NR2X1 gate2385(.O (n646gat), .I1 (n93gat), .I2 (n2669gat));
NR2X1 gate2386(.O (n1383gat), .I1 (n1280gat), .I2 (n1225gat));
NR2X1 gate2387(.O (n1327gat), .I1 (n1281gat), .I2 (n1224gat));
NR2X1 gate2388(.O (n651gat), .I1 (n93gat), .I2 (n2778gat));
NR2X1 gate2389(.O (n652gat), .I1 (n2789gat), .I2 (n93gat));
NR2X1 gate2390(.O (n765gat), .I1 (n2781gat), .I2 (n93gat));
NR3X1 gate2391(.O (n1202gat), .I1 (n1206gat), .I2 (n1207gat), .I3 (n1208gat));
NR3X1 gate2392(.O (n1203gat), .I1 (n1206gat), .I2 (n1209gat), .I3 (n1210gat));
NR3X1 gate2393(.O (n1204gat), .I1 (n1211gat), .I2 (n1207gat), .I3 (n1210gat));
NR3X1 gate2394(.O (n1205gat), .I1 (n1211gat), .I2 (n1209gat), .I3 (n1208gat));
NR3X1 gate2395(.O (n1270gat), .I1 (n1274gat), .I2 (n1275gat), .I3 (n1276gat));
NR3X1 gate2396(.O (n1271gat), .I1 (n1274gat), .I2 (n1277gat), .I3 (n1278gat));
NR3X1 gate2397(.O (n1272gat), .I1 (n1279gat), .I2 (n1275gat), .I3 (n1278gat));
NR3X1 gate2398(.O (n1273gat), .I1 (n1279gat), .I2 (n1277gat), .I3 (n1276gat));
NR2X1 gate2399(.O (n763gat), .I1 (n2672gat), .I2 (n93gat));
NR2X1 gate2400(.O (n1287gat), .I1 (n1284gat), .I2 (n1195gat));
NR2X1 gate2401(.O (n1285gat), .I1 (n1196gat), .I2 (n1269gat));
NR2X1 gate2402(.O (n853gat), .I1 (n740gat), .I2 (n2148gat));
NR2X1 gate2403(.O (n793gat), .I1 (n2852gat), .I2 (n851gat));
NR2X1 gate2404(.O (n854gat), .I1 (n2148gat), .I2 (n374gat));
NR2X1 gate2405(.O (n556gat), .I1 (n2672gat), .I2 (n852gat));
NR2X1 gate2406(.O (n795gat), .I1 (n2731gat), .I2 (n852gat));
NR2X1 gate2407(.O (n656gat), .I1 (n851gat), .I2 (n2718gat));
NR2X1 gate2408(.O (n794gat), .I1 (n852gat), .I2 (n2775gat));
NR2X1 gate2409(.O (n773gat), .I1 (n851gat), .I2 (n2838gat));
NR2X1 gate2410(.O (n965gat), .I1 (n2711gat), .I2 (n851gat));
NR2X1 gate2411(.O (n960gat), .I1 (n2734gat), .I2 (n852gat));
NR3X1 gate2412(.O (n780gat), .I1 (n784gat), .I2 (n785gat), .I3 (n786gat));
NR3X1 gate2413(.O (n781gat), .I1 (n784gat), .I2 (n787gat), .I3 (n788gat));
NR3X1 gate2414(.O (n782gat), .I1 (n789gat), .I2 (n785gat), .I3 (n788gat));
NR3X1 gate2415(.O (n783gat), .I1 (n789gat), .I2 (n787gat), .I3 (n786gat));
NR2X1 gate2416(.O (n555gat), .I1 (n852gat), .I2 (n2792gat));
NR2X1 gate2417(.O (n450gat), .I1 (n851gat), .I2 (n2846gat));
NR2X1 gate2418(.O (n654gat), .I1 (n851gat), .I2 (n2844gat));
NR2X1 gate2419(.O (n557gat), .I1 (n2669gat), .I2 (n852gat));
NR2X1 gate2420(.O (n874gat), .I1 (n559gat), .I2 (n365gat));
NR2X1 gate2421(.O (n132gat), .I1 (n560gat), .I2 (n364gat));
NR2X1 gate2422(.O (n649gat), .I1 (n2778gat), .I2 (n852gat));
NR2X1 gate2423(.O (n449gat), .I1 (n2836gat), .I2 (n851gat));
NR2X1 gate2424(.O (n791gat), .I1 (n851gat), .I2 (n2840gat));
NR2X1 gate2425(.O (n650gat), .I1 (n852gat), .I2 (n2789gat));
NR2X1 gate2426(.O (n774gat), .I1 (n2842gat), .I2 (n851gat));
NR2X1 gate2427(.O (n764gat), .I1 (n852gat), .I2 (n2781gat));
NR3X1 gate2428(.O (n222gat), .I1 (n226gat), .I2 (n227gat), .I3 (n228gat));
NR3X1 gate2429(.O (n223gat), .I1 (n226gat), .I2 (n229gat), .I3 (n230gat));
NR3X1 gate2430(.O (n224gat), .I1 (n231gat), .I2 (n227gat), .I3 (n230gat));
NR3X1 gate2431(.O (n225gat), .I1 (n231gat), .I2 (n229gat), .I3 (n228gat));
NR3X1 gate2432(.O (n121gat), .I1 (n125gat), .I2 (n126gat), .I3 (n127gat));
NR3X1 gate2433(.O (n122gat), .I1 (n125gat), .I2 (n128gat), .I3 (n129gat));
NR3X1 gate2434(.O (n123gat), .I1 (n130gat), .I2 (n126gat), .I3 (n129gat));
NR3X1 gate2435(.O (n124gat), .I1 (n130gat), .I2 (n128gat), .I3 (n127gat));
NR2X1 gate2436(.O (n2460gat), .I1 (n666gat), .I2 (n120gat));
NR2X1 gate2437(.O (n2423gat), .I1 (n665gat), .I2 (n1601gat));
NR3X1 gate2438(.O (n2594gat), .I1 (n3017gat), .I2 (n2520gat), .I3 (n2597gat));
NR3X1 gate2439(.O (n2569gat), .I1 (n2573gat), .I2 (n2574gat), .I3 (n2575gat));
NR3X1 gate2440(.O (n2570gat), .I1 (n2573gat), .I2 (n2576gat), .I3 (n2577gat));
NR3X1 gate2441(.O (n2571gat), .I1 (n2578gat), .I2 (n2574gat), .I3 (n2577gat));
NR3X1 gate2442(.O (n2572gat), .I1 (n2578gat), .I2 (n2576gat), .I3 (n2575gat));
NR3X1 gate2443(.O (n2410gat), .I1 (n2414gat), .I2 (n2415gat), .I3 (n2416gat));
NR3X1 gate2444(.O (n2411gat), .I1 (n2414gat), .I2 (n2417gat), .I3 (n2418gat));
NR3X1 gate2445(.O (n2412gat), .I1 (n2419gat), .I2 (n2415gat), .I3 (n2418gat));
NR3X1 gate2446(.O (n2413gat), .I1 (n2419gat), .I2 (n2417gat), .I3 (n2416gat));
NR2X1 gate2447(.O (n2583gat), .I1 (n2582gat), .I2 (n2585gat));
NR2X1 gate2448(.O (n2580gat), .I1 (n2582gat), .I2 (n2583gat));
NR2X1 gate2449(.O (n2581gat), .I1 (n2583gat), .I2 (n2585gat));
NR2X1 gate2450(.O (n2567gat), .I1 (n2493gat), .I2 (n2388gat));
NR2X1 gate2451(.O (n2499gat), .I1 (n2389gat), .I2 (n2494gat));
NR2X1 gate2452(.O (n299gat), .I1 (n2268gat), .I2 (n2338gat));
NR2X1 gate2453(.O (n207gat), .I1 (n2337gat), .I2 (n2269gat));
NR2X1 gate2454(.O (n2650gat), .I1 (n2649gat), .I2 (n2652gat));
NR2X1 gate2455(.O (n2647gat), .I1 (n2649gat), .I2 (n2650gat));
NR2X1 gate2456(.O (n2648gat), .I1 (n2650gat), .I2 (n2652gat));
NR3X1 gate2457(.O (n2602gat), .I1 (n2606gat), .I2 (n2607gat), .I3 (n2608gat));
NR3X1 gate2458(.O (n2603gat), .I1 (n2606gat), .I2 (n2609gat), .I3 (n2610gat));
NR3X1 gate2459(.O (n2604gat), .I1 (n2611gat), .I2 (n2607gat), .I3 (n2610gat));
NR3X1 gate2460(.O (n2605gat), .I1 (n2611gat), .I2 (n2609gat), .I3 (n2608gat));
NR3X1 gate2461(.O (n2546gat), .I1 (n2550gat), .I2 (n2551gat), .I3 (n2552gat));
NR3X1 gate2462(.O (n2547gat), .I1 (n2550gat), .I2 (n2553gat), .I3 (n2554gat));
NR3X1 gate2463(.O (n2548gat), .I1 (n2555gat), .I2 (n2551gat), .I3 (n2554gat));
NR3X1 gate2464(.O (n2549gat), .I1 (n2555gat), .I2 (n2553gat), .I3 (n2552gat));
NR2X1 gate2465(.O (n2617gat), .I1 (n2616gat), .I2 (n2619gat));
NR2X1 gate2466(.O (n2614gat), .I1 (n2616gat), .I2 (n2617gat));
NR2X1 gate2467(.O (n2615gat), .I1 (n2617gat), .I2 (n2619gat));
NR4X1 gate2468(.O (n2655gat), .I1 (n2508gat), .I2 (n2656gat), .I3 (n2500gat), .I4 (n2504gat));
NR3X1 gate2469(.O (n2293gat), .I1 (n2353gat), .I2 (n2284gat), .I3 (n2443gat));
NR2X1 gate2470(.O (n2219gat), .I1 (n2354gat), .I2 (n2214gat));
NR2X1 gate2471(.O (n1529gat), .I1 (n1528gat), .I2 (n1523gat));
NR2X1 gate2472(.O (n1704gat), .I1 (n3027gat), .I2 (n1706gat));
NR2X1 gate2473(.O (n2461gat), .I1 (n120gat), .I2 (n2666gat));
NR2X1 gate2474(.O (n2421gat), .I1 (n1601gat), .I2 (n1704gat));
NR2X1 gate2475(.O (n1598gat), .I1 (n1592gat), .I2 (n2422gat));
NR2X1 gate2476(.O (n2218gat), .I1 (n2214gat), .I2 (n2290gat));
NR3X1 gate2477(.O (n2358gat), .I1 (n2285gat), .I2 (n2356gat), .I3 (n2355gat));
NR2X1 gate2478(.O (n1415gat), .I1 (n2081gat), .I2 (n2359gat));
NR2X1 gate2479(.O (n1153gat), .I1 (n1414gat), .I2 (n566gat));
NR3X1 gate2480(.O (n2292gat), .I1 (n2443gat), .I2 (n2284gat), .I3 (n2285gat));
NR2X1 gate2481(.O (n1416gat), .I1 (n2081gat), .I2 (n1480gat));
NR2X1 gate2482(.O (n1151gat), .I1 (n1301gat), .I2 (n1150gat));
NR3X1 gate2483(.O (n2306gat), .I1 (n2356gat), .I2 (n2284gat), .I3 (n2285gat));
NR2X1 gate2484(.O (n1481gat), .I1 (n2081gat), .I2 (n2011gat));
NR2X1 gate2485(.O (n982gat), .I1 (n873gat), .I2 (n1478gat));
NR3X1 gate2486(.O (n2357gat), .I1 (n2285gat), .I2 (n2355gat), .I3 (n2443gat));
NR2X1 gate2487(.O (n1347gat), .I1 (n2081gat), .I2 (n1410gat));
NR2X1 gate2488(.O (n877gat), .I1 (n875gat), .I2 (n876gat));
NR2X1 gate2489(.O (n1484gat), .I1 (n2081gat), .I2 (n1528gat));
NR2X1 gate2490(.O (n1159gat), .I1 (n1160gat), .I2 (n1084gat));
NR3X1 gate2491(.O (n2363gat), .I1 (n2353gat), .I2 (n2356gat), .I3 (n2355gat));
NR2X1 gate2492(.O (n1483gat), .I1 (n2081gat), .I2 (n1482gat));
NR2X1 gate2493(.O (n1158gat), .I1 (n983gat), .I2 (n1157gat));
NR3X1 gate2494(.O (n2364gat), .I1 (n2353gat), .I2 (n2284gat), .I3 (n2356gat));
NR2X1 gate2495(.O (n1308gat), .I1 (n2081gat), .I2 (n1530gat));
NR2X1 gate2496(.O (n1156gat), .I1 (n985gat), .I2 (n1307gat));
NR3X1 gate2497(.O (n2291gat), .I1 (n2353gat), .I2 (n2355gat), .I3 (n2443gat));
NR2X1 gate2498(.O (n1349gat), .I1 (n1479gat), .I2 (n2081gat));
NR2X1 gate2499(.O (n1155gat), .I1 (n1085gat), .I2 (n1348gat));
NR3X1 gate2500(.O (n1154gat), .I1 (n1598gat), .I2 (n2930gat), .I3 (n2957gat));
NR2X1 gate2501(.O (n1703gat), .I1 (n1705gat), .I2 (n3028gat));
NR2X1 gate2502(.O (n1608gat), .I1 (n1704gat), .I2 (n1703gat));
NR2X1 gate2503(.O (n1411gat), .I1 (n1154gat), .I2 (n1608gat));
NR2X1 gate2504(.O (n2223gat), .I1 (n2354gat), .I2 (n2217gat));
NR2X1 gate2505(.O (n1438gat), .I1 (n1591gat), .I2 (n1480gat));
NR2X1 gate2506(.O (n1625gat), .I1 (n3021gat), .I2 (n1628gat));
NR2X1 gate2507(.O (n1626gat), .I1 (n1627gat), .I2 (n3022gat));
NR3X1 gate2508(.O (n1831gat), .I1 (n1832gat), .I2 (n1765gat), .I3 (n1878gat));
NR2X1 gate2509(.O (n1443gat), .I1 (n1442gat), .I2 (n706gat));
NR2X1 gate2510(.O (n1325gat), .I1 (n1444gat), .I2 (n164gat));
NR2X1 gate2511(.O (n1441gat), .I1 (n1437gat), .I2 (n1378gat));
NR2X1 gate2512(.O (n1321gat), .I1 (n1442gat), .I2 (n837gat));
NR2X1 gate2513(.O (n1320gat), .I1 (n1444gat), .I2 (n278gat));
NR2X1 gate2514(.O (n1486gat), .I1 (n1482gat), .I2 (n1591gat));
NR2X1 gate2515(.O (n1440gat), .I1 (n1322gat), .I2 (n1439gat));
NR2X1 gate2516(.O (n1426gat), .I1 (n2011gat), .I2 (n1591gat));
NR2X1 gate2517(.O (n1368gat), .I1 (n1442gat), .I2 (n613gat));
NR2X1 gate2518(.O (n1258gat), .I1 (n274gat), .I2 (n1444gat));
NR2X1 gate2519(.O (n1371gat), .I1 (n1370gat), .I2 (n1369gat));
NR2X1 gate2520(.O (n1365gat), .I1 (n1479gat), .I2 (n1591gat));
NR2X1 gate2521(.O (n1373gat), .I1 (n833gat), .I2 (n1442gat));
NR2X1 gate2522(.O (n1372gat), .I1 (n282gat), .I2 (n1444gat));
NR2X1 gate2523(.O (n1367gat), .I1 (n1366gat), .I2 (n1374gat));
NR2X1 gate2524(.O (n2220gat), .I1 (n2290gat), .I2 (n2217gat));
NR2X1 gate2525(.O (n1423gat), .I1 (n2162gat), .I2 (n1530gat));
NR2X1 gate2526(.O (n1498gat), .I1 (n1609gat), .I2 (n1427gat));
NR2X1 gate2527(.O (n1504gat), .I1 (n1450gat), .I2 (n1498gat));
NR2X1 gate2528(.O (n1607gat), .I1 (n2082gat), .I2 (n1609gat));
NR2X1 gate2529(.O (n1494gat), .I1 (n1528gat), .I2 (n2162gat));
NR2X1 gate2530(.O (n1502gat), .I1 (n1607gat), .I2 (n1449gat));
NR2X1 gate2531(.O (n1250gat), .I1 (n1603gat), .I2 (n815gat));
NR2X1 gate2532(.O (n1103gat), .I1 (n956gat), .I2 (n1590gat));
NR2X1 gate2533(.O (n1417gat), .I1 (n2162gat), .I2 (n1480gat));
NR2X1 gate2534(.O (n1352gat), .I1 (n1248gat), .I2 (n1418gat));
NR2X1 gate2535(.O (n1304gat), .I1 (n1590gat), .I2 (n1067gat));
NR2X1 gate2536(.O (n1249gat), .I1 (n679gat), .I2 (n1603gat));
NR2X1 gate2537(.O (n1419gat), .I1 (n2162gat), .I2 (n1479gat));
NR2X1 gate2538(.O (n1351gat), .I1 (n1306gat), .I2 (n1353gat));
NR2X1 gate2539(.O (n1246gat), .I1 (n864gat), .I2 (n1590gat));
NR2X1 gate2540(.O (n1161gat), .I1 (n583gat), .I2 (n1603gat));
NR2X1 gate2541(.O (n1422gat), .I1 (n2011gat), .I2 (n2162gat));
NR2X1 gate2542(.O (n1303gat), .I1 (n1247gat), .I2 (n1355gat));
NR2X1 gate2543(.O (n1291gat), .I1 (n1603gat), .I2 (n579gat));
NR2X1 gate2544(.O (n1245gat), .I1 (n1590gat), .I2 (n860gat));
NR2X1 gate2545(.O (n1485gat), .I1 (n1482gat), .I2 (n2162gat));
NR2X1 gate2546(.O (n1302gat), .I1 (n1300gat), .I2 (n1487gat));
NR2X1 gate2547(.O (n1163gat), .I1 (n882gat), .I2 (n1603gat));
NR2X1 gate2548(.O (n1102gat), .I1 (n1297gat), .I2 (n1590gat));
NR2X1 gate2549(.O (n1354gat), .I1 (n1591gat), .I2 (n1530gat));
NR2X1 gate2550(.O (n1360gat), .I1 (n1164gat), .I2 (n1356gat));
NR2X1 gate2551(.O (n1435gat), .I1 (n1591gat), .I2 (n1528gat));
NR2X1 gate2552(.O (n1101gat), .I1 (n1590gat), .I2 (n1293gat));
NR2X1 gate2553(.O (n996gat), .I1 (n1603gat), .I2 (n823gat));
NR2X1 gate2554(.O (n1359gat), .I1 (n1436gat), .I2 (n1106gat));
NR2X1 gate2555(.O (n1421gat), .I1 (n2162gat), .I2 (n2359gat));
NR2X1 gate2556(.O (n1104gat), .I1 (n1079gat), .I2 (n1590gat));
NR2X1 gate2557(.O (n887gat), .I1 (n1603gat), .I2 (n683gat));
NR2X1 gate2558(.O (n1358gat), .I1 (n1425gat), .I2 (n1105gat));
NR2X1 gate2559(.O (n1420gat), .I1 (n1410gat), .I2 (n2162gat));
NR2X1 gate2560(.O (n1305gat), .I1 (n1147gat), .I2 (n1590gat));
NR2X1 gate2561(.O (n1162gat), .I1 (n698gat), .I2 (n1603gat));
NR2X1 gate2562(.O (n1357gat), .I1 (n1424gat), .I2 (n1309gat));
NR4X1 gate2563(.O (n1428gat), .I1 (n2978gat), .I2 (n2982gat), .I3 (n2973gat), .I4 (n2977gat));
NR2X1 gate2564(.O (n1794gat), .I1 (n1673gat), .I2 (n1719gat));
NR2X1 gate2565(.O (n1796gat), .I1 (n1858gat), .I2 (n1635gat));
NR2X1 gate2566(.O (n1792gat), .I1 (n1794gat), .I2 (n1796gat));
NR3X1 gate2567(.O (n1865gat), .I1 (n1989gat), .I2 (n1918gat), .I3 (n1986gat));
NR3X1 gate2568(.O (n1861gat), .I1 (n1866gat), .I2 (n2216gat), .I3 (n1988gat));
NR2X1 gate2569(.O (n1793gat), .I1 (n1792gat), .I2 (n1735gat));
NR2X1 gate2570(.O (n1406gat), .I1 (n1428gat), .I2 (n1387gat));
NR3X1 gate2571(.O (n1780gat), .I1 (n1777gat), .I2 (n1625gat), .I3 (n1626gat));
NR2X1 gate2572(.O (n2016gat), .I1 (n2019gat), .I2 (n1878gat));
NR2X1 gate2573(.O (n2664gat), .I1 (n2850gat), .I2 (n3018gat));
NR3X1 gate2574(.O (n1666gat), .I1 (n1986gat), .I2 (n2212gat), .I3 (n1991gat));
NR3X1 gate2575(.O (n1578gat), .I1 (n2152gat), .I2 (n2351gat), .I3 (n1665gat));
NR2X1 gate2576(.O (n1516gat), .I1 (n1551gat), .I2 (n1517gat));
NR3X1 gate2577(.O (n1864gat), .I1 (n1858gat), .I2 (n1495gat), .I3 (n2090gat));
NR2X1 gate2578(.O (n1565gat), .I1 (n1735gat), .I2 (n1552gat));
NR2X1 gate2579(.O (n1921gat), .I1 (n1738gat), .I2 (n1673gat));
NR2X1 gate2580(.O (n1798gat), .I1 (n1739gat), .I2 (n1673gat));
NR3X1 gate2581(.O (n1920gat), .I1 (n1864gat), .I2 (n1921gat), .I3 (n1798gat));
NR2X1 gate2582(.O (n1926gat), .I1 (n1925gat), .I2 (n1635gat));
NR2X1 gate2583(.O (n1916gat), .I1 (n1917gat), .I2 (n1859gat));
NR2X1 gate2584(.O (n1994gat), .I1 (n1719gat), .I2 (n1922gat));
NR2X1 gate2585(.O (n1924gat), .I1 (n1743gat), .I2 (n1923gat));
NR4X1 gate2586(.O (n2078gat), .I1 (n1926gat), .I2 (n1916gat), .I3 (n1994gat), .I4 (n1924gat));
NR2X1 gate2587(.O (n1690gat), .I1 (n1700gat), .I2 (n1702gat));
NR3X1 gate2588(.O (n1660gat), .I1 (n1918gat), .I2 (n1986gat), .I3 (n2212gat));
NR3X1 gate2589(.O (n1576gat), .I1 (n2351gat), .I2 (n1988gat), .I3 (n1661gat));
NR2X1 gate2590(.O (n1733gat), .I1 (n1673gat), .I2 (n1572gat));
NR3X1 gate2591(.O (n1582gat), .I1 (n2283gat), .I2 (n1991gat), .I3 (n2212gat));
NR3X1 gate2592(.O (n1577gat), .I1 (n1520gat), .I2 (n2351gat), .I3 (n1988gat));
NR2X1 gate2593(.O (n1581gat), .I1 (n1858gat), .I2 (n1580gat));
NR3X1 gate2594(.O (n2129gat), .I1 (n2189gat), .I2 (n2134gat), .I3 (n2261gat));
NR4X1 gate2595(.O (n2079gat), .I1 (n2078gat), .I2 (n2178gat), .I3 (n1990gat), .I4 (n2128gat));
NR4X1 gate2596(.O (n1695gat), .I1 (n1609gat), .I2 (n1778gat), .I3 (n1704gat), .I4 (n1703gat));
NR3X1 gate2597(.O (n2073gat), .I1 (n2078gat), .I2 (n1990gat), .I3 (n2181gat));
NR2X1 gate2598(.O (n1696gat), .I1 (n1707gat), .I2 (n1698gat));
NR2X1 gate2599(.O (n1758gat), .I1 (n1311gat), .I2 (n1773gat));
NR3X1 gate2600(.O (n1574gat), .I1 (n1719gat), .I2 (n1673gat), .I3 (n1444gat));
NR3X1 gate2601(.O (n1573gat), .I1 (n1444gat), .I2 (n1858gat), .I3 (n1635gat));
NR2X1 gate2602(.O (n1521gat), .I1 (n2283gat), .I2 (n1991gat));
NR2X1 gate2603(.O (n1737gat), .I1 (n2212gat), .I2 (n2152gat));
NR3X1 gate2604(.O (n1732gat), .I1 (n1515gat), .I2 (n1736gat), .I3 (n1658gat));
NR3X1 gate2605(.O (n1723gat), .I1 (n1659gat), .I2 (n1722gat), .I3 (n1724gat));
NR2X1 gate2606(.O (n1663gat), .I1 (n1986gat), .I2 (n1918gat));
NR3X1 gate2607(.O (n1655gat), .I1 (n1736gat), .I2 (n1662gat), .I3 (n1658gat));
NR3X1 gate2608(.O (n1647gat), .I1 (n1656gat), .I2 (n1659gat), .I3 (n1554gat));
NR2X1 gate2609(.O (n1667gat), .I1 (n1991gat), .I2 (n1986gat));
NR3X1 gate2610(.O (n1570gat), .I1 (n1736gat), .I2 (n1658gat), .I3 (n1670gat));
NR3X1 gate2611(.O (n1646gat), .I1 (n1569gat), .I2 (n1659gat), .I3 (n1566gat));
NR2X1 gate2612(.O (n1575gat), .I1 (n1918gat), .I2 (n2283gat));
NR3X1 gate2613(.O (n1728gat), .I1 (n1568gat), .I2 (n1736gat), .I3 (n1658gat));
NR3X1 gate2614(.O (n1650gat), .I1 (n1727gat), .I2 (n1659gat), .I3 (n1640gat));
NR2X1 gate2615(.O (n1801gat), .I1 (n2152gat), .I2 (n1989gat));
NR3X1 gate2616(.O (n1731gat), .I1 (n1658gat), .I2 (n1515gat), .I3 (n1797gat));
NR3X1 gate2617(.O (n1649gat), .I1 (n1560gat), .I2 (n1659gat), .I3 (n1730gat));
NR3X1 gate2618(.O (n1571gat), .I1 (n1670gat), .I2 (n1658gat), .I3 (n1797gat));
NR3X1 gate2619(.O (n1563gat), .I1 (n1561gat), .I2 (n1562gat), .I3 (n1659gat));
NR2X1 gate2620(.O (n1734gat), .I1 (n1988gat), .I2 (n2212gat));
NR3X1 gate2621(.O (n1669gat), .I1 (n1668gat), .I2 (n1742gat), .I3 (n1670gat));
NR2X1 gate2622(.O (n1654gat), .I1 (n1671gat), .I2 (n1659gat));
NR3X1 gate2623(.O (n1657gat), .I1 (n1662gat), .I2 (n1797gat), .I3 (n1658gat));
NR3X1 gate2624(.O (n1653gat), .I1 (n1651gat), .I2 (n1652gat), .I3 (n1659gat));
NR3X1 gate2625(.O (n1729gat), .I1 (n1658gat), .I2 (n1797gat), .I3 (n1568gat));
NR3X1 gate2626(.O (n1644gat), .I1 (n1643gat), .I2 (n1648gat), .I3 (n1659gat));
NR3X1 gate2627(.O (n1726gat), .I1 (n2992gat), .I2 (n2986gat), .I3 (n2991gat));
NR2X1 gate2628(.O (n1929gat), .I1 (n1758gat), .I2 (n1790gat));
NR3X1 gate2629(.O (n2009gat), .I1 (n2016gat), .I2 (n2664gat), .I3 (n2004gat));
NR3X1 gate2630(.O (n1413gat), .I1 (n1869gat), .I2 (n672gat), .I3 (n2591gat));
NR2X1 gate2631(.O (n1636gat), .I1 (n1584gat), .I2 (n1718gat));
NR2X1 gate2632(.O (n1401gat), .I1 (n1584gat), .I2 (n1590gat));
NR3X1 gate2633(.O (n1408gat), .I1 (n1507gat), .I2 (n1396gat), .I3 (n1393gat));
NR2X1 gate2634(.O (n1476gat), .I1 (n1858gat), .I2 (n1590gat));
NR3X1 gate2635(.O (n1407gat), .I1 (n1393gat), .I2 (n1409gat), .I3 (n1677gat));
NR3X1 gate2636(.O (n1412gat), .I1 (n1411gat), .I2 (n1406gat), .I3 (n2981gat));
NR3X1 gate2637(.O (n2663gat), .I1 (n2586gat), .I2 (n2660gat), .I3 (n2307gat));
NR2X1 gate2638(.O (n2662gat), .I1 (n2660gat), .I2 (n2586gat));
NR2X1 gate2639(.O (n2238gat), .I1 (n2448gat), .I2 (n2444gat));
NR3X1 gate2640(.O (n87gat), .I1 (n743gat), .I2 (n17gat), .I3 (n293gat));
NR2X1 gate2641(.O (n200gat), .I1 (n199gat), .I2 (n92gat));
NR3X1 gate2642(.O (n184gat), .I1 (n189gat), .I2 (n188gat), .I3 (n179gat));
NR2X1 gate2643(.O (n196gat), .I1 (n297gat), .I2 (n195gat));
NR2X1 gate2644(.O (n204gat), .I1 (n200gat), .I2 (n196gat));
NR4X1 gate2645(.O (n2163gat), .I1 (n1790gat), .I2 (n1310gat), .I3 (n2664gat), .I4 (n2168gat));
NR2X1 gate2646(.O (n2258gat), .I1 (n2260gat), .I2 (n2189gat));
NR2X1 gate2647(.O (n2255gat), .I1 (n2261gat), .I2 (n2188gat));
NR3X1 gate2648(.O (n2015gat), .I1 (n2039gat), .I2 (n1774gat), .I3 (n1315gat));
NR2X1 gate2649(.O (n2017gat), .I1 (n1790gat), .I2 (n2016gat));
NR2X1 gate2650(.O (n2018gat), .I1 (n2016gat), .I2 (n2097gat));
NR4X1 gate2651(.O (n2014gat), .I1 (n2035gat), .I2 (n2093gat), .I3 (n2018gat), .I4 (n2664gat));
NR2X1 gate2652(.O (n2194gat), .I1 (n2187gat), .I2 (n1855gat));
NR2X1 gate2653(.O (n2192gat), .I1 (n2184gat), .I2 (n1855gat));
NR2X1 gate2654(.O (n2185gat), .I1 (n2261gat), .I2 (n2189gat));
NR2X1 gate2655(.O (n2132gat), .I1 (n2133gat), .I2 (n2131gat));
NR2X1 gate2656(.O (n2130gat), .I1 (n2134gat), .I2 (n2185gat));
NR2X1 gate2657(.O (n2057gat), .I1 (n2049gat), .I2 (n1855gat));
NR2X1 gate2658(.O (n2250gat), .I1 (n2248gat), .I2 (n2264gat));
NR2X1 gate2659(.O (n2249gat), .I1 (n2265gat), .I2 (n3006gat));
NR2X1 gate2660(.O (n2329gat), .I1 (n1855gat), .I2 (n3007gat));
NR2X1 gate2661(.O (n1958gat), .I1 (n1963gat), .I2 (n1886gat));
NR3X1 gate2662(.O (n1895gat), .I1 (n1845gat), .I2 (n1891gat), .I3 (n1968gat));
NR2X1 gate2663(.O (n1710gat), .I1 (n1709gat), .I2 (n1629gat));
NR2X1 gate2664(.O (n1630gat), .I1 (n1895gat), .I2 (n1631gat));
NR2X1 gate2665(.O (n2195gat), .I1 (n2200gat), .I2 (n1855gat));
NR2X1 gate2666(.O (n2556gat), .I1 (n1711gat), .I2 (n2437gat));
NR2X1 gate2667(.O (n2539gat), .I1 (n2048gat), .I2 (n2437gat));
NR3X1 gate2668(.O (n1894gat), .I1 (n1968gat), .I2 (n1891gat), .I3 (n1969gat));
NR2X1 gate2669(.O (n1847gat), .I1 (n1958gat), .I2 (n1845gat));
NR2X1 gate2670(.O (n1846gat), .I1 (n1845gat), .I2 (n1893gat));
NR2X1 gate2671(.O (n2436gat), .I1 (n2437gat), .I2 (n1892gat));
NR2X1 gate2672(.O (n2055gat), .I1 (n1891gat), .I2 (n1958gat));
NR2X1 gate2673(.O (n1967gat), .I1 (n1893gat), .I2 (n1968gat));
NR2X1 gate2674(.O (n2387gat), .I1 (n2056gat), .I2 (n2437gat));
NR2X1 gate2675(.O (n1959gat), .I1 (n1956gat), .I2 (n1963gat));
NR2X1 gate2676(.O (n1957gat), .I1 (n1886gat), .I2 (n1887gat));
NR2X1 gate2677(.O (n2330gat), .I1 (n2437gat), .I2 (n1961gat));
NR2X1 gate2678(.O (n2147gat), .I1 (n2988gat), .I2 (n1855gat));
NR2X1 gate2679(.O (n2498gat), .I1 (n2199gat), .I2 (n2328gat));
NR2X1 gate2680(.O (n2193gat), .I1 (n2393gat), .I2 (n2439gat));
NR2X1 gate2681(.O (n2211gat), .I1 (n2193gat), .I2 (n2402gat));
NR2X1 gate2682(.O (n2210gat), .I1 (n2401gat), .I2 (n2151gat));
NR2X1 gate2683(.O (n2396gat), .I1 (n2199gat), .I2 (n2209gat));
NR2X1 gate2684(.O (n2053gat), .I1 (n2393gat), .I2 (n2438gat));
NR2X1 gate2685(.O (n1964gat), .I1 (n2392gat), .I2 (n2439gat));
NR2X1 gate2686(.O (n2198gat), .I1 (n2199gat), .I2 (n2058gat));
NR3X1 gate2687(.O (n2215gat), .I1 (n2346gat), .I2 (n2151gat), .I3 (n2402gat));
NR2X1 gate2688(.O (n2350gat), .I1 (n2405gat), .I2 (n2349gat));
NR2X1 gate2689(.O (n2282gat), .I1 (n2406gat), .I2 (n2215gat));
NR2X1 gate2690(.O (n2197gat), .I1 (n2199gat), .I2 (n2281gat));
NR3X1 gate2691(.O (n2213gat), .I1 (n2402gat), .I2 (n2151gat), .I3 (n2345gat));
NR2X1 gate2692(.O (n2150gat), .I1 (n2401gat), .I2 (n2346gat));
NR2X1 gate2693(.O (n2149gat), .I1 (n2193gat), .I2 (n2346gat));
NR2X1 gate2694(.O (n2196gat), .I1 (n2199gat), .I2 (n2146gat));
NR3X1 gate2695(.O (n1882gat), .I1 (n2124gat), .I2 (n2115gat), .I3 (n2239gat));
NR2X1 gate2696(.O (n1962gat), .I1 (n1963gat), .I2 (n1893gat));
NR2X1 gate2697(.O (n1896gat), .I1 (n2995gat), .I2 (n1895gat));
NR2X1 gate2698(.O (n1972gat), .I1 (n1974gat), .I2 (n1970gat));
NR2X1 gate2699(.O (n1971gat), .I1 (n1896gat), .I2 (n1973gat));
NR2X1 gate2700(.O (n2559gat), .I1 (n2999gat), .I2 (n2437gat));
NR2X1 gate2701(.O (n2331gat), .I1 (n2393gat), .I2 (n2401gat));
NR2X1 gate2702(.O (n2352gat), .I1 (n3011gat), .I2 (n2215gat));
NR2X1 gate2703(.O (n2566gat), .I1 (n2643gat), .I2 (n2564gat));
NR2X1 gate2704(.O (n2565gat), .I1 (n2352gat), .I2 (n2642gat));
NR2X1 gate2705(.O (n2637gat), .I1 (n3015gat), .I2 (n2199gat));
NR3X1 gate2706(.O (n84gat), .I1 (n296gat), .I2 (n17gat), .I3 (n294gat));
NR2X1 gate2707(.O (n89gat), .I1 (n88gat), .I2 (n2784gat));
NR2X1 gate2708(.O (n110gat), .I1 (n182gat), .I2 (n89gat));
NR2X1 gate2709(.O (n1074gat), .I1 (n2775gat), .I2 (n110gat));
NR3X1 gate2710(.O (n141gat), .I1 (n155gat), .I2 (n253gat), .I3 (n150gat));
NR2X1 gate2711(.O (n38gat), .I1 (n151gat), .I2 (n233gat));
NR2X1 gate2712(.O (n37gat), .I1 (n151gat), .I2 (n154gat));
NR2X1 gate2713(.O (n872gat), .I1 (n375gat), .I2 (n800gat));
NR2X1 gate2714(.O (n234gat), .I1 (n155gat), .I2 (n233gat));
NR2X1 gate2715(.O (n137gat), .I1 (n154gat), .I2 (n253gat));
NR2X1 gate2716(.O (n378gat), .I1 (n375gat), .I2 (n235gat));
NR2X1 gate2717(.O (n377gat), .I1 (n110gat), .I2 (n2778gat));
NR2X1 gate2718(.O (n869gat), .I1 (n219gat), .I2 (n2792gat));
NR2X1 gate2719(.O (n212gat), .I1 (n182gat), .I2 (n78gat));
NR3X1 gate2720(.O (n250gat), .I1 (n329gat), .I2 (n387gat), .I3 (n334gat));
NR2X1 gate2721(.O (n249gat), .I1 (n386gat), .I2 (n330gat));
NR2X1 gate2722(.O (n248gat), .I1 (n330gat), .I2 (n1490gat));
NR2X1 gate2723(.O (n453gat), .I1 (n372gat), .I2 (n452gat));
NR2X1 gate2724(.O (n448gat), .I1 (n111gat), .I2 (n2846gat));
NR2X1 gate2725(.O (n974gat), .I1 (n2844gat), .I2 (n111gat));
NR2X1 gate2726(.O (n251gat), .I1 (n1490gat), .I2 (n387gat));
NR2X1 gate2727(.O (n244gat), .I1 (n334gat), .I2 (n386gat));
NR2X1 gate2728(.O (n973gat), .I1 (n372gat), .I2 (n333gat));
NR2X1 gate2729(.O (n870gat), .I1 (n2669gat), .I2 (n219gat));
NR2X1 gate2730(.O (n975gat), .I1 (n111gat), .I2 (n2852gat));
NR3X1 gate2731(.O (n246gat), .I1 (n330gat), .I2 (n325gat), .I3 (n334gat));
NR2X1 gate2732(.O (n245gat), .I1 (n386gat), .I2 (n334gat));
NR2X1 gate2733(.O (n460gat), .I1 (n462gat), .I2 (n2884gat));
NR2X1 gate2734(.O (n459gat), .I1 (n457gat), .I2 (n461gat));
NR2X1 gate2735(.O (n972gat), .I1 (n372gat), .I2 (n458gat));
NR2X1 gate2736(.O (n969gat), .I1 (n219gat), .I2 (n2672gat));
NR2X1 gate2737(.O (n971gat), .I1 (n111gat), .I2 (n2840gat));
NR3X1 gate2738(.O (n247gat), .I1 (n334gat), .I2 (n387gat), .I3 (n330gat));
NR2X1 gate2739(.O (n145gat), .I1 (n144gat), .I2 (n325gat));
NR2X1 gate2740(.O (n143gat), .I1 (n326gat), .I2 (n247gat));
NR2X1 gate2741(.O (n970gat), .I1 (n372gat), .I2 (n878gat));
NR2X1 gate2742(.O (n968gat), .I1 (n2789gat), .I2 (n219gat));
NR2X1 gate2743(.O (n772gat), .I1 (n111gat), .I2 (n2842gat));
NR3X1 gate2744(.O (n142gat), .I1 (n382gat), .I2 (n326gat), .I3 (n144gat));
NR2X1 gate2745(.O (n40gat), .I1 (n325gat), .I2 (n383gat));
NR2X1 gate2746(.O (n39gat), .I1 (n383gat), .I2 (n247gat));
NR2X1 gate2747(.O (n451gat), .I1 (n134gat), .I2 (n372gat));
NR2X1 gate2748(.O (n446gat), .I1 (n219gat), .I2 (n2781gat));
NR3X1 gate2749(.O (n139gat), .I1 (n253gat), .I2 (n151gat), .I3 (n254gat));
NR2X1 gate2750(.O (n136gat), .I1 (n253gat), .I2 (n154gat));
NR2X1 gate2751(.O (n391gat), .I1 (n252gat), .I2 (n468gat));
NR2X1 gate2752(.O (n390gat), .I1 (n469gat), .I2 (n2877gat));
NR2X1 gate2753(.O (n1083gat), .I1 (n381gat), .I2 (n375gat));
NR2X1 gate2754(.O (n1077gat), .I1 (n110gat), .I2 (n2672gat));
NR3X1 gate2755(.O (n140gat), .I1 (n151gat), .I2 (n253gat), .I3 (n155gat));
NR2X1 gate2756(.O (n242gat), .I1 (n254gat), .I2 (n241gat));
NR2X1 gate2757(.O (n240gat), .I1 (n255gat), .I2 (n140gat));
NR2X1 gate2758(.O (n871gat), .I1 (n802gat), .I2 (n375gat));
NR2X1 gate2759(.O (n797gat), .I1 (n110gat), .I2 (n2734gat));
NR3X1 gate2760(.O (n324gat), .I1 (n255gat), .I2 (n146gat), .I3 (n241gat));
NR2X1 gate2761(.O (n238gat), .I1 (n147gat), .I2 (n254gat));
NR2X1 gate2762(.O (n237gat), .I1 (n140gat), .I2 (n147gat));
NR2X1 gate2763(.O (n1082gat), .I1 (n375gat), .I2 (n380gat));
NR2X1 gate2764(.O (n796gat), .I1 (n2731gat), .I2 (n110gat));
NR3X1 gate2765(.O (n85gat), .I1 (n17gat), .I2 (n294gat), .I3 (n637gat));
NR3X1 gate2766(.O (n180gat), .I1 (n286gat), .I2 (n188gat), .I3 (n287gat));
NR2X1 gate2767(.O (n68gat), .I1 (n85gat), .I2 (n180gat));
NR3X1 gate2768(.O (n186gat), .I1 (n189gat), .I2 (n287gat), .I3 (n288gat));
NR2X1 gate2769(.O (n357gat), .I1 (n2726gat), .I2 (n2860gat));
NR3X1 gate2770(.O (n82gat), .I1 (n16gat), .I2 (n295gat), .I3 (n637gat));
NR2X1 gate2771(.O (n12gat), .I1 (n186gat), .I2 (n82gat));
NR2X1 gate2772(.O (n1599gat), .I1 (n1691gat), .I2 (n336gat));
NR2X1 gate2773(.O (n1613gat), .I1 (n1544gat), .I2 (n1698gat));
NR3X1 gate2774(.O (n1756gat), .I1 (n2512gat), .I2 (n1769gat), .I3 (n1773gat));
NR2X1 gate2775(.O (n1586gat), .I1 (n1869gat), .I2 (n1683gat));
NR3X1 gate2776(.O (n1755gat), .I1 (n1769gat), .I2 (n1773gat), .I3 (n2512gat));
NR3X1 gate2777(.O (n2538gat), .I1 (n2620gat), .I2 (n2625gat), .I3 (n2488gat));
NR3X1 gate2778(.O (n2483gat), .I1 (n2537gat), .I2 (n2482gat), .I3 (n2486gat));
NR2X1 gate2779(.O (n1391gat), .I1 (n1513gat), .I2 (n2442gat));
NR3X1 gate2780(.O (n1471gat), .I1 (n1334gat), .I2 (n1858gat), .I3 (n1604gat));
NR2X1 gate2781(.O (n1469gat), .I1 (n1858gat), .I2 (n1608gat));
NR3X1 gate2782(.O (n1472gat), .I1 (n1476gat), .I2 (n1471gat), .I3 (n1469gat));
NR2X1 gate2783(.O (n1927gat), .I1 (n1790gat), .I2 (n1635gat));
NR2X1 gate2784(.O (n1470gat), .I1 (n1472gat), .I2 (n1747gat));
NR3X1 gate2785(.O (n1402gat), .I1 (n1858gat), .I2 (n1393gat), .I3 (n1604gat));
NR2X1 gate2786(.O (n1400gat), .I1 (n1674gat), .I2 (n1403gat));
NR2X1 gate2787(.O (n1567gat), .I1 (n1634gat), .I2 (n1735gat));
NR3X1 gate2788(.O (n1399gat), .I1 (n1806gat), .I2 (n1338gat), .I3 (n1584gat));
NR4X1 gate2789(.O (n1564gat), .I1 (n1584gat), .I2 (n1719gat), .I3 (n1790gat), .I4 (n1576gat));
NR2X1 gate2790(.O (n1600gat), .I1 (n1685gat), .I2 (n1427gat));
NR3X1 gate2791(.O (n1519gat), .I1 (n1584gat), .I2 (n1339gat), .I3 (n1600gat));
NR2X1 gate2792(.O (n1397gat), .I1 (n1519gat), .I2 (n1401gat));
NR2X1 gate2793(.O (n1398gat), .I1 (n1455gat), .I2 (n1397gat));
NR2X1 gate2794(.O (n2008gat), .I1 (n2012gat), .I2 (n1774gat));
NR2X1 gate2795(.O (n2005gat), .I1 (n2002gat), .I2 (n2857gat));
NR2X1 gate2796(.O (n1818gat), .I1 (n1823gat), .I2 (n2005gat));
NR3X1 gate2797(.O (n1759gat), .I1 (n1818gat), .I2 (n1935gat), .I3 (n2765gat));
NR3X1 gate2798(.O (n1686gat), .I1 (n1774gat), .I2 (n1869gat), .I3 (n1684gat));
NR2X1 gate2799(.O (n1533gat), .I1 (n1524gat), .I2 (n1403gat));
NR3X1 gate2800(.O (n1863gat), .I1 (n1991gat), .I2 (n2283gat), .I3 (n1989gat));
NR3X1 gate2801(.O (n1860gat), .I1 (n1988gat), .I2 (n2216gat), .I3 (n1862gat));
NR2X1 gate2802(.O (n1915gat), .I1 (n1859gat), .I2 (n1919gat));
NR2X1 gate2803(.O (n1510gat), .I1 (n1584gat), .I2 (n1460gat));
NR2X1 gate2804(.O (n1800gat), .I1 (n1635gat), .I2 (n1919gat));
NR2X1 gate2805(.O (n1459gat), .I1 (n1595gat), .I2 (n1454gat));
NR2X1 gate2806(.O (n1458gat), .I1 (n1510gat), .I2 (n1459gat));
NR2X1 gate2807(.O (n1532gat), .I1 (n1677gat), .I2 (n1458gat));
NR2X1 gate2808(.O (n1467gat), .I1 (n2289gat), .I2 (n1468gat));
NR3X1 gate2809(.O (n1466gat), .I1 (n1392gat), .I2 (n1461gat), .I3 (n1396gat));
NR2X1 gate2810(.O (n1531gat), .I1 (n1507gat), .I2 (n1477gat));
NR2X1 gate2811(.O (n1593gat), .I1 (n1551gat), .I2 (n1310gat));
NR3X1 gate2812(.O (n1602gat), .I1 (n1594gat), .I2 (n1587gat), .I3 (n2989gat));
NR3X1 gate2813(.O (n1761gat), .I1 (n2985gat), .I2 (n1602gat), .I3 (n1681gat));
NR3X1 gate2814(.O (n1760gat), .I1 (n1681gat), .I2 (n1602gat), .I3 (n2985gat));
NR3X1 gate2815(.O (n1721gat), .I1 (n2442gat), .I2 (n1690gat), .I3 (n1978gat));
NR2X1 gate2816(.O (n520gat), .I1 (n374gat), .I2 (n2862gat));
NR2X1 gate2817(.O (n519gat), .I1 (n2854gat), .I2 (n374gat));
NR2X1 gate2818(.O (n518gat), .I1 (n520gat), .I2 (n519gat));
NR2X1 gate2819(.O (n418gat), .I1 (n374gat), .I2 (n2723gat));
NR2X1 gate2820(.O (n411gat), .I1 (n374gat), .I2 (n2726gat));
NR2X1 gate2821(.O (n522gat), .I1 (n374gat), .I2 (n2859gat));
NR2X1 gate2822(.O (n516gat), .I1 (n374gat), .I2 (n2715gat));
NR4X1 gate2823(.O (n410gat), .I1 (n417gat), .I2 (n413gat), .I3 (n412gat), .I4 (n406gat));
NR2X1 gate2824(.O (n354gat), .I1 (n411gat), .I2 (n522gat));
NR3X1 gate2825(.O (n355gat), .I1 (n517gat), .I2 (n410gat), .I3 (n354gat));
NR2X1 gate2826(.O (n408gat), .I1 (n516gat), .I2 (n407gat));
NR2X1 gate2827(.O (n526gat), .I1 (n2859gat), .I2 (n740gat));
NR2X1 gate2828(.O (n531gat), .I1 (n740gat), .I2 (n2854gat));
NR2X1 gate2829(.O (n530gat), .I1 (n2862gat), .I2 (n740gat));
NR3X1 gate2830(.O (n525gat), .I1 (n526gat), .I2 (n531gat), .I3 (n530gat));
NR2X1 gate2831(.O (n356gat), .I1 (n2726gat), .I2 (n740gat));
NR2X1 gate2832(.O (n415gat), .I1 (n2723gat), .I2 (n740gat));
NR2X1 gate2833(.O (n521gat), .I1 (n740gat), .I2 (n2715gat));
NR3X1 gate2834(.O (n532gat), .I1 (n527gat), .I2 (n416gat), .I3 (n528gat));
NR2X1 gate2835(.O (n359gat), .I1 (n290gat), .I2 (n358gat));
NR2X1 gate2836(.O (n420gat), .I1 (n408gat), .I2 (n359gat));
NR2X1 gate2837(.O (n523gat), .I1 (n522gat), .I2 (n356gat));
NR2X1 gate2838(.O (n634gat), .I1 (n418gat), .I2 (n521gat));
NR2X1 gate2839(.O (n414gat), .I1 (n411gat), .I2 (n415gat));
NR3X1 gate2840(.O (n635gat), .I1 (n639gat), .I2 (n634gat), .I3 (n414gat));
NR2X1 gate2841(.O (n1100gat), .I1 (n1297gat), .I2 (n1111gat));
NR3X1 gate2842(.O (n630gat), .I1 (n634gat), .I2 (n523gat), .I3 (n524gat));
NR2X1 gate2843(.O (n994gat), .I1 (n1112gat), .I2 (n882gat));
NR3X1 gate2844(.O (n629gat), .I1 (n414gat), .I2 (n634gat), .I3 (n523gat));
NR2X1 gate2845(.O (n989gat), .I1 (n721gat), .I2 (n741gat));
NR3X1 gate2846(.O (n632gat), .I1 (n414gat), .I2 (n523gat), .I3 (n633gat));
NR2X1 gate2847(.O (n880gat), .I1 (n926gat), .I2 (n566gat));
NR3X1 gate2848(.O (n636gat), .I1 (n414gat), .I2 (n633gat), .I3 (n639gat));
NR2X1 gate2849(.O (n801gat), .I1 (n672gat), .I2 (n670gat));
NR2X1 gate2850(.O (n879gat), .I1 (n2931gat), .I2 (n801gat));
NR2X1 gate2851(.O (n1003gat), .I1 (n420gat), .I2 (n879gat));
NR2X1 gate2852(.O (n1255gat), .I1 (n1123gat), .I2 (n1225gat));
NR2X1 gate2853(.O (n1012gat), .I1 (n1007gat), .I2 (n918gat));
NR2X1 gate2854(.O (n905gat), .I1 (n625gat), .I2 (n1006gat));
NR2X1 gate2855(.O (n1009gat), .I1 (n1255gat), .I2 (n2943gat));
NR2X1 gate2856(.O (n409gat), .I1 (n406gat), .I2 (n407gat));
NR2X1 gate2857(.O (n292gat), .I1 (n415gat), .I2 (n356gat));
NR2X1 gate2858(.O (n291gat), .I1 (n290gat), .I2 (n292gat));
NR2X1 gate2859(.O (n419gat), .I1 (n409gat), .I2 (n291gat));
NR2X1 gate2860(.O (n902gat), .I1 (n1009gat), .I2 (n419gat));
NR2X1 gate2861(.O (n1099gat), .I1 (n1111gat), .I2 (n1293gat));
NR2X1 gate2862(.O (n998gat), .I1 (n725gat), .I2 (n741gat));
NR2X1 gate2863(.O (n995gat), .I1 (n823gat), .I2 (n1112gat));
NR2X1 gate2864(.O (n980gat), .I1 (n875gat), .I2 (n926gat));
NR2X1 gate2865(.O (n1001gat), .I1 (n420gat), .I2 (n1002gat));
NR2X1 gate2866(.O (n1175gat), .I1 (n621gat), .I2 (n1006gat));
NR2X1 gate2867(.O (n1174gat), .I1 (n845gat), .I2 (n1007gat));
NR2X1 gate2868(.O (n1243gat), .I1 (n1281gat), .I2 (n1123gat));
NR2X1 gate2869(.O (n1171gat), .I1 (n2960gat), .I2 (n1243gat));
NR2X1 gate2870(.O (n999gat), .I1 (n419gat), .I2 (n1171gat));
NR2X1 gate2871(.O (n1244gat), .I1 (n1123gat), .I2 (n1134gat));
NR2X1 gate2872(.O (n1323gat), .I1 (n1007gat), .I2 (n401gat));
NR2X1 gate2873(.O (n1264gat), .I1 (n1006gat), .I2 (n617gat));
NR2X1 gate2874(.O (n1265gat), .I1 (n1244gat), .I2 (n2969gat));
NR2X1 gate2875(.O (n892gat), .I1 (n419gat), .I2 (n1265gat));
NR2X1 gate2876(.O (n981gat), .I1 (n926gat), .I2 (n873gat));
NR2X1 gate2877(.O (n890gat), .I1 (n741gat), .I2 (n702gat));
NR2X1 gate2878(.O (n889gat), .I1 (n1111gat), .I2 (n1079gat));
NR2X1 gate2879(.O (n886gat), .I1 (n683gat), .I2 (n1112gat));
NR2X1 gate2880(.O (n891gat), .I1 (n420gat), .I2 (n888gat));
NR2X1 gate2881(.O (n904gat), .I1 (n1006gat), .I2 (n490gat));
NR2X1 gate2882(.O (n903gat), .I1 (n1007gat), .I2 (n397gat));
NR2X1 gate2883(.O (n1254gat), .I1 (n1123gat), .I2 (n1044gat));
NR2X1 gate2884(.O (n1008gat), .I1 (n2942gat), .I2 (n1254gat));
NR2X1 gate2885(.O (n900gat), .I1 (n419gat), .I2 (n1008gat));
NR2X1 gate2886(.O (n1152gat), .I1 (n926gat), .I2 (n1150gat));
NR2X1 gate2887(.O (n1092gat), .I1 (n1147gat), .I2 (n1111gat));
NR2X1 gate2888(.O (n997gat), .I1 (n741gat), .I2 (n393gat));
NR2X1 gate2889(.O (n993gat), .I1 (n1112gat), .I2 (n698gat));
NR2X1 gate2890(.O (n895gat), .I1 (n420gat), .I2 (n898gat));
NR2X1 gate2891(.O (n1094gat), .I1 (n1112gat), .I2 (n583gat));
NR2X1 gate2892(.O (n1093gat), .I1 (n1111gat), .I2 (n864gat));
NR2X1 gate2893(.O (n988gat), .I1 (n340gat), .I2 (n741gat));
NR2X1 gate2894(.O (n984gat), .I1 (n926gat), .I2 (n983gat));
NR2X1 gate2895(.O (n1178gat), .I1 (n420gat), .I2 (n1179gat));
NR2X1 gate2896(.O (n1267gat), .I1 (n613gat), .I2 (n1006gat));
NR2X1 gate2897(.O (n1257gat), .I1 (n1007gat), .I2 (n274gat));
NR2X1 gate2898(.O (n1253gat), .I1 (n930gat), .I2 (n1123gat));
NR2X1 gate2899(.O (n1266gat), .I1 (n2965gat), .I2 (n1253gat));
NR2X1 gate2900(.O (n1116gat), .I1 (n419gat), .I2 (n1266gat));
NR2X1 gate2901(.O (n1375gat), .I1 (n1006gat), .I2 (n706gat));
NR2X1 gate2902(.O (n1324gat), .I1 (n164gat), .I2 (n1007gat));
NR2X1 gate2903(.O (n1200gat), .I1 (n1120gat), .I2 (n1123gat));
NR2X1 gate2904(.O (n1172gat), .I1 (n2961gat), .I2 (n1200gat));
NR2X1 gate2905(.O (n899gat), .I1 (n419gat), .I2 (n1172gat));
NR2X1 gate2906(.O (n1091gat), .I1 (n1111gat), .I2 (n956gat));
NR2X1 gate2907(.O (n1088gat), .I1 (n1085gat), .I2 (n926gat));
NR2X1 gate2908(.O (n992gat), .I1 (n815gat), .I2 (n1112gat));
NR2X1 gate2909(.O (n987gat), .I1 (n741gat), .I2 (n159gat));
NR2X1 gate2910(.O (n896gat), .I1 (n897gat), .I2 (n420gat));
NR2X1 gate2911(.O (n1262gat), .I1 (n837gat), .I2 (n1006gat));
NR2X1 gate2912(.O (n1260gat), .I1 (n1007gat), .I2 (n278gat));
NR2X1 gate2913(.O (n1251gat), .I1 (n1123gat), .I2 (n1071gat));
NR2X1 gate2914(.O (n1259gat), .I1 (n2967gat), .I2 (n1251gat));
NR2X1 gate2915(.O (n901gat), .I1 (n419gat), .I2 (n1259gat));
NR2X1 gate2916(.O (n1098gat), .I1 (n336gat), .I2 (n741gat));
NR2X1 gate2917(.O (n1090gat), .I1 (n1111gat), .I2 (n860gat));
NR2X1 gate2918(.O (n986gat), .I1 (n985gat), .I2 (n926gat));
NR2X1 gate2919(.O (n885gat), .I1 (n579gat), .I2 (n1112gat));
NR2X1 gate2920(.O (n893gat), .I1 (n894gat), .I2 (n420gat));
NR2X1 gate2921(.O (n1097gat), .I1 (n270gat), .I2 (n741gat));
NR2X1 gate2922(.O (n1089gat), .I1 (n1067gat), .I2 (n1111gat));
NR2X1 gate2923(.O (n1087gat), .I1 (n926gat), .I2 (n1084gat));
NR2X1 gate2924(.O (n991gat), .I1 (n1112gat), .I2 (n679gat));
NR2X1 gate2925(.O (n1177gat), .I1 (n1180gat), .I2 (n420gat));
NR2X1 gate2926(.O (n1212gat), .I1 (n1123gat), .I2 (n1034gat));
NR2X1 gate2927(.O (n1326gat), .I1 (n1007gat), .I2 (n282gat));
NR2X1 gate2928(.O (n1261gat), .I1 (n833gat), .I2 (n1006gat));
NR2X1 gate2929(.O (n1263gat), .I1 (n1212gat), .I2 (n2968gat));
NR2X1 gate2930(.O (n1115gat), .I1 (n1263gat), .I2 (n419gat));
NR2X1 gate2931(.O (n977gat), .I1 (n670gat), .I2 (n671gat));
NR3X1 gate2932(.O (n631gat), .I1 (n523gat), .I2 (n633gat), .I3 (n524gat));
NR2X1 gate2933(.O (n1096gat), .I1 (n819gat), .I2 (n1112gat));
NR2X1 gate2934(.O (n1095gat), .I1 (n1240gat), .I2 (n1111gat));
NR2X1 gate2935(.O (n990gat), .I1 (n841gat), .I2 (n741gat));
NR2X1 gate2936(.O (n979gat), .I1 (n1601gat), .I2 (n926gat));
NR2X1 gate2937(.O (n978gat), .I1 (n2944gat), .I2 (n2945gat));
NR2X1 gate2938(.O (n1004gat), .I1 (n978gat), .I2 (n420gat));
NR2X1 gate2939(.O (n1199gat), .I1 (n1123gat), .I2 (n1284gat));
NR2X1 gate2940(.O (n1176gat), .I1 (n829gat), .I2 (n1006gat));
NR2X1 gate2941(.O (n1173gat), .I1 (n1007gat), .I2 (n1025gat));
NR2X1 gate2942(.O (n1252gat), .I1 (n1199gat), .I2 (n2962gat));
NR2X1 gate2943(.O (n1000gat), .I1 (n419gat), .I2 (n1252gat));
NR2X1 gate2944(.O (n1029gat), .I1 (n978gat), .I2 (n455gat));
NR2X1 gate2945(.O (n1028gat), .I1 (n455gat), .I2 (n879gat));
NR2X1 gate2946(.O (n1031gat), .I1 (n1002gat), .I2 (n455gat));
NR2X1 gate2947(.O (n1030gat), .I1 (n455gat), .I2 (n888gat));
NR2X1 gate2948(.O (n1011gat), .I1 (n455gat), .I2 (n898gat));
NR2X1 gate2949(.O (n1181gat), .I1 (n455gat), .I2 (n1179gat));
NR2X1 gate2950(.O (n1010gat), .I1 (n897gat), .I2 (n455gat));
NR2X1 gate2951(.O (n1005gat), .I1 (n894gat), .I2 (n455gat));
NR2X1 gate2952(.O (n1182gat), .I1 (n1180gat), .I2 (n455gat));
NR2X1 gate2953(.O (n1757gat), .I1 (n1773gat), .I2 (n1769gat));
NR2X1 gate2954(.O (n1745gat), .I1 (n1869gat), .I2 (n1757gat));
NR2X1 gate2955(.O (n73gat), .I1 (n67gat), .I2 (n2784gat));
NR2X1 gate2956(.O (n70gat), .I1 (n71gat), .I2 (n2720gat));
NR2X1 gate2957(.O (n77gat), .I1 (n76gat), .I2 (n2784gat));
NR2X1 gate2958(.O (n13gat), .I1 (n2720gat), .I2 (n14gat));
endmodule