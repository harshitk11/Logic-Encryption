
module s5378_0 ( clk, n3065gat, n3066gat, n3067gat, n3068gat, n3069gat, 
        n3070gat, n3071gat, n3072gat, n3073gat, n3074gat, n3075gat, n3076gat, 
        n3077gat, n3078gat, n3079gat, n3080gat, n3081gat, n3082gat, n3083gat, 
        n3084gat, n3085gat, n3086gat, n3087gat, n3088gat, n3089gat, n3090gat, 
        n3091gat, n3092gat, n3093gat, n3094gat, n3095gat, n3097gat, n3098gat, 
        n3099gat, n3100gat, key_1, key_2, key_3, key_4, key_5, key_6, key_7, 
        key_8, key_9, key_10, key_11, key_12, key_13, key_14, key_15, key_16, 
        key_17, key_18, key_19, key_20, key_21, key_22, key_23, key_24, key_25, 
        key_26, key_27, key_28, key_29, key_30, key_31, key_32, key_33, key_34, 
        key_35, key_36, key_37, key_38, key_39, key_40, key_41, key_42, key_43, 
        key_44, key_45, key_46, key_47, key_48, key_49, key_50, key_51, key_52, 
        key_53, key_54, key_55, key_56, key_57, key_58, key_59, key_60, key_61, 
        key_62, key_63, key_64, key_65, key_66, key_67, key_68, key_69, key_70, 
        key_71, key_72, key_73, key_74, key_75, key_76, key_77, key_78, key_79, 
        key_80, key_81, key_82, key_83, key_84, key_85, key_86, key_87, key_88, 
        key_89, key_90, key_91, key_92, key_93, key_94, key_95, key_96, key_97, 
        key_98, key_99, key_100, key_101, key_102, key_103, key_104, key_105, 
        key_106, key_107, key_108, key_109, key_110, key_111, key_112, key_113, 
        key_114, key_115, key_116, key_117, key_118, key_119, key_120, key_121, 
        key_122, key_123, key_124, key_125, key_126, key_127, key_128, 
        n3104gat, n3105gat, n3106gat, n3107gat, n3108gat, n3109gat, n3110gat, 
        n3111gat, n3112gat, n3113gat, n3114gat, n3115gat, n3116gat, n3117gat, 
        n3118gat, n3119gat, n3120gat, n3121gat, n3122gat, n3123gat, n3124gat, 
        n3125gat, n3126gat, n3127gat, n3128gat, n3129gat, n3130gat, n3131gat, 
        n3132gat, n3133gat, n3134gat, n3135gat, n3136gat, n3137gat, n3138gat, 
        n3139gat, n3140gat, n3141gat, n3142gat, n3143gat, n3144gat, n3145gat, 
        n3146gat, n3147gat, n3148gat, n3149gat, n3150gat, n3151gat, n3152gat, 
        test_si, test_so, test_se );
  input clk, n3065gat, n3066gat, n3067gat, n3068gat, n3069gat, n3070gat,
         n3071gat, n3072gat, n3073gat, n3074gat, n3075gat, n3076gat, n3077gat,
         n3078gat, n3079gat, n3080gat, n3081gat, n3082gat, n3083gat, n3084gat,
         n3085gat, n3086gat, n3087gat, n3088gat, n3089gat, n3090gat, n3091gat,
         n3092gat, n3093gat, n3094gat, n3095gat, n3097gat, n3098gat, n3099gat,
         n3100gat, key_1, key_2, key_3, key_4, key_5, key_6, key_7, key_8,
         key_9, key_10, key_11, key_12, key_13, key_14, key_15, key_16, key_17,
         key_18, key_19, key_20, key_21, key_22, key_23, key_24, key_25,
         key_26, key_27, key_28, key_29, key_30, key_31, key_32, key_33,
         key_34, key_35, key_36, key_37, key_38, key_39, key_40, key_41,
         key_42, key_43, key_44, key_45, key_46, key_47, key_48, key_49,
         key_50, key_51, key_52, key_53, key_54, key_55, key_56, key_57,
         key_58, key_59, key_60, key_61, key_62, key_63, key_64, key_65,
         key_66, key_67, key_68, key_69, key_70, key_71, key_72, key_73,
         key_74, key_75, key_76, key_77, key_78, key_79, key_80, key_81,
         key_82, key_83, key_84, key_85, key_86, key_87, key_88, key_89,
         key_90, key_91, key_92, key_93, key_94, key_95, key_96, key_97,
         key_98, key_99, key_100, key_101, key_102, key_103, key_104, key_105,
         key_106, key_107, key_108, key_109, key_110, key_111, key_112,
         key_113, key_114, key_115, key_116, key_117, key_118, key_119,
         key_120, key_121, key_122, key_123, key_124, key_125, key_126,
         key_127, key_128, test_si, test_se;
  output n3104gat, n3105gat, n3106gat, n3107gat, n3108gat, n3109gat, n3110gat,
         n3111gat, n3112gat, n3113gat, n3114gat, n3115gat, n3116gat, n3117gat,
         n3118gat, n3119gat, n3120gat, n3121gat, n3122gat, n3123gat, n3124gat,
         n3125gat, n3126gat, n3127gat, n3128gat, n3129gat, n3130gat, n3131gat,
         n3132gat, n3133gat, n3134gat, n3135gat, n3136gat, n3137gat, n3138gat,
         n3139gat, n3140gat, n3141gat, n3142gat, n3143gat, n3144gat, n3145gat,
         n3146gat, n3147gat, n3148gat, n3149gat, n3150gat, n3151gat, n3152gat,
         test_so;
  wire   n1821gat, n3146gat, n2579gat, n2874gat, n2885gat, n2875gat, n2881gat,
         n3108gat, n3094gat, n1827gat, n1793gat, n2009gat, n2015gat, n2017gat,
         n2194gat, n2396gat, n2198gat, n2197gat, n2196gat, n153, n157, n256,
         n268, n273, n3139gat, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n329, n333,
         n339, n352, n354, n359, n360, n361, n362, n363, n364, n368, n369,
         n370, n371, n373, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461;
  assign n3105gat = n3146gat;
  assign n3124gat = n3146gat;
  assign n3141gat = n3146gat;
  assign n3142gat = n3146gat;
  assign n3129gat = n3146gat;
  assign n3137gat = n3146gat;
  assign n3117gat = n3146gat;
  assign n3130gat = n3146gat;
  assign n3119gat = n3146gat;
  assign n3132gat = n3146gat;
  assign n3131gat = n3146gat;
  assign n3136gat = n3146gat;
  assign n3133gat = n3146gat;
  assign n3135gat = n3146gat;
  assign n3134gat = n3146gat;
  assign n3138gat = n3146gat;
  assign n3150gat = n3108gat;
  assign n3147gat = n3108gat;
  assign n3143gat = n3108gat;
  assign n3113gat = n3108gat;
  assign n3111gat = n3108gat;
  assign n3110gat = n3108gat;
  assign n3109gat = n3108gat;
  assign n3115gat = n3108gat;
  assign n3152gat = n3108gat;
  assign n3151gat = n3108gat;
  assign n3112gat = n3108gat;
  assign n3120gat = n3108gat;
  assign n3118gat = n3108gat;
  assign n3116gat = n3108gat;
  assign n3148gat = n3108gat;
  assign n3145gat = n3108gat;
  assign n3107gat = n3108gat;
  assign n3123gat = n3108gat;
  assign n3149gat = n3108gat;
  assign n3114gat = n3108gat;
  assign n3104gat = n3094gat;
  assign n3140gat = n3139gat;

  DFZX1 gate19 ( .D(n1827gat), .TD(test_si), .SEL(test_se), .CK(clk), .Q(
        n1821gat) );
  DFZX1 gate20 ( .D(n1827gat), .TD(n1821gat), .SEL(test_se), .CK(clk), .Q(n425), .QB(n373) );
  DFZX1 gate21 ( .D(n311), .TD(n425), .SEL(test_se), .CK(clk), .Q(n461), .QB(
        n312) );
  DFZX1 gate22 ( .D(n312), .TD(n461), .SEL(test_se), .CK(clk), .Q(n460), .QB(
        n256) );
  DFZX1 gate43 ( .D(n2881gat), .TD(n460), .SEL(test_se), .CK(clk), .Q(n421), 
        .QB(n313) );
  DFZX1 gate44 ( .D(n2874gat), .TD(n421), .SEL(test_se), .CK(clk), .Q(n419), 
        .QB(n314) );
  DFZX1 gate45 ( .D(n363), .TD(n419), .SEL(test_se), .CK(clk), .Q(n422), .QB(
        n315) );
  DFZX1 gate46 ( .D(n364), .TD(n422), .SEL(test_se), .CK(clk), .Q(n416), .QB(
        n316) );
  DFZX1 gate47 ( .D(n359), .TD(n416), .SEL(test_se), .CK(clk), .Q(n420), .QB(
        n317) );
  DFZX1 gate52 ( .D(n2885gat), .TD(n420), .SEL(test_se), .CK(clk), .Q(n435), 
        .QB(n318) );
  DFZX1 gate53 ( .D(n361), .TD(n435), .SEL(test_se), .CK(clk), .Q(n436), .QB(
        n319) );
  DFZX1 gate54 ( .D(n360), .TD(n436), .SEL(test_se), .CK(clk), .Q(n417), .QB(
        n320) );
  DFZX1 gate56 ( .D(n362), .TD(n417), .SEL(test_se), .CK(clk), .Q(n459), .QB(
        n321) );
  DFZX1 gate57 ( .D(n2875gat), .TD(n459), .SEL(test_se), .CK(clk), .Q(n418), 
        .QB(n322) );
  DFZX1 gate59 ( .D(n2396gat), .TD(n418), .SEL(test_se), .CK(clk), .Q(n426), 
        .QB(n323) );
  DFZX1 gate60 ( .D(n2198gat), .TD(n426), .SEL(test_se), .CK(clk), .Q(n427), 
        .QB(n324) );
  DFZX1 gate61 ( .D(n2196gat), .TD(n427), .SEL(test_se), .CK(clk), .Q(n428), 
        .QB(n325) );
  DFZX1 gate62 ( .D(n153), .TD(n428), .SEL(test_se), .CK(clk), .Q(n458), .QB(
        n326) );
  DFZX1 gate63 ( .D(n2197gat), .TD(n458), .SEL(test_se), .CK(clk), .Q(n429), 
        .QB(n327) );
  DFZX1 gate94 ( .D(n329), .TD(n429), .SEL(test_se), .CK(clk), .Q(n423), .QB(
        n333) );
  DFZX1 gate97 ( .D(n157), .TD(n423), .SEL(test_se), .CK(clk), .Q(n457), .QB(
        n3128gat) );
  DFZX1 gate98 ( .D(n2194gat), .TD(n457), .SEL(test_se), .CK(clk), .Q(n456), 
        .QB(n3127gat) );
  DFZX1 gate99 ( .D(n3146gat), .TD(n456), .SEL(test_se), .CK(clk), .Q(n455), 
        .QB(n3126gat) );
  DFZX1 gate111 ( .D(n323), .TD(n455), .SEL(test_se), .CK(clk), .Q(n454), .QB(
        n368) );
  DFZX1 gate112 ( .D(n324), .TD(n454), .SEL(test_se), .CK(clk), .Q(n430), .QB(
        n369) );
  DFZX1 gate113 ( .D(n326), .TD(n430), .SEL(test_se), .CK(clk), .Q(n431), .QB(
        n371) );
  DFZX1 gate114 ( .D(n327), .TD(n431), .SEL(test_se), .CK(clk), .Q(n432) );
  DFZX1 gate115 ( .D(n325), .TD(n432), .SEL(test_se), .CK(clk), .Q(n433), .QB(
        n370) );
  DFZX1 gate116 ( .D(n1793gat), .TD(n433), .SEL(test_se), .CK(clk), .Q(n453), 
        .QB(n273) );
  DFZX1 gate128 ( .D(n3146gat), .TD(n453), .SEL(test_se), .CK(clk), .Q(n452), 
        .QB(n339) );
  DFZX1 gate129 ( .D(n339), .TD(n452), .SEL(test_se), .CK(clk), .Q(n424) );
  DFZX1 gate133 ( .D(n2009gat), .TD(n424), .SEL(test_se), .CK(clk), .Q(n451), 
        .QB(n3106gat) );
  DFZX1 gate145 ( .D(n2015gat), .TD(n451), .SEL(test_se), .CK(clk), .Q(n450), 
        .QB(n352) );
  DFZX1 gate146 ( .D(n352), .TD(n450), .SEL(test_se), .CK(clk), .Q(n434) );
  DFZX1 gate147 ( .D(n2017gat), .TD(n434), .SEL(test_se), .CK(clk), .Q(n449), 
        .QB(n354) );
  DFZX1 gate148 ( .D(n354), .TD(n449), .SEL(test_se), .CK(clk), .Q(n448), .QB(
        n268) );
  DFZX1 gate156 ( .D(n333), .TD(n448), .SEL(test_se), .CK(clk), .Q(n415) );
  DFZX1 gate157 ( .D(n317), .TD(n415), .SEL(test_se), .CK(clk), .Q(n447), .QB(
        n359) );
  DFZX1 gate158 ( .D(n314), .TD(n447), .SEL(test_se), .CK(clk), .Q(n446), .QB(
        n2874gat) );
  DFZX1 gate159 ( .D(n318), .TD(n446), .SEL(test_se), .CK(clk), .Q(n445), .QB(
        n2885gat) );
  DFZX1 gate160 ( .D(n320), .TD(n445), .SEL(test_se), .CK(clk), .Q(n444), .QB(
        n360) );
  DFZX1 gate161 ( .D(n319), .TD(n444), .SEL(test_se), .CK(clk), .Q(n443), .QB(
        n361) );
  DFZX1 gate162 ( .D(n321), .TD(n443), .SEL(test_se), .CK(clk), .Q(n442), .QB(
        n362) );
  DFZX1 gate163 ( .D(n322), .TD(n442), .SEL(test_se), .CK(clk), .Q(n441), .QB(
        n2875gat) );
  DFZX1 gate164 ( .D(n315), .TD(n441), .SEL(test_se), .CK(clk), .Q(n440), .QB(
        n363) );
  DFZX1 gate165 ( .D(n316), .TD(n440), .SEL(test_se), .CK(clk), .Q(n439), .QB(
        n364) );
  DFZX1 gate166 ( .D(n313), .TD(n439), .SEL(test_se), .CK(clk), .Q(test_so), 
        .QB(n2881gat) );
  TIE1X1 U171 ( .O(n3108gat) );
  TIE0X1 U172 ( .O(n3146gat) );
  MOAI1X1 U173 ( .A1(n395), .A2(n396), .B1(n3108gat), .B2(n397), .O(n394) );
  INVCKX2 U174 ( .I(n395), .O(n393) );
  INVCKX2 U175 ( .I(n405), .O(n2194gat) );
  XOR4XLP U176 ( .I1(n418), .I2(n321), .I3(n417), .I4(n3108gat), .O(n383) );
  AN2B1X2 U177 ( .I1(n431), .B1(n368), .O(n414) );
  AN4B2X1 U178 ( .I1(n411), .I2(n3108gat), .B1(n433), .B2(n3146gat), .O(n409)
         );
  INVCKX2 U179 ( .I(n413), .O(n1793gat) );
  NR2X2 U180 ( .I1(n390), .I2(n273), .O(n389) );
  OA22X1 U181 ( .A1(n3128gat), .A2(n3146gat), .B1(n3126gat), .B2(n3127gat), 
        .O(n3125gat) );
  INVCKX2 U182 ( .I(n3099gat), .O(n1827gat) );
  INVCKX2 U183 ( .I(n422), .O(n382) );
  INVCKX2 U184 ( .I(n378), .O(n3139gat) );
  INVCKX2 U185 ( .I(n410), .O(n2009gat) );
  INVCKX2 U186 ( .I(n424), .O(n2015gat) );
  OR4X1 U187 ( .I1(n379), .I2(n3098gat), .I3(n380), .I4(n3146gat), .O(n378) );
  XOR2X2 U188 ( .I1(n436), .I2(n435), .O(n384) );
  XNR2X2 U189 ( .I1(n384), .I2(n383), .O(n3121gat) );
  XOR4XLP U190 ( .I1(n420), .I2(n421), .I3(n416), .I4(n3146gat), .O(n381) );
  INVCKX2 U191 ( .I(n323), .O(n396) );
  INVCKX2 U192 ( .I(n426), .O(n399) );
  INVCKX2 U193 ( .I(n323), .O(n398) );
  INVCKX2 U194 ( .I(n373), .O(n379) );
  INVCKX2 U195 ( .I(n409), .O(n2017gat) );
  OAI12X1 U196 ( .B1(n3146gat), .B2(n268), .A1(n434), .O(n405) );
  ND2X1 U197 ( .I1(n375), .I2(n153), .O(n329) );
  XOR2X1 U198 ( .I1(n376), .I2(n415), .O(n375) );
  OAI112X1 U199 ( .C1(n430), .C2(n368), .A1(n377), .B1(n371), .O(n376) );
  XOR3X1 U200 ( .I1(n381), .I2(n382), .I3(n419), .O(n3122gat) );
  ND2X1 U201 ( .I1(n2579gat), .I2(n386), .O(n3144gat) );
  INVCKX1 U202 ( .I(n389), .O(n386) );
  OA13X1 U203 ( .B1(n428), .B2(n327), .B3(n391), .A1(n392), .O(n390) );
  MXL2XLP U204 ( .A(n393), .B(n394), .S(n427), .OB(n392) );
  MXL2XLP U205 ( .A(n398), .B(n399), .S(n427), .OB(n391) );
  XOR4XLP U206 ( .I1(n423), .I2(n427), .I3(n326), .I4(n402), .O(n2579gat) );
  MUXB2X1 U207 ( .EB(n397), .A(n403), .B(n404), .S(n426), .O(n402) );
  ND2X1 U208 ( .I1(n428), .I2(n327), .O(n404) );
  OA12X1 U209 ( .B1(n429), .B2(n428), .A1(n395), .O(n403) );
  ND2X1 U210 ( .I1(n428), .I2(n429), .O(n395) );
  NR3X1 U211 ( .I1(n323), .I2(n428), .I3(n327), .O(n397) );
  NR2X1 U212 ( .I1(n406), .I2(n401), .O(n2396gat) );
  XNR2X1 U213 ( .I1(n368), .I2(n407), .O(n401) );
  NR2X1 U214 ( .I1(n400), .I2(n406), .O(n2198gat) );
  NR2X1 U215 ( .I1(n406), .I2(n388), .O(n2197gat) );
  XNR2X1 U216 ( .I1(n377), .I2(n432), .O(n388) );
  NR2X1 U217 ( .I1(n406), .I2(n387), .O(n2196gat) );
  ND2X1 U218 ( .I1(n377), .I2(n408), .O(n387) );
  AO12X1 U219 ( .B1(n368), .B2(n407), .A1(n370), .O(n408) );
  ND3X1 U220 ( .I1(n370), .I2(n368), .I3(n407), .O(n377) );
  NR2X1 U221 ( .I1(n430), .I2(n431), .O(n407) );
  INVCKX1 U222 ( .I(n2017gat), .O(n410) );
  AN2B1XLP U223 ( .I1(n256), .B1(n311), .O(n380) );
  ND2X1 U224 ( .I1(n425), .I2(n1821gat), .O(n311) );
  ND3X1 U225 ( .I1(n431), .I2(n369), .I3(n412), .O(n413) );
  AN3X1 U226 ( .I1(n432), .I2(n370), .I3(n368), .O(n412) );
  INVCKX1 U227 ( .I(n406), .O(n153) );
  ND2X1 U228 ( .I1(n157), .I2(n385), .O(n406) );
  OR4B2XLP U229 ( .I1(n432), .I2(n400), .B1(n370), .B2(n414), .O(n385) );
  INVCKX1 U230 ( .I(n405), .O(n157) );
  AN3B2X1 U231 ( .I1(n400), .B1(n368), .B2(n432), .O(n411) );
  NR2X1 U232 ( .I1(n369), .I2(n371), .O(n400) );
endmodule

