module s9234(clk, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23, key_1, key_2, key_3, key_4, key_5, key_6, key_7, key_8, key_9, key_10, key_11, key_12, key_13, key_14, key_15, key_16, key_17, key_18, key_19, key_20, key_21, key_22, key_23, key_24, key_25, key_26, key_27, key_28, key_29, key_30, key_31, key_32, key_33, key_34, key_35, key_36, key_37, key_38, key_39, key_40, key_41, key_42, key_43, key_44, key_45, key_46, key_47, key_48, key_49, key_50, key_51, key_52, key_53, key_54, key_55, key_56, key_57, key_58, key_59, key_60, key_61, key_62, key_63, key_64, key_65, key_66, key_67, key_68, key_69, key_70, key_71, key_72, key_73, key_74, key_75, key_76, key_77, key_78, key_79, key_80, key_81, key_82, key_83, key_84, key_85, key_86, key_87, key_88, key_89, key_90, key_91, key_92, key_93, key_94, key_95, key_96, key_97, key_98, key_99, key_100, key_101, key_102, key_103, key_104, key_105, key_106, key_107, key_108, key_109, key_110, key_111, key_112, key_113, key_114, key_115, key_116, key_117, key_118, key_119, key_120, key_121, key_122, key_123, key_124, key_125, key_126, key_127, key_128, g2584, g3222, g3600, g4307, g4321, g4422, g4809, g5137, g5468, g5469, g5692, g6282, g6284, g6360, g6362, g6364, g6366, g6368, g6370, g6372, g6374, g6728, g1290, g4121, g4108, g4106, g4103, g1293, g4099, g4102, g4109, g4100, g4112, g4105, g4101, g4110, g4104, g4107, g4098);
input clk, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23, key_1, key_2, key_3, key_4, key_5, key_6, key_7, key_8, key_9, key_10, key_11, key_12, key_13, key_14, key_15, key_16, key_17, key_18, key_19, key_20, key_21, key_22, key_23, key_24, key_25, key_26, key_27, key_28, key_29, key_30, key_31, key_32, key_33, key_34, key_35, key_36, key_37, key_38, key_39, key_40, key_41, key_42, key_43, key_44, key_45, key_46, key_47, key_48, key_49, key_50, key_51, key_52, key_53, key_54, key_55, key_56, key_57, key_58, key_59, key_60, key_61, key_62, key_63, key_64, key_65, key_66, key_67, key_68, key_69, key_70, key_71, key_72, key_73, key_74, key_75, key_76, key_77, key_78, key_79, key_80, key_81, key_82, key_83, key_84, key_85, key_86, key_87, key_88, key_89, key_90, key_91, key_92, key_93, key_94, key_95, key_96, key_97, key_98, key_99, key_100, key_101, key_102, key_103, key_104, key_105, key_106, key_107, key_108, key_109, key_110, key_111, key_112, key_113, key_114, key_115, key_116, key_117, key_118, key_119, key_120, key_121, key_122, key_123, key_124, key_125, key_126, key_127, key_128;
output g2584, g3222, g3600, g4307, g4321, g4422, g4809, g5137, g5468, g5469, g5692, g6282, g6284, g6360, g6362, g6364, g6366, g6368, g6370, g6372, g6374, g6728, g1290, g4121, g4108, g4106, g4103, g1293, g4099, g4102, g4109, g4100, g4112, g4105, g4101, g4110, g4104, g4107, g4098;
wire clk, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23, key_1, key_2, key_3, key_4, key_5, key_6, key_7, key_8, key_9, key_10, key_11, key_12, key_13, key_14, key_15, key_16, key_17, key_18, key_19, key_20, key_21, key_22, key_23, key_24, key_25, key_26, key_27, key_28, key_29, key_30, key_31, key_32, key_33, key_34, key_35, key_36, key_37, key_38, key_39, key_40, key_41, key_42, key_43, key_44, key_45, key_46, key_47, key_48, key_49, key_50, key_51, key_52, key_53, key_54, key_55, key_56, key_57, key_58, key_59, key_60, key_61, key_62, key_63, key_64, key_65, key_66, key_67, key_68, key_69, key_70, key_71, key_72, key_73, key_74, key_75, key_76, key_77, key_78, key_79, key_80, key_81, key_82, key_83, key_84, key_85, key_86, key_87, key_88, key_89, key_90, key_91, key_92, key_93, key_94, key_95, key_96, key_97, key_98, key_99, key_100, key_101, key_102, key_103, key_104, key_105, key_106, key_107, key_108, key_109, key_110, key_111, key_112, key_113, key_114, key_115, key_116, key_117, key_118, key_119, key_120, key_121, key_122, key_123, key_124, key_125, key_126, key_127, key_128;
wire g678, g332, g123, g207, g695, g461, g18, g292, g331, g689, g24;
wire g465, g84, g291, g676, key_out_112, g622, g117, g278, g128, g598, g554;
wire g496, g179, g48, g590, g551, g682, g11, g606, g188, g646, g327;
wire g361, g289, g398, g684, g619, g208, g248, g390, g625, g681, g437;
wire g276, g3, g323, g224, g685, g43, g157, g282, g697, g206, g449;
wire g118, g528, g284, g426, g634, g669, g520, g281, g175, g15, g631;
wire g69, g693, g337, g457, g486, g471, g328, g285, g418, g402, g297;
wire g212, g410, g430, g33, g662, g453, g269, g574, g441, g664, g349;
wire g211, g586, g571, g29, g326, g698, g654, g293, g690, g445, g374;
wire g6, g687, g357, g386, g504, g665, g166, g541, g74, g338, g696;
wire g516, g536, g683, g353, g545, g254, g341, g290, g2, g287, g336;
wire g345, g628, g679, g28, g688, g283, g613, g10, g14, g680, g143;
wire g672, g667, g366, g279, g492, g170, g686, g288, g638, g602, g642;
wire g280, g663, g610, g148, g209, g675, g478, g122, g54, g594, g286;
wire g489, g616, g79, g218, g242, g578, g184, g119, g668, g139, g422;
wire g210, g394, g230, g25, g204, g658, g650, g378, g508, g548, g370;
wire g406, g236, g500, g205, g197, g666, g114, g524, g260, g111, g131;
wire g7, g19, g677, g582, g485, g699, g193, g135, g382, g414, g434;
wire g266, g49, g152, g692, g277, g127, g161, g512, g532, g64, g694;
wire g691, g1, g59, I8854, g1289, key_out_103, I9125, I6783, I4424, g6895, g1835;
wire I3040, g6837, I7466, I4809, g3537, g5457, g6062, g4040, I6001, g5549, I4477;
wire g3612, I7055, g2892, I5264, I2225, g4123, g4323, g908, I5933, I8252, I2473;
wire I7333, I8812, g1674, I3528, I8958, I5050, g3234, I2324, g2945, g5121, g1997;
wire g3128, I8005, g1541, g5670, g2738, g6842, g4528, g2244, g6192, g2709, g1332;
wire g4530, g1680, g2078, g1209, key_out_128, I3010, g5813, I7509, I5379, g3800, g2907;
wire g6854, g2035, g2959, g6941, g4010, I2287, I4273, I8270, g5740, I5777, g2876;
wire g873, g4839, I5882, g2656, I8473, I2199, g900, g6708, I2399, I3278, g6520;
wire g940, I6677, g3902, g5687, g2915, g847, I3235, I3343, g6431, g709, g6812;
wire I6576, g749, g3090, I9107, g2214, g4618, g6376, g4143, key_out_95, I6349, g4343;
wire I5674, I8177, g2110, I3134, g6405, I3334, I7197, g4566, I7397, I4534, g1714;
wire I4961, g2663, g3456, g5141, g922, g4693, g4134, g5570, g5860, g4334, I3804;
wire I2207, I5153, g3355, g5645, g6733, g5691, g4804, I9047, I4414, g6610, g2877;
wire I4903, g6796, g3063, I3313, g5879, g3463, I4513, g1623, g5358, I3202, I2215;
wire g4113, g1076, g6069, I7817, g6540, I6352, I1865, g4202, I6867, I5511, g5587;
wire I8144, g1175, g1375, g3118, g3318, g2464, g3872, g4494, I2870, g4518, I4288;
wire g5615, g4567, I4382, I3776, g3057, I5600, I3593, I2825, g1285, g3457, g5174;
wire I6386, I3965, I8488, g6849, I6599, I2408, g3834, g2295, g1384, g1339, g5545;
wire I6170, I9128, g6898, g1838, g6900, g2194, g6797, g2394, I3050, I3641, I2943;
wire I5736, g6510, I6280, g4933, g5420, g4521, g1672, I7058, I2887, I2122, g1477;
wire g3232, I2228, g5794, g1643, I4495, I4437, g2705, g3813, I8650, I3379, g2242;
wire g1205, I2033, I5871, g774, g6819, g6694, g4379, g5905, g3519, I7856, g921;
wire g1551, g1742, I4752, g6488, g2254, I8594, g2814, g4289, g4658, I6756, g6701;
wire I8972, I3271, I2845, g5300, g2350, I8806, I3611, I2137, I8943, I2337, I2913;
wire g1754, g6886, g2409, g894, g1273, I5424, I6403, g6314, g4799, I9155, g2836;
wire g2212, I6763, g3860, g2967, g6825, g5440, g3710, I5523, g843, g1543, g4132;
wire g6408, g4153, I6359, g6136, g2822, I8891, I8913, I2692, g6594, g946, g1729;
wire I5551, g4802, g3962, I2154, I4189, I5499, g5151, g3158, g6806, I4706, g5875;
wire g5530, I9167, I5926, g2921, g6065, I6315, I4371, g6887, I4429, g6122, g6465;
wire g6322, g1660, g1946, g6230, g5010, g4511, I6874, g2895, g6033, key_out_16, g2837;
wire I2979, I3864, g5884, I8342, I2218, g1513, I2312, I3714, I4297, I8255, I8815;
wire g4492, I1868, I7608, I5862, g1679, g1378, g4714, I2293, g5278, g3284, I4684;
wire I8497, g3239, I6537, g3545, g2788, g6137, g5667, g6891, g1831, g1335, g3380;
wire I4791, g6337, I4309, I2828, g3832, g1288, g5566, g3853, I3736, I6612, I7161;
wire I7361, g2842, g1805, I6417, I3623, g4262, I7051, I2221, g3559, key_out_9, g4736;
wire g2485, I7451, I2703, I8267, g4623, g1947, I5885, I7999, g878, I7146, I6330;
wire I7346, I3871, I8329, g4375, g4871, I8761, g3204, g4722, g710, I4498, g829;
wire g5113, g1632, g1037, g3100, I8828, g6726, g6497, g1653, g2640, I8727, g2031;
wire I5436, g2252, g5908, g2958, I7472, g2176, I2716, I5831, I2349, g4139, I5182;
wire g5518, g5567, I5382, g2405, I2848, g1917, g2829, g2765, I7116, I4019, g4424;
wire I6090, I4362, I3672, g3040, I3077, g4809, g5593, g3440, g3969, g6312, I6366;
wire I4452, g2974, g6401, g895, I6456, g4523, g1233, I6649, g4643, g5264, I9158;
wire g1054, g5160, g2796, I6355, g2473, I3099, I8576, g1770, I8866, I3304, I4486;
wire g5521, I3499, I8716, g1725, I7596, g6727, g3875, g2324, I4504, I2119, g5450;
wire I5037, g5996, key_out_18, g4104, g6592, g4099, g4499, I2352, I6063, g6746, I2867;
wire I8699, g2177, g5179, g5379, I2893, g5878, I3044, g1189, g3839, g6932, g4273;
wire g5658, g6624, I6118, I6318, I3983, g2849, I3572, g1787, I5442, I4678, I6057;
wire I8524, I4331, I8644, I3543, I6989, I2614, g1675, I2370, I2125, g3235, g3343;
wire I5233, I2821, g4712, g985, g6576, I6549, I8258, I8818, I3534, g2245, I3729;
wire I3961, I5454, g2291, g5997, g4534, I3927, I5532, g1684, g6699, g1639, g1338;
wire g1963, I8186, I6321, I4226, g1109, g1791, I8975, I3946, g889, I2306, g3792;
wire I6625, g2819, g4014, I8426, I5412, g4660, I6253, g2088, g2923, I4173, I8614;
wire I3513, g2488, g1759, I2756, g2701, I7190, I8821, g6524, I6740, g4513, I8984;
wire I7501, g1957, g2215, g6119, I2904, g6319, g1049, g5901, g2886, I6552, I4059;
wire g4036, g3094, I4459, I8544, g4679, g6352, g6818, g6577, I1847, I3288, g3567;
wire key_out_7, I3382, g1715, g4135, I7704, g848, g5092, g1498, I2763, g2870, I3022;
wire I4261, I2391, g4382, g3776, g6893, g1833, I3422, g5574, I3749, g3593, key_out_6;
wire g6211, g2650, g5714, g932, I8061, g4805, g4022, g1584, g4422, g6599, g1539;
wire I5109, g2408, I2159, I6570, g2136, I4664, I8027, I4246, g2336, g5580, g716;
wire I3560, g736, I6525, g2768, g6370, g2594, g4798, g6325, g6821, g4560, g2806;
wire I3632, g3450, I3037, g6939, g1052, I3653, I3102, I2115, I2315, I2811, g6083;
wire g2887, I2047, g6544, I6607, g4632, g5889, g5476, g2934, g2230, g4437, g4102;
wire g4302, I5865, g6106, g4579, g4869, g6306, I3752, g5375, I8107, g4719, g1730;
wire g3289, g1504, g3777, I6587, I8159, I6111, g3835, I6311, I8223, g2096, I9143;
wire g3882, g1070, g2550, I6615, g3271, key_out_5, I4671, I2880, g2845, g1897, g6622;
wire I2537, I5896, g2195, g4265, g2891, g2913, g5139, I3364, g5384, I9134, I2272;
wire g6904, g4786, g3799, g6514, g4364, I8447, I3770, I5019, I2417, g6403, g5809;
wire I7683, g6841, g3541, I2982, g1678, g4770, g1006, I2234, g1331, g4296, I2128;
wire g3238, I3553, I6020, g3332, g5477, I6420, g6695, I2330, g3209, I6507, g4532;
wire g1682, g6107, I9113, I1856, g1305, g6536, g3802, I5728, g2481, I7475, g931;
wire g1748, g2692, I4217, g2097, I4066, g5551, g5742, g2726, g5099, g2497, I5385;
wire g5304, g2154, g1755, g4189, I8978, g4706, g6416, I8243, I8417, g3901, I6630;
wire I7646, I3675, g6522, g6115, g1045, I3281, I7039, I7484, g1173, I4455, I8629;
wire g5273, I4133, g1491, g760, g2783, g4281, g3600, g2112, g1283, g2312, g1369;
wire I6750, g6654, g3714, I7583, I3684, I5006, I8800, g1059, g1578, g2001, I5406;
wire g5572, I3109, I3791, g2293, g6880, g6595, g4138, g1535, g4639, g6537, g5543;
wire I3808, I7276, I5487, I2355, g4109, g4309, g2828, g2830, g2727, g4808, I2964;
wire g821, g6612, g5534, g5729, I6666, I9179, g1415, g4707, g6417, I7404, g3076;
wire I8512, g3889, I6528, g1664, g1246, g6234, I3575, g5885, g6328, g1203, I5445;
wire g5946, g6542, g6330, g1721, key_out_46, I5091, I8056, g2932, I8456, g5903, I3833;
wire I2318, g4715, I2367, I1924, g6800, I5169, I6410, g4098, g3500, g4498, I2057;
wire g1502, I5059, I5920, I2457, I3584, I5868, I2989, I2193, g5436, g3384, g1940;
wire g2576, g2866, g5135, g2716, g3838, I7906, I3268, I3019, g3424, g5382, I5793;
wire I3419, g6902, I6143, I6343, g846, g1671, g5805, I5415, g6512, I3452, g4162;
wire g5022, g1030, I8279, g3231, g6490, I2321, g6823, g3477, g6166, g6366, I6334;
wire I8872, g2241, g1564, I7892, I3086, g6529, I8843, g6649, I6555, g1741, I6792;
wire g3104, I3385, g2524, g2644, I8834, g6698, g1638, g839, key_out_31, I6621, g2119;
wire I5502, g1108, I3025, I2552, g5437, g4385, I3425, I9092, I4441, g2818, g2867;
wire g1883, g5579, I7478, g4425, I7035, I5388, I7517, g2893, g5752, I8232, g5917;
wire I6567, g6720, I3678, g2975, I5030, I3331, g1861, g6367, g1048, I5430, g2599;
wire g5042, g1711, key_out_43, I3635, g6652, g5442, g1055, I2570, I2860, g6057, g4131;
wire I4743, I3105, g2170, g2370, g4406, g6193, g1333, g2125, I8552, g1774, g4766;
wire g4105, g1846, g5054, g4801, g6834, g4487, I7110, g3534, I5910, g5770, I3755;
wire g5296, I8687, I6933, g2544, g6598, I5609, I4474, I2358, g3014, g6121, I7002;
wire g766, g3885, g4226, g2106, g2306, I3373, g2790, g6232, I5217, I8570, I8860;
wire I4480, g1994, g1290, I2275, g6938, I5466, g4173, I8710, g2461, I7590, I3602;
wire I3007, g2756, g2622, I3059, I3578, I3868, g5888, g1256, g6519, I6289, I9024;
wire I5448, I3767, g5787, g2904, g6552, g6606, g2446, I5333, I2284, g1381, g4718;
wire g4767, I3261, g1847, I4688, I5774, I9077, I8659, g4535, I4976, g1685, g2145;
wire I8506, g2841, g4582, g3022, g2391, g6586, g952, g1263, g964, I2420, g2695;
wire g2637, g1950, g5138, g4227, I7295, g5791, g3798, I9104, g5309, g2159, g6570;
wire g4246, I6132, I8174, g6525, g6710, I5418, I6680, g4721, g1631, g2416, g3095;
wire g3037, I3502, g1257, g1101, I2204, I2630, I5493, I8180, I4220, I7966, I8591;
wire g2315, g5957, g6879, g6607, I6558, g4502, g5049, I9044, g927, I1942, I4023;
wire g3719, g6506, g5575, I8420, I3388, g2874, g3752, I5397, I3028, g4188, g6587;
wire g4388, I5421, I3428, I2973, I7254, I7814, I3247, g3042, g6615, I7150, I4327;
wire g4428, g3786, g5584, g5539, g5896, g1673, g6374, I3826, g3364, g3233, I8515;
wire g4564, g3054, I5562, I4303, g2612, I8300, g6284, g2243, g3770, I9014, I3638;
wire g1772, I5723, g4741, g6591, g5052, g6832, g4910, I2648, g2234, g6853, g1890;
wire I3883, g6420, I4240, g2330, g4108, g4609, g6507, g4308, g1011, g1734, I3758;
wire g5086, g897, I8040, g951, I8969, g2800, g5730, g2554, g4758, I2839, I3861;
wire g6905, g3029, I3711, I9182, g3787, g2213, g5897, g5025, key_out_89, g6515, g4861;
wire g5425, I4347, I2172, I2278, g4711, g6100, I4681, g1480, g2902, I8875, I2143;
wire I2343, I6139, g4133, g3297, g2512, g2090, g4846, I2134, I6795, I6737, I2334;
wire I6809, I5743, g5331, I5890, I3509, g3963, g3791, I8884, I5505, g1688, I6672;
wire g4780, g6040, g1857, I6231, I3662, g4509, g5087, I9095, g5801, g2155, I9208;
wire g4662, I3093, g965, I3493, I3816, g1326, I8235, I6099, I8282, g3049, g6528;
wire g1760, g4493, g6351, I1850, g6875, g834, I8988, g6530, g3575, g5045, I8693;
wire g6655, g5445, I5713, g3604, I8548, g5491, g3498, g4381, g4847, g2118, g2619;
wire I8555, g2367, g2872, g1608, g1220, g4700, g6410, I9164, g4397, I9233, I2776;
wire I7640, g5407, g6884, I2593, g5059, g5920, g6839, g2457, g5578, I6444, I6269;
wire g1423, g923, I5857, I7176, g1588, I8113, g5582, g1161, key_out_126, g6278, g2686;
wire g6372, g3162, g5261, g3019, I4294, I6543, g6618, g1665, I7829, I3723, g6143;
wire g4562, g6235, g2598, g3052, g1327, I2521, I3301, g5415, g3452, g6282, I2050;
wire I5400, g6566, I8494, I4501, I6534, I8518, I3605, g4723, I8567, g4101, g6134;
wire g5664, g2625, I7270, g2232, g6548, I6927, g3086, I2724, g2253, I2179, g3486;
wire g2813, I2379, g1696, key_out_44, I7073, I7796, I6885, I6414, g3504, I6946, g1732;
wire g3881, g2740, I2658, I3441, I7069, g3070, I8264, g6621, I2835, I7469, g3897;
wire I5023, g1472, g1043, I5977, I8521, I6036, I8641, I2611, g893, g2687, I8450;
wire I3669, g1116, g2586, I3531, I5451, I6182, g6518, g6567, I8724, I6382, g996;
wire g3331, I3890, g4772, g5247, g4531, I5633, I8878, g1681, I3505, g6593, g3766;
wire g1533, g5564, I5103, g2525, g3801, g3487, g1914, I5696, g2691, g4011, I6798;
wire g4856, g5741, I2802, I3074, I3474, I5753, g5638, g6160, g3226, I5508, g6360;
wire g6933, I5944, g2962, g6521, I9098, g2158, I5472, I8981, g2506, I3080, I8674;
wire g1820, I5043, I6495, g1936, I6437, g3173, I6102, I6302, I8997, g1117, I8541;
wire g1317, g3491, key_out_10, g2587, I6579, I5116, I7852, I5316, g6724, I3569, g2111;
wire g2275, g5466, I8332, g4713, I7701, g3369, I8153, g3007, g2615, g6878, I2864;
wire g4569, g5571, g5861, g3868, g2174, g3459, g815, g1775, g5448, g1922, g835;
wire g5711, g6835, g1581, g6882, I6042, g1060, g2284, I6786, g1460, g5774, g4857;
wire g3793, g6611, g2591, g3015, g3227, g1739, I6054, g5538, I6296, I4646, I2623;
wire g4126, g5509, g4400, g1937, g6541, I9185, I2476, I7336, I8600, g2931, g4760;
wire g1294, key_out_39, I1877, g6332, g5067, g1190, I2175, g6353, g5994, I3608, g2905;
wire I6012, g6744, I3779, g6802, g2628, g1156, g2515, g5493, I7065, g5256, I6706;
wire g4220, g3940, I6371, I4276, g4423, I3161, I3361, g5381, g3388, I9131, I6956;
wire g6901, I5460, I5597, I8623, g3216, I3665, g5685, g6511, I8476, I2424, g743;
wire g862, g2973, g1954, g3030, g1250, I5739, g1363, I4986, I3999, g3247, g4127;
wire key_out_30, I3346, g5950, g1053, g2040, g6600, g6574, I2231, I1844, g2440, g3564;
wire key_out_1, g6714, I2643, g4146, key_out_99, I5668, g4633, I8285, I5840, I8500, g791;
wire g4103, g6580, I7859, g5631, g3638, g5723, I9173, I3240, g4732, g3108, g3308;
wire I6759, g2875, g4753, g4508, g917, I8809, I7342, g6623, g6076, I7081, g6889;
wire g5751, I3316, g3589, key_out_8, I7481, I3034, g3466, g2410, I7692, I3434, I4516;
wire I7497, g4116, g6375, g2884, I2044, g3571, key_out_4, g2839, g3861, g6722, g4034;
wire I7960, g852, I2269, g6651, g3448, g4565, I3681, I5053, g3455, g6285, g4147;
wire key_out_100, g6500, g2172, I2712, I9227, I5568, g4533, g3846, g2618, I3596, g2667;
wire g1683, g2343, g5168, I3013, g6339, g3196, g4914, g3803, g4210, I7267, g1894;
wire I5157, g6838, I9203, I2961, g6424, g2134, I6362, g1735, key_out_47, I8273, g6809;
wire g5890, g1782, I4340, I6452, I5929, g1661, I8044, g2555, g6231, g5011, I8444;
wire g3067, I2414, g729, g5411, g6523, g861, I2946, g2792, g1627, g4117, g1292;
wire I5626, g3093, g898, g1998, g1646, g5992, g4601, g1084, g6104, g854, g1039;
wire g1484, I3581, g6499, g1439, I9028, I8961, g4775, I6470, g5573, g3847, g5480;
wire I6425, I2831, g2494, I2182, g2518, g1583, g1702, I2382, I8414, g3263, I8946;
wire g1919, I2805, I2916, g2776, I2749, g4784, g6044, g1276, I4402, I3294, I3840;
wire I6406, I5475, g6572, I4762, I7349, I6635, g2264, g6712, g851, I6766, I6087;
wire I6105, g6543, g4840, I6305, I6801, g2360, g2933, g3723, g1647, g4190, I5526;
wire I5998, I8335, I8831, I9217, g1546, I2873, I2037, g6534, g6729, g3605, I5084;
wire I5603, g2996, I2653, I5484, I3942, g1503, I5439, I8916, g1925, I8749, g2179;
wire g6014, key_out_19, g6885, I6045, g4704, g6414, I5702, g1320, g3041, g5383, g5924;
wire g5220, I7119, g6903, g2777, g3441, g2835, I3053, I1958, g4250, g6513, g913;
wire I6283, I7258, I5952, g4810, g2882, I7352, g3673, key_out_11, I2442, g1789, g6036;
wire I8632, I2364, g980, I8653, g1771, g3772, I6582, g5051, g2981, I8579, I8869;
wire I4489, g3458, g865, I2296, g3890, g2997, I6015, g2541, I8752, I4471, I7170;
wire g6422, g2353, g4929, I4955, I3626, g2744, g909, g1738, g2802, g3074, g949;
wire g1991, g6560, I5320, g4626, g1340, I2029, I9021, g3480, g1690, g6653, g6102;
wire I2281, I7061, I7187, g6579, g5116, I5987, g5316, g1656, I6689, g5434, g2574;
wire g2864, g4778, g855, g5147, I3782, g4894, I2745, I8189, I4229, I6430, g3976;
wire I2791, I6247, I7514, I2309, I9101, g1110, I8888, g2580, g5210, g6786, I6564;
wire I8171, I2808, I8429, g5596, g6164, g6364, g6233, I5991, I2707, g4292, I7695;
wire I7637, g2968, I5078, g1824, g4526, I5478, g1236, key_out_120, I7107, I5907, g6725;
wire g1762, g2889, I6108, g4603, g6532, I6308, I5517, I9041, I2449, g4439, g5117;
wire g6553, g4850, I8684, I5876, I8745, g2175, g2871, I2604, g3183, g2722, I4462;
wire I8309, g1556, I6066, g3779, g1222, key_out_124, g4702, g6412, g896, g3023, I7251;
wire g1928, I7811, g6706, g5922, I8707, g1064, I2584, I5214, g6888, g1899, I6048;
wire g5581, I6448, g6371, g4276, I4249, g5597, I3004, I1825, g4561, g2838, I3647;
wire g3451, I2162, g1563, I9011, I4192, g2809, I3764, g5784, I3546, I5002, g4527;
wire g4404, g1295, g4647, g3346, I5236, g2672, g2231, g4764, g5995, key_out_17, I9074;
wire g5479, g2643, I6780, g6745, g1394, g4503, I7612, g1731, I2728, g1557, g2634;
wire g1966, g4224, I5556, I2185, g2104, g2099, g3240, I2385, g6707, g1471, g4120;
wire I4031, g4320, I4252, I3617, I3906, I6093, I8162, g3043, g971, I5899, I4176;
wire I6816, I3516, g2754, g4617, g3034, g1254, g1814, g6575, g4516, g6715, g4771;
wire g2044, I6685, g5250, g6604, g1038, I6397, g6498, g1773, I2131, g5432, g4299;
wire g6833, I8730, g5453, I4270, g2862, I2635, g2712, I8881, I5394, g1769, g3914;
wire g6584, I1859, g6539, g6896, g1836, g5568, I8070, I5731, I8470, I8897, g1918;
wire I3244, I7490, I4980, g5912, I4324, I3140, g2961, I5071, I3340, I5705, g6162;
wire I3478, g6362, g6419, I6723, g4140, g6052, g2927, I5948, I9220, g2885, I7355;
wire I8678, I2445, g2660, g2946, g938, g4435, I2373, g4517, I7698, I3656, g3601;
wire I2491, g2903, I8635, g6728, g6486, I2169, g942, g6730, I9161, g3775, g6504;
wire g3922, I7463, I2578, g6385, g6881, I5409, g2036, g706, I6441, g4915, g2178;
wire g2436, g2679, g6070, g2378, g3060, I3310, g6897, g1837, I8755, g3460, I8226;
wire g6425, g2135, I4510, I9146, g4110, I7167, I7318, I4291, g5894, g2805, g910;
wire g1788, g2422, I6772, I7193, I8491, g3079, I6531, g4402, g784, g1249, g4824;
wire g837, g5661, g3840, g719, I3590, g6406, g5475, I7686, g1842, I2721, g1192;
wire I8459, g6105, g6087, g6801, g6305, g5292, I8767, g6487, I3556, g3501, I3222;
wire I8535, g4657, I8582, g1854, I9116, I8261, g5084, g4222, g2437, g2653, I6992;
wire I1932, g2102, g5439, I3785, I2940, I5837, g2869, I2388, I6573, I3563, g5702;
wire I8246, g1219, g1640, g2752, g6373, g3363, g6491, g5919, I2671, g1812, I8721;
wire I2428, g4563, g3053, g1176, g2265, g3453, g6283, g6369, g2042, g6602, I5249;
wire g6407, g6578, g4844, g2164, g1286, g2364, g2233, g4194, g1911, g4394, g6535;
wire I6976, g3912, I2741, g5527, g6582, I8940, g4731, I2910, I3071, g5647, I3705;
wire I3471, g2296, g1733, I2638, g1270, g5546, I5854, I4465, g6015, g4705, g6415;
wire I6126, I6400, g4242, I2883, I8671, g5925, I8030, I4433, g1324, I5708, I5520;
wire g6721, I5640, g5120, I8564, g2706, I5252, I3773, g1177, key_out_125, g4150, I2165;
wire g1206, g4350, g2888, I7358, I4195, g2029, I7506, I5376, g2171, I4337, I8910;
wire g2787, g6502, g2956, I6023, I8638, g1287, g2675, I3836, I3212, I7587, g6940;
wire g4769, g1849, g3778, g6188, I2196, g5299, g1781, I6051, g1898, g3782, I8217;
wire I8758, I8066, g5892, I6327, g6428, g3075, g4229, g2109, I7284, I4255, I6346;
wire I8165, g4822, g1291, I5124, I2067, g6564, I5324, I7832, g6826, I5469, I2290;
wire g1344, I4354, g5140, I5177, g3084, g5478, g1819, I6753, g2957, I8803, g1088;
wire g1852, I6072, g6609, g5435, g6308, I3062, g5082, g2449, I3620, I3462, I8538;
wire g2575, g2865, g6883, g5876, g4837, I8509, I2700, g2604, I4267, g2098, I4312;
wire g4620, g4462, g6589, g945, I8662, I3788, g6466, g5915, g3952, I6434, I8467;
wire I8994, I8290, g1114, g6165, g6571, g6365, g2584, g4788, g6048, I1841, g6711;
wire I8093, g5110, g4249, g5310, I3298, g1825, g6827, g1650, I3485, g3527, g809;
wire I6697, g4842, g849, g2268, g4192, g4392, g3546, key_out_3, g4485, I2817, g5824;
wire g1336, g6803, g3970, g1594, g4854, g6538, g1972, I5923, g6509, g1806, g5877;
wire g5590, g1943, I3708, g3224, g2086, g2728, I3031, I4468, g3320, g6067, g1887;
wire I3431, g1122, g6418, g6467, g1322, g4520, g1934, I2041, I3376, g4431, g4252;
wire I1874, I3405, g3906, g2470, g3789, g5064, g2025, g6493, g5899, I6775, g4376;
wire g4405, g3771, I5825, g872, g1550, I6060, g4286, g4765, I1880, I4198, g3299;
wire g5563, I4398, g4911, I3733, g6700, g1395, g1891, g1337, g5237, g3892, g2678;
wire I3225, g6421, I2890, I8585, I5594, g4270, I7372, g1807, g4225, g2682, g2766;
wire I6995, I1935, g2087, g2105, I6937, I7143, I8441, g2801, I2411, g5089, g5489;
wire I5065, g4124, g714, I3540, g4980, g2748, g6562, I3206, g5705, I2992, g3478;
wire g1142, g2755, I4258, g5242, I8168, g6723, g1255, I5033, g6101, g6817, I5433;
wire g4206, g3082, g3482, I8531, g1692, key_out_48, g6605, g1726, key_out_45, g3876, g2173;
wire I6942, g2091, I5496, g1960, g2491, g5150, g4849, g2169, g2283, I7113, I8411;
wire I5337, I5913, g2602, g6585, g2007, g5773, g4399, I3797, I6250, g2059, g2920;
wire I4170, g4781, g6441, I8074, g2767, g4900, g1783, g3110, I4821, I2688, I2857;
wire g2535, I3291, g1979, g1112, g1267, I7494, g4510, I3144, g5918, g1001, g3002;
wire I8573, I8863, I4483, g1293, g6368, g4144, key_out_98, I8713, I7593, I3819, g3236;
wire g1329, I3694, g1761, g857, g5993, g6531, I5081, I3923, I4306, I2760, g2664;
wire I5481, I3488, g6743, g6890, g1830, I5692, I7264, g4852, g6505, I3215, g1221;
wire g6411, g6734, g3222, I3886, I8857, g1703, key_out_41, I2608, g5921, g4215, I2779;
wire I7996, g6074, g3064, g3785, g1624, g1953, I4003, g5895, g4114, g4314, I2588;
wire I3650, g6080, I2361, g6573, I4391, g6713, I3408, g3237, I7835, I2327, g6569;
wire g2030, g5788, g2430, I2346, g4136, I8183, I4223, I8220, g4768, g1848, I9140;
wire g2826, g1699, key_out_42, g1747, g838, I6075, I2696, I4757, I7799, I3065, g3557;
wire I5746, g4806, g5392, I8423, I9035, I6949, g4943, I3465, I3322, I9082, g3705;
wire I8588, I4522, I2753, g842, I6292, I4315, g3242, g4122, g4228, g4322, I2240;
wire I1938, g2108, g2609, I6646, g2308, I8665, I8051, I7153, g2883, I6084, I6039;
wire I5068, I3096, g1644, I3496, g715, I3550, I7802, g5708, g1119, g1319, g2066;
wire g3150, g5219, I3137, I8103, I3395, I3337, g4496, g1352, I9110, g1577, g4550;
wire g3773, g4845, I4537, I8696, g2165, g5958, I2147, g6608, g4195, g4137, g830;
wire I5716, g3769, I9002, g2827, I6952, I5848, g3836, g3212, g6423, I4243, g2333;
wire I8240, g1975, I5699, g4807, I9236, g3967, I6561, g6588, I4935, I2596, g6161;
wire g1274, g6361, g1426, g2196, I7600, g2803, I6004, g3229, I6986, g6051, key_out_14;
wire g5270, g804, I3255, g2538, g1325, g1821, g844, I3481, I8034, g4142, key_out_93;
wire g4248, g2509, I6546, I3726, g4815, I5644, I8147, g5124, g6103, I5119, g4692;
wire g2467, I8681, g4726, g5469, g4154, I2601, g6696, g1636, g3921, g5540, I5577;
wire g1106, g6732, g853, g2256, g1790, I2922, g6508, I5893, I3979, I2581, I3112;
wire g1461, g3462, g1756, g2381, I6789, g4783, g6043, key_out_15, I7871, I2460, I3001;
wire g4112, g4218, g2197, g4267, I4166, g2397, I4366, g5199, g5399, g1046, I3761;
wire g3788, g6034, key_out_13, g6434, g6565, I6299, g4293, g4129, g5797, I3830, I2995;
wire g6147, g1345, g1841, g6347, I1832, I2479, I7339, g1191, I2668, g1391, I1853;
wire g3192, g6533, g3085, I3746, I7838, g4727, I4964, g3485, I2190, g1695, g6697;
wire g1637, g1107, g2631, g6596, g3854, I5106, I8597, g2817, I6244, I7077, g4703;
wire g6413, I5790, g1858, I6078, I6340, I7643, I3068, g5923, I9038, I3468, I4279;
wire I5756, g6820, g4624, I6959, I5622, g3219, I5027, I4318, I7634, I5427, g3031;
wire g1115, g6117, g1315, g1811, g1642, I8479, g2585, I7104, I5904, I8668, g5886;
wire I8840, g2041, g6601, I5514, I3349, I2053, g5114, I5403, g5314, I2453, g1654;
wire g4716, g4149, key_out_92, g6922, I8156, I3198, I3855, I5391, g3911, g6581, g4848;
wire I5637, g1880, g4198, g4699, g6597, g4855, g4398, g2772, I4321, g5136, g3225;
wire I5223, g2743, g6784, g2890, g3073, g1978, g3796, g1017, I2929, g798, g2505;
wire I3644, g3124, g1935, g3980, g2856, g2734, I8432, I3319, g1982, g754, g4524;
wire g836, I8453, g6840, I4519, g4644, I3152, I3258, g3540, I3352, g1328, g5887;
wire g4119, g5465, g1542, g1330, g3177, I3717, g5230, g845, g4152, g6501, g4577;
wire g4717, g5433, I5654, I6930, g2863, I6464, I3599, g2713, I3274, g4386, g3199;
wire g5550, I3614, g3781, I3370, g5137, g5395, g5891, g3898, g3900, I3325, g4426;
wire key_out_102, I2735, g3797, I9085, g1902, g6163, g4614, I2782, I7679, g6363, g4370;
wire I8626, g3510, I5612, g6032, g4125, g2688, g2857, g3291, I3083, g2976, g1823;
wire I2949, g1366, g5266, I2627, g1056, g6568, I5328, g1529, I7805, I5542, I2998;
wire g1649, g1348, g3259, I4358, g5248, g4636, g1355, g4106, g5255, g3852, I9031;
wire g2760, g3488, I8894, g4790, g5692, I4587, g5097, g5726, g4187, I9176, g4387;
wire I9005, g1063, g3886, g4622, g2608, I2919, g2779, g4904, g3114, I2952, g1279;
wire g4514, g1720, g4003, g1118, I3391, g1318, g4403, I5490, g5112, g2588, g4145;
wire key_out_97, g4841, I8603, g2361, I6769, g4763, g4191, g4391, I5056, I2986, I3307;
wire g1193, key_out_127, I5529, I4420, I5148, g3136, g2327, I6918, I4507, g5329, g1549;
wire g4107, I7042, g947, g6894, g1834, I4794, g4307, I5851, g4536, I3858, I8702;
wire g2346, g6735, I3016, I2970, g5727, I7164, g2103, g858, I2925, g4858, I3522;
wire g4016, I3115, I3251, I3811, I8276, g1321, I3047, g1670, g3228, g3465, g3322;
wire I5463, g3230, g4522, g4115, g2753, g4251, g1232, I4300, g6526, g1813, I8527;
wire I8647, I2617, I5720, g2043, g6039, key_out_20, I8764, g2443, g6484, g3096, g5468;
wire g1519, g1740, I7012, g6850, I6895, I1835, g3845, I5843, g2316, I3537, I8503;
wire g1552, I5457, g2565, g6583, g850, g5576, g4537, I7029, g2347, I5686, I4123;
wire g3807, g1586, g3859, g6276, g4612, g2914, g6616, I3629, g6561, I3328, I2738;
wire I8617, g1341, g2413, I4351, g3342, g4128, g1710, g4629, I6485, g6527, g6404;
wire g4328, I2140, g1645, I2340, g4130, I5938, I7963, I3800, g3481, I2907, g2820;
wire g2936, g5524, g6503, g3354, I4410, I7808, g2117, g3960, g2317, g5119, g6925;
wire I7707, I5606, g1659, g1358, g5352, g5577, g4213, g5717, I3902, g6120, g2922;
wire g1587, I6812, I8991, g3783, g1111, I3090, I9008, g5893, g1275, g6277, g2581;
wire I3823, g3267, key_out_2, I4667, g3312, I7865, I4343, g2060, g6617, g6906, g5975;
wire g4512, I4282, g2460, I7604, I8907, I3056, g3001, g1174, g4823, I2663, g4166;
wire g6516, g5274, I8435, I3148, I8690, g1985, I4334, I8482, g2739, g3761, I3155;
wire I3355, I2402, g4529, g1284, g4148, key_out_96, I6733, I8656, g3830, I9122, g2079;
wire g4155, g4851, g6892, g1832, I9230, g1853, g2840, I2877, I5879, g5544, g2390;
wire I6324, g1559, I6069, I8110, g4463, g943, g1931, g6709, g3932, I6540, I3720;
wire g6078, I1871, I6377, g5061, g6478, I2464, I3367, g5387, I9137, g1905, I8002;
wire g866, I2785, I7086, I5615, g6035, key_out_21, g4720, I3843, g4118, g4619, g6517;
wire g1204, g3677, g6876, g4843, g3866, g2954, I4593, g5046, g2163, g6656, g4193;
wire I2237, g2032, g4393, I5545, g5403, I1838, g3848, I5591, I4264, I2394, g5391;
wire g2568, I2731, I4050, g3241, g2912, g4121, g1969, I3232, g4321, g5307, g2157;
wire g5536, g2357, g1123, key_out_122, g1323, g4625, I3909, g4232, g6402, g6824, g1666;
wire g4938, I6819, g6236, I3519, I8295, I2955, I7487, g856, I6923, g1528, I5204;
wire I5630, I6488, g1351, g1648, I2814, g1875, g4519, g5115, g6590, g5251, g6877;
wire g3258, I4777, I6701, g5315, g3867, I2150, g1655, g6657, g4606, I3687, I8089;
wire I2773, g5874, g1410, I8966, I5750, I7045, I6114, g3975, I7173, g1884, I7091;
wire g6899, I4799, I2212, g929, g6785, g5880, I5040, I2967, g5537, g2778, I1862;
wire I3525, g3370, g2894, I7007, g1372, g4141, g6563, I6008, I3691, g4525, g1143;
wire key_out_123, g3984, I8150, g1282, I8438, g3083, g1988, I4802, I6972, g3483, I7261;
wire g6194, g1334, I3158, I3659, I3358, g5328, I1927, g6489, g5542, g5330, key_out_38;
wire g3306, g2998, g4158, g4659, g1555, key_out_113, g3790, I3587, g1792, g2603, g2039;
wire g3187, g2484, g3387, g3461, g4587, I6033, g5554, g3622, g4111, I8229, I9149;
wire I2620, g1113, I4492, g4615, g2583, g3904, g3200, I6096, g3046, g899, g4374;
wire I3284, g2919, g1908, I2788, g1094, I5618, g2952, I6337, I5343, g2276, g1567;
wire g4284, g5512, g4545, g5090, g6409, g5490, I7689, g4380, I2842, g1776, g1593;
wire g2004, g4853, g6836, I2485, I3794, g2986, g4020, g6212, I5548, g5456, g2647;
wire I8837, g5148, g5649, g4507, g3223, I4623, I1947, g2764, I8620, I8462, I9119;
wire I2854, g4559, g5155, g5355, I9152, g3016, g6229, g1160, g5260, I6081, I4375;
wire g6822, g1641, g3251, I6692, g1450, g5063, I7910, I8249, g4628, g4515, g2120;
wire I4285, g2320, g4100, g1724, g3874, I2958, I5094, I2376, I8485, g5720, I2405;
wire g2906, g2789, g1878, g5118, I9170, I1917, g2771, g6620, g5193, I5360, g5598;
wire g6249, g4666, g3629, g3328, g6085, g4351, g4648, g5232, g2340, g5938, g5909;
wire g1802, g3554, g4410, g6640, g4172, g4372, g3512, g3490, g4667, g3166, g3366;
wire g6829, g3649, g6911, g3155, g3698, g6270, key_out_54, g4792, g6473, g4621, g5158;
wire g6124, g6324, g6469, g3279, g3619, g3167, g5311, g3367, g3652, g3843, g4593;
wire g3686, g5180, g5380, g4160, g3321, g2089, g6245, g4360, g3670, g3625, g6291;
wire g4050, g5559, g6144, g6344, g2948, g6259, key_out_51, g4179, g2955, g6088, g6852;
wire g6923, g5515, g1499, g4835, g3687, g4271, g4611, g3341, g6650, g4541, g3645;
wire g5123, g3691, g4209, g4353, g6336, g6768, g4744, g3659, g5351, g3358, g5648;
wire g6934, g3275, g3311, g5410, g3615, g2062, g3374, g4600, g6096, g1436, g5172;
wire g3180, g5618, g5143, g6913, g5235, g4580, g2085, g6266, key_out_55, g5555, g2941;
wire g6248, g6342, g5621, g3628, g6255, g6081, g3630, g6692, g3300, g6154, g6354;
wire g4184, g5494, g4384, g4339, g4838, g3123, g3323, g4672, g2733, g3666, g6129;
wire g6329, g2073, g5360, g6828, g5050, g3351, g6830, g3648, g3655, g1706, g6068;
wire key_out_66, g4044, g6468, g3172, g3278, g3372, g2781, g3618, g3667, g3143, g3282;
wire g6716, g6149, g3693, g3134, g3334, g6848, g5153, g5209, g5353, g6241, g1808;
wire g3113, g5558, g6644, g6152, g6258, g4178, g1575, g4378, g4831, g4182, g5492;
wire g5600, g6614, g4947, g3360, g6125, g1419, g3641, g4873, g4037, g3724, g4495;
wire g3379, g5175, g3658, g6061, key_out_69, g5500, g3611, g2137, g4042, g5184, g4442;
wire g4164, g2807, g5424, g6145, g2859, g3997, g4054, g6345, g3132, g3680, g6637;
wire g3353, g2142, g2255, g6159, g2081, g3558, g5499, g4389, g4171, g6315, g4371;
wire g4429, g4787, g6047, key_out_63, g6874, g2267, g5444, g5269, g1407, g4684, g4791;
wire g6243, g6935, g2746, g4759, g6128, g5414, g6130, g5660, g3375, g4449, g3651;
wire g4865, g2953, g2068, g3285, g4833, g5178, g5679, g5378, g3339, g1689, g5182;
wire g2699, g2747, g6090, g4362, g3672, g4052, g3643, g4452, g6056, key_out_70, g1826;
wire g6148, g6348, g5560, g3634, g6155, g6851, g3551, g3099, g3304, g4486, g3499;
wire g4730, g5632, g5095, g6260, key_out_50, g4185, g1609, g5495, g2577, g3613, g6619;
wire g6318, g2026, g5164, g5364, g5233, g2821, g3729, g5454, g5553, g6321, g3660;
wire g6625, g4045, g4445, g6253, g4373, g5189, g4491, g6909, g4169, g5171, g4369;
wire g3679, g4602, g5371, g3378, g5429, g4407, g5956, g4868, g5675, g3135, g4459;
wire g3335, g3831, g3182, g3288, g3382, g4793, g4015, g2107, g6141, g6341, g6645;
wire g3632, g3437, g3653, g5201, g3208, g3302, g6158, g5449, g5604, g5098, g5498;
wire g1585, g6275, key_out_56, g6311, g4671, g4247, g3454, g4826, g5162, g5362, g3296;
wire g5419, g3725, g2935, g5452, g6559, g5728, g5486, g5185, g3171, g3371, g6628;
wire g4165, g4048, g4448, g3281, g4827, g4333, I2566, g2166, g3684, g4396, g3338;
wire g2056, g5406, g3309, g5635, g5682, g5487, g6123, g6323, g3759, g5226, g6151;
wire g3449, g6648, g5173, g5373, g4181, g2720, g4685, g5169, g5369, g5602, g2834;
wire g3362, g6343, g2121, g2670, g6693, g1633, g6334, g3728, g6555, g3730, g2909;
wire g4041, g3425, g6313, g5940, g4673, g5188, g6908, g5216, g6094, g4168, g4368;
wire g5671, g3678, g5428, g4058, g3635, g2860, g3682, g3305, g5910, g3755, g2659;
wire g5883, key_out_68, g3373, g5217, g4863, g3283, g3602, I2574, g5165, g6777, g3718;
wire g3767, g4688, g1784, g2853, g6799, g2794, g3203, g6132, key_out_49, g6238, g6153;
wire g4183, g4383, g6558, g5181, g3689, g4588, g5197, g4161, g4361, g3671, g4051;
wire g6092, g4346, g2323, g5562, g3910, g3609, g6262, g6736, g3758, g4043, g3365;
wire g5441, g5673, g4347, g3133, g3333, g3774, g4697, g3780, g6737, g6077, key_out_64;
wire g3662, g6643, g3290, g6634, g3816, g2113, g6099, g6304, g3181, g3381, g3685;
wire g3700, g3421, g5569, g4460, g4597, g6613, g4739, g6269, g4937, g4668, g3631;
wire g2160, g4390, g3301, g4501, g4156, g4356, g4942, g5183, g4163, g5023, g4363;
wire g4032, g4053, g4453, g5161, g3669, g5361, g3368, g6135, g5665, g6831, g5451;
wire g6288, g4157, g4357, g5146, g6916, g5633, g3505, g6749, g6798, g5944, g5240;
wire g5043, g5443, g6302, g6719, g2092, g4683, g5681, g3688, g4735, g6265, g4782;
wire g4661, g4949, g3326, g6770, g3760, g5936, g4039, g5317, g3383, g5601, g3608;
wire g3924, g4583, g3161, g2339, g3361, g4616, g3665, g3127, g3327, g3146, g3633;
wire g5937, g3103, g3303, g5668, g6338, g5190, g5501, g2551, g5156, g5356, g4277;
wire g5942, g4789, g3316, g3434, g5954, g5163, g6098, g3147, g5363, g3681, g5053;
wire g3697, key_out_101, g5157, g5357, g4244, g4340, g3936, g3117, g3317, g4035, g918;
wire g6086, g4214, g1620, g3784, g2916, g3479, g6131, g3668, g6331, g4236, g3294;
wire g5949, g3190, g6766, g3156, g3356, g5646, g2873, g6748, g5603, g5484, g4928;
wire g3704, g4464, g4785, g6091, g3810, g5952, g5616, g6718, g6767, g3157, g3357;
wire g4489, g2770, g4471, g5503, g3626, g4038, g5617, g3683, g4836, g2138, g3661;
wire g6247, g3627, g5945, g2808, g3292, g3646, g2759, g6910, g3603, g3484, g5482;
wire g3702, g6066, key_out_65, g5214, g3616, g6055, key_out_67, g6133, g5663, g6333, g2419;
wire g3764, g5402, g5236, g4708, g5556, g4219, g3277, g3617, g6093, g2897, g6256;
wire key_out_53, g4176, g6816, g4829, g6263, key_out_52, g5194, g3709, g5557, g3340, g6631;
wire g3907, g4177, g5948, g4377, g3690, g5955, g5350, g4199, g5438, g2868, g3310;
wire g4797, g5212, g3663, g2793, g2015, g4344, g5229, g6772, g3762, g4694, g3657;
wire g2721, g4488, g4701, g3928, g6474, g3899, g3464, g5620, g4870, g3295, g2671;
wire g1576, g3844, g1716, g3089, g3731, g3489, g5192, g5485, g5941, g4230, g6126;
wire g6326, g4033, g3814, g2758, g3350, g2861, g6924, g5176, g4395, g5376, g5911;
wire g2846, g6127, g6327, g5225, g4342, g6146, g6346, g2018, g4354, I5352, g5177;
wire g6240, g3620, g1027, g2685, g2700, g2021, g6316, g5898, g4401, g1514, g5900;
wire g2950, g4761, g5245, g1763, g4828, g3298, g4830, g5144, g4592, g6914, g2101;
wire g5488, g4932, g1416, g5701, g6317, g5215, g5951, g4677, g3176, g3376, g3286;
wire g3765, g4349, g6060, key_out_71, g1595, I5359, g3610, g6739, g1612, g3324, g6079;
wire g5122, g3377, g4352, g4867, g6156, g3287, g5096, g4186, g5496, g6250, key_out_57;
wire g4170, g4280, g3144, g3344, g5142, g3819, g6912, g3694, g6157, g5481, g3701;
wire g5497, g5154, g5354, g4461, g4756, g4046, g5218, g3650, g4345, g3336, g3768;
wire g4159, g4359, g3806, g4416, g3887, g3122, g2732, g4047, g6646, g3433, g5953;
wire g6084, g6603, g4874, g5677, g3195, g3337, I4040, g5149, g5349, g5198, g5398;
wire g1570, g6647, g1691, g3692, g3726, g3154, g4800, g5152, g6320, g5211, g5186;
wire g5599, g4490, g3293, g6771, g3329, g5170, g4456, g6299, g4348, g3727, g2937;
wire g4355, g5939, g2294, g4698, g5483, g3703, g6738, g2156, g6244, g2356, g6140;
wire g3953, g6340, g5187, g1628, g4167, g6082, g4367, g4872, g4057, g5904, g5200;
wire g4457, g5446, g3349, g2053, g5145, g6915, g4834, g4686, g5191, g3699, g4598;
wire g5637, g5159, g5359, g4253, g3644, g3319, g3352, g5047, g5447, g4687, g3186;
wire g3170, g3614, g3325, g4341, g2782, g6295, g3280, g5017, g4691, g5935, g2949;
wire I5351, g5234, g3636, g2292, g6089, g6731, g6557, g4358, g2084, g2850, g5213;
wire g6254, g6150, g5902, g3145, g3345, g6773, g3763, g3191, g4180, g5166, g3637;
wire g4832, g6769, g3307, g3359, g4794, g3757, g3522, g3315, g3642, g3654, g5619;
wire g5167, g3880, g4440, g3978, g6788, g3935, g3982, I8376, g5625, g6298, g6485;
wire g4655, g6252, g6176, I8377, g6286, g3851, g3964, g5659, g2928, g6287, g3989;
wire g5374, g3971, g6781, g3598, g4641, g4450, g3740, I8136, g5628, g5630, g6114;
wire g5323, g5666, I8137, I8395, key_out_119, g3879, I9057, g4092, I8081, g4864, g6845;
wire g5372, g5693, g5804, g6142, I8129, g6481, g4651, g4285, g4500, g5202, key_out_87;
wire g3750, g6267, g4231, g6676, g6293, g4205, g4634, I8349, key_out_121, g6703, g3884;
wire g4444, g4862, I8119, g3988, g5674, g6747, g6855, I8211, I8386, g5680, g4946;
wire I8370, key_out_117, g4436, I8387, key_out_118, g6274, g6426, g6170, g3996, I8345, g5623;
wire g6483, g4653, g3878, g6790, I8359, g4752, g6461, g3981, g5024, g4233, g4454;
wire g5672, g5077, g5231, g6307, g3744, g6251, g6447, I8128, g3864, g5044, g4745;
wire g6272, g5014, g3871, I7970, I8348, g6554, I7987, g5916, I8118, I8367, g6456;
wire I8393, g4086, g1589, g6118, g6167, g3862, g6457, g4635, g6549, g6686, g5532;
wire g6670, g5012, g4059, g5281, I8358, g6687, g3749, g5808, g6691, g3873, g3869;
wire g6659, g4430, g6239, g6545, g4638, g6794, g6931, g3990, g5385, g3888, g5470;
wire g6300, g4455, g6750, g5678, g3745, g6440, g3865, g3833, g4021, g3896, g5535;
wire g5015, g4631, g5246, g6792, I7980, I8360, key_out_94, g4441, g6113, g5388, I8379;
wire key_out_116, g5430, g4458, g3748, g6264, g4074, g6450, g4080, g5066, g6179, I8209;
wire g6289, g6658, g6271, g5662, g5018, I7972, g5467, g5816, g5700, g4451, g6864;
wire g5817, g3883, g5605, I9059, key_out_115, g4443, g4434, g5669, g5368, I7979, g5531;
wire g5458, g6795, g4936, g5074, g5474, g6926, g6754, g6273, g6444, I8378, I8135;
wire g5326, I9066, key_out_114, g6927, g3751, g6660, g6679, I8208, g6182, g5327, g3743;
wire g3856, g5303, g5696, g3992, g5472, g3863, g6437, g6917, g3857, g5533, g5697;
wire g5013, g4627, g6454, g6296, g4646, I8138, g6189, g3977, I9058, g6787, g5060;
wire g6297, g3999, g6684, I7978, g6109, g6791, g6309, g3732, g3533, I8385, g6268;
wire g3820, g6452, g5626, g4656, g6185, g3739, I7989, g3995, I8369, I7971, g5627;
wire g6682, g3942, g5583, g6173, g3954, g6920, g6261, g6793, g4948, g6246, g5224;
wire g5277, g4438, g4773, g6689, g3998, I8774, g3850, g6108, g6758, g2896, g6455;
wire g3986, g6846, g3503, I7969, g4941, g6290, g3987, g6847, g6685, g5295, g4473;
wire g3991, I7988, g5471, I8368, g6257, g6301, g6673, I8080, g6669, g3877, I8126;
wire g5062, g6480, I8779, g6688, g5085, I7981, I8127, g4433, I8346, g5812, g4859;
wire g6665, g5473, I8347, g6303, g5069, I9064, g4497, I8210, g5377, g3837, g6116;
wire I8117, g4001, g3842, g5291, g3941, g5694, g6936, g4068, I8079, g4468, g4866;
wire g3829, I8356, g3733, g6937, g6479, g6294, g5065, g5228, I8357, g3849, g6704;
wire g4599, g6453, g4544, I8778, g2924, g4427, g4446, g3870, g6683, g5676, g4637;
wire g3972, g6782, g6661, g4757, g6292, g4811, g4642, g4447, g5624, g5068, g4654;
wire g3891, g3913, I7990, g6702, g6919, I8120, g4243, g5699, g5241, g4234, g3815;
wire g5386, g6789, I8082, g5370, g3828, I9065, g3746, g5083, g6907, g5622, g6690;
wire g6482, g4652, g4549, g3747, g3855, g5695, g6110, g6310, g5016, g6762, g4740;
wire I8394, g6556, g6930, g3599, g3821, g4860, g6237, g4645, g6844, I8773, g5629;
wire g4607, g6705, g5800, g6242, g3841, g6918, g5348, g3858, g5698, g4630, g6921;
wire g5367, g1777, I7217, I7571, g5686, I2073, I2796, g948, I4205, I3875, g3330;
wire g4151, g2435, I5658, g1558, I4444, I5271, I2898, I2797, I2245, I3988, g1574;
wire g3529, I1963, I5209, key_out_72, I7562, g5506, g5111, I4182, I6186, key_out_75, I7441;
wire I6026, I2768, I3933, g5853, g2731, g5507, g2966, I2934, I3179, I6187, key_out_73;
wire I6027, g2009, I4233, g2769, g1044, key_out_106, g4674, I7569, I6391, g3525, g4680;
wire I2081, I8195, g1534, I2497, g939, I5269, key_out_22, g3985, g1036, key_out_108, I2676;
wire g1749, g6097, g6783, g5776, I7434, g1042, key_out_109, I7210, g3530, I6964, I5208;
wire key_out_78, I5302, g5777, g4613, I2544, g1138, I1994, I4445, I2061, I5189, g4903;
wire I3178, I4920, g2951, g3518, I2003, g6717, I3916, g5864, g2008, I5309, I7432;
wire I4203, g3521, I5759, I6962, I6659, key_out_33, I4940, I2935, g2266, I2542, I3412;
wire I3189, g5634, I3990, g2960, g5926, g3511, I7439, I2090, g5862, I9050, I5766;
wire key_out_34, g1582, g1793, g3968, key_out_110, I7527, I5226, key_out_29, g4049, I7224, I5767;
wire key_out_77, I5535, I5227, g5947, g3742, g5873, g4504, I7244, g5869, I5188, key_out_60;
wire g3983, key_out_105, g4678, g6843, g3961, I5308, I2506, I3445, g2061, I3169, g6740;
wire I7556, g4007, I5196, key_out_76, I7563, g5684, I2507, I1995, g2307, I7237, g2858;
wire g2757, I6744, I4183, I7557, I2300, I3188, g5865, I5197, key_out_74, I4161, I3741;
wire g5019, I5257, key_out_27, g3532, I2528, I5301, g1743, g1411, g3012, g5504, I6175;
wire I3455, I6500, g1573, I3846, I4210, g4803, g3109, g2698, g3957, I6499, key_out_91;
wire g4816, I3847, I7520, I4784, I1952, g3539, I8202, I1986, I2933, I5760, g4301;
wire I1970, I7225, I6660, g5502, I3168, I1987, g1316, I2674, g4669, I3411, I7245;
wire g2607, g5308, g2311, g3535, g5455, I4782, I9052, I3126, I3400, I4526, g5780;
wire g3246, g3502, g4608, I4919, g2100, I7230, I7433, I3127, g3028, I2795, I5784;
wire I4527, I7550, I4546, I6745, I5294, I6963, g3741, g1157, I2499, g937, g4472;
wire g2010, g928, I7097, I4547, I3697, I3914, I2543, I3413, I7218, I7312, g3538;
wire g5505, g1075, I2014, g2804, g6742, I6185, key_out_36, g5863, I3739, I2022, I5782;
wire I7576, g5688, g5857, I3190, I5292, g1764, I3954, g5779, I7577, I5647, g3531;
wire I1980, g5508, I4150, g6873, g6095, I4009, I2675, g926, I3894, I4212, g5565;
wire I6028, I2109, I5244, g1402, I4921, I7536, I7223, I2498, I1951, I7522, I3952;
wire g5775, I8201, g2024, g2795, g4004, I6196, I3970, I4941, I5657, I7542, I2897;
wire I2682, I2766, g3013, I5242, key_out_28, I7529, g1822, I3876, I2091, I3915, I9051;
wire I2767, I1979, g3597, g2831, g5683, g5778, I2015, g930, g5782, g4002, I2246;
wire I6743, I7549, g2947, g4762, g2095, g944, I6474, I7232, I1953, g2719, I8203;
wire I4008, g4237, g1829, g901, g941, I7570, I2108, g1540, g4814, I7311, I5270;
wire g2745, g1797, g2791, I7239, g3526, g6741, I8196, I3895, I4783, I2021, g905;
wire g3276, g6774, I5207, key_out_37, I2301, I5259, I7440, I7528, g4640, g4812, g1845;
wire g6397, I5768, key_out_88, I1978, g4610, I5228, I2074, g3140, I6390, key_out_59, I3177;
wire I4152, I6501, key_out_90, I7548, g1815, I7555, g3517, I2080, key_out_24, I4211, I3399;
wire I5195, key_out_35, I7313, g2582, I4939, g950, g4819, I7521, I2023, I4446, I5783;
wire g2940, g4825, I5293, I5761, I1971, I3972, I4159, I6661, key_out_62, g1398, I6475;
wire I3934, I7541, I2508, g5854, g4465, I2072, key_out_25, I7238, g3955, I7209, g5431;
wire I2681, I2013, I4234, g2780, g2067, I1962, I5258, g1387, I2060, key_out_26, g5781;
wire g2263, g4221, g1359, I7231, I3953, I5187, key_out_61, g5852, g3520, g1047, key_out_107;
wire I7099, I3848, I3699, I3398, I1969, I5307, g3974, key_out_111, I5536, g1417, I7543;
wire g5943, I7534, g4319, I3893, g2080, I2683, I5537, I3170, I3125, I5243, I1988;
wire I6194, g3207, I2526, g6929, g3215, I3446, I7208, g5783, I4545, I2004, I2527;
wire I5649, g6778, g1686, g4223, I1996, I3447, I4204, I3874, g2944, g1253, g2434;
wire I2299, g5866, g1687, I3935, g4017, I4528, I2244, I4151, I6392, key_out_58, I4010;
wire I2082, g5818, g3979, key_out_104, I6176, I4235, I2110, I7098, I3456, g5821, I3698;
wire g2995, I6473, I5659, g5636, I6177, I2899, I3457, I3989, I3971, I4160, I2089;
wire key_out_23, g4670, g4813, I3740, I8194, I5300, g3893, g6928, I7578, I7535, I1961;
wire g3544, g6394, I5648, I7246, g3756, I2062, I6195, I7216, g3536, I7564, g4300;
wire I4184, I2005, g5318, g5872, g5552, g4235, g6073, g4776, g4777, g4238, g6433;
wire g6496, g1422, g3931, g1560, g3905, g5094, g3973, g3528, g5541, g3621, g1449;
wire g3965, g3933, g6280, key_out_86, g2433, g1470, g6427, g6446, g6359, key_out_81, g1459;
wire g4584, g3926, g6279, key_out_82, g5265, g3927, g3903, g1418, g4578, g4261, g6358;
wire key_out_84, g4589, g1474, g3956, g4774, g5091, g4950, g5227, g4585, g6494, g5048;
wire g3664, g4000, g5418, g5093, g4779, g6492, g4240, g4596, g1603, g2908, g4581;
wire g5423, g4432, g6436, g4568, g6335, key_out_80, g5753, g6495, g6442, g6429, g6281;
wire key_out_85, g6449, g4590, g4877, g6445, g5561, g3929, g1473, g4967, g6430, g4993;
wire g6448, g3647, g3925, g5731, g3959, g1481, g3656, g4245, g3930, g5249, g3966;
wire g6400, key_out_79, g4266, g6451, g5324, g6443, g5088, g3958, g4241, g6432, g6357;
wire key_out_83, g3923, g6075, g3934, g6439, g4272, g1879, g5325, g6435, g4586, g3939;
wire g6438, g1518, g4239, g4591;
wire line1, line2, line3, line4, line5, line6, line7, line8, line9, line10, line11;
wire line12, line13, line14, line15, line16, line17, line18, line19, line20, line21, line22;
wire line23, line24, line25, line26, line27, line28, line29, line30, line31, line32, line33;
wire line34, line35, line36, line37, line38, line39, line40, line41, line42, line43, line44;
wire line45, line46, line47, line48, line49, line50, line51, line52, line53, line54, line55;
wire line56, line57, line58, line59, line60, line61, line62, line63, line64, line65, line66;
wire line67, line68, line69, line70, line71, line72, line73, line74, line75, line76, line77;
wire line78, line79, line80, line81, line82, line83, line84, line85, line86, line87, line88;
wire line89, line90, line91, line92, line93, line94, line95, line96, line97, line98, line99;
wire line100, line101, line102, line103, line104, line105, line106, line107, line108, line109, line110;
wire line111, line112, line113, line114, line115, line116, line117, line118, line119, line120, line121;
wire line122, line123, line124, line125, line126, line127, line128, line129, line130, line131, line132;
wire line133, line134, line135, line136, line137, line138, line139, line140, line141, line142, line143;
wire line144, line145, line146, line147, line148, line149, line150, line151, line152, line153, line154;
wire line155, line156, line157, line158, line159, line160, line161, line162, line163, line164, line165;
wire line166, line167, line168, line169, line170, line171, line172, line173, line174, line175, line176;
wire line177, line178, line179, line180, line181, line182, line183, line184, line185, line186, line187;
wire line188, line189, line190, line191, line192, line193, line194, line195, line196, line197, line198;
wire line199, line200, line201, line202, line203, line204, line205, line206, line207, line208, line209;
wire line210, line211;
DFFX1 gate1(.Q (g678), .QB (line1), .D(g4130), .CK(clk));
DFFX1 gate2(.Q (g332), .QB (line2), .D(g6823), .CK(clk));
DFFX1 gate3(.Q (g123), .QB (line3), .D(g6940), .CK(clk));
DFFX1 gate4(.Q (g207), .QB (line4), .D(g6102), .CK(clk));
DFFX1 gate5(.Q (g695), .QB (line5), .D(key_out_100), .CK(clk));
DFFX1 gate6(.Q (g461), .QB (line6), .D(g4841), .CK(clk));
DFFX1 gate7(.Q (g18), .QB (line7), .D(g6725), .CK(clk));
DFFX1 gate8(.Q (g292), .QB (line8), .D(g3232), .CK(clk));
DFFX1 gate9(.Q (g331), .QB (line9), .D(g4119), .CK(clk));
DFFX1 gate10(.Q (g689), .QB (line10), .D(g4141), .CK(clk));
DFFX1 gate11(.Q (g24), .QB (line11), .D(g6726), .CK(clk));
DFFX1 gate12(.Q (g465), .QB (line12), .D(g6507), .CK(clk));
DFFX1 gate13(.Q (g84), .QB (line13), .D(g6590), .CK(clk));
DFFX1 gate14(.Q (g291), .QB (line14), .D(g3231), .CK(clk));
DFFX1 gate15(.Q (g676), .QB (line15), .D(key_out_38), .CK(clk));
DFFX1 gate16(.Q (g622), .QB (line16), .D(g5147), .CK(clk));
DFFX1 gate17(.Q (g117), .QB (line17), .D(g4839), .CK(clk));
DFFX1 gate18(.Q (g278), .QB (line18), .D(g6105), .CK(clk));
DFFX1 gate19(.Q (g128), .QB (line19), .D(g5138), .CK(clk));
DFFX1 gate20(.Q (g598), .QB (line20), .D(g4122), .CK(clk));
DFFX1 gate21(.Q (g554), .QB (line21), .D(g6827), .CK(clk));
DFFX1 gate22(.Q (g496), .QB (line22), .D(g6745), .CK(clk));
DFFX1 gate23(.Q (g179), .QB (line23), .D(g6405), .CK(clk));
DFFX1 gate24(.Q (g48), .QB (line24), .D(g6729), .CK(clk));
DFFX1 gate25(.Q (g590), .QB (line25), .D(g6595), .CK(clk));
DFFX1 gate26(.Q (g551), .QB (line26), .D(g6826), .CK(clk));
DFFX1 gate27(.Q (g682), .QB (line27), .D(g4134), .CK(clk));
DFFX1 gate28(.Q (g11), .QB (line28), .D(g6599), .CK(clk));
DFFX1 gate29(.Q (g606), .QB (line29), .D(g4857), .CK(clk));
DFFX1 gate30(.Q (g188), .QB (line30), .D(g6406), .CK(clk));
DFFX1 gate31(.Q (g646), .QB (line31), .D(g5148), .CK(clk));
DFFX1 gate32(.Q (g327), .QB (line32), .D(g4117), .CK(clk));
DFFX1 gate33(.Q (g361), .QB (line33), .D(g6582), .CK(clk));
DFFX1 gate34(.Q (g289), .QB (line34), .D(g3229), .CK(clk));
DFFX1 gate35(.Q (g398), .QB (line35), .D(g5700), .CK(clk));
DFFX1 gate36(.Q (g684), .QB (line36), .D(g4136), .CK(clk));
DFFX1 gate37(.Q (g619), .QB (line37), .D(g4858), .CK(clk));
DFFX1 gate38(.Q (g208), .QB (line38), .D(g5876), .CK(clk));
DFFX1 gate39(.Q (g248), .QB (line39), .D(g3239), .CK(clk));
DFFX1 gate40(.Q (g390), .QB (line40), .D(g5698), .CK(clk));
DFFX1 gate41(.Q (g625), .QB (line41), .D(g5328), .CK(clk));
DFFX1 gate42(.Q (g681), .QB (line42), .D(g4133), .CK(clk));
DFFX1 gate43(.Q (g437), .QB (line43), .D(g4847), .CK(clk));
DFFX1 gate44(.Q (g276), .QB (line44), .D(g5877), .CK(clk));
DFFX1 gate45(.Q (g3), .QB (line45), .D(g6597), .CK(clk));
DFFX1 gate46(.Q (g323), .QB (line46), .D(g4120), .CK(clk));
DFFX1 gate47(.Q (g224), .QB (line47), .D(g3235), .CK(clk));
DFFX1 gate48(.Q (g685), .QB (line48), .D(g4137), .CK(clk));
DFFX1 gate49(.Q (g43), .QB (line49), .D(g6407), .CK(clk));
DFFX1 gate50(.Q (g157), .QB (line50), .D(g5470), .CK(clk));
DFFX1 gate51(.Q (g282), .QB (line51), .D(g6841), .CK(clk));
DFFX1 gate52(.Q (g697), .QB (line52), .D(key_out_92), .CK(clk));
DFFX1 gate53(.Q (g206), .QB (line53), .D(g6101), .CK(clk));
DFFX1 gate54(.Q (g449), .QB (line54), .D(g4844), .CK(clk));
DFFX1 gate55(.Q (g118), .QB (line55), .D(g4113), .CK(clk));
DFFX1 gate56(.Q (g528), .QB (line56), .D(g6504), .CK(clk));
DFFX1 gate57(.Q (g284), .QB (line57), .D(g3224), .CK(clk));
DFFX1 gate58(.Q (g426), .QB (line58), .D(g4855), .CK(clk));
DFFX1 gate59(.Q (g634), .QB (line59), .D(g4424), .CK(clk));
DFFX1 gate60(.Q (g669), .QB (line60), .D(g5582), .CK(clk));
DFFX1 gate61(.Q (g520), .QB (line61), .D(g6502), .CK(clk));
DFFX1 gate62(.Q (g281), .QB (line62), .D(g6107), .CK(clk));
DFFX1 gate63(.Q (g175), .QB (line63), .D(g5472), .CK(clk));
DFFX1 gate64(.Q (g15), .QB (line64), .D(g6602), .CK(clk));
DFFX1 gate65(.Q (g631), .QB (line65), .D(g5581), .CK(clk));
DFFX1 gate66(.Q (g69), .QB (line66), .D(g6587), .CK(clk));
DFFX1 gate67(.Q (g693), .QB (line67), .D(key_out_97), .CK(clk));
DFFX1 gate68(.Q (g337), .QB (line68), .D(g2585), .CK(clk));
DFFX1 gate69(.Q (g457), .QB (line69), .D(g4842), .CK(clk));
DFFX1 gate70(.Q (g486), .QB (line70), .D(g2586), .CK(clk));
DFFX1 gate71(.Q (g471), .QB (line71), .D(g1291), .CK(clk));
DFFX1 gate72(.Q (g328), .QB (line72), .D(g4118), .CK(clk));
DFFX1 gate73(.Q (g285), .QB (line73), .D(g3225), .CK(clk));
DFFX1 gate74(.Q (g418), .QB (line74), .D(g4853), .CK(clk));
DFFX1 gate75(.Q (g402), .QB (line75), .D(g4849), .CK(clk));
DFFX1 gate76(.Q (g297), .QB (line76), .D(g6512), .CK(clk));
DFFX1 gate77(.Q (g212), .QB (line77), .D(g3233), .CK(clk));
DFFX1 gate78(.Q (g410), .QB (line78), .D(g4851), .CK(clk));
DFFX1 gate79(.Q (g430), .QB (line79), .D(g4856), .CK(clk));
DFFX1 gate80(.Q (g33), .QB (line80), .D(g6854), .CK(clk));
DFFX1 gate81(.Q (g662), .QB (line81), .D(g1831), .CK(clk));
DFFX1 gate82(.Q (g453), .QB (line82), .D(g4843), .CK(clk));
DFFX1 gate83(.Q (g269), .QB (line83), .D(g6510), .CK(clk));
DFFX1 gate84(.Q (g574), .QB (line84), .D(g6591), .CK(clk));
DFFX1 gate85(.Q (g441), .QB (line85), .D(g4846), .CK(clk));
DFFX1 gate86(.Q (g664), .QB (line86), .D(g1288), .CK(clk));
DFFX1 gate87(.Q (g349), .QB (line87), .D(g5478), .CK(clk));
DFFX1 gate88(.Q (g211), .QB (line88), .D(g6840), .CK(clk));
DFFX1 gate89(.Q (g586), .QB (line89), .D(g6594), .CK(clk));
DFFX1 gate90(.Q (g571), .QB (line90), .D(g5580), .CK(clk));
DFFX1 gate91(.Q (g29), .QB (line91), .D(g6853), .CK(clk));
DFFX1 gate92(.Q (g326), .QB (line92), .D(g4840), .CK(clk));
DFFX1 gate93(.Q (g698), .QB (line93), .D(g4150), .CK(clk));
DFFX1 gate94(.Q (g654), .QB (line94), .D(g5490), .CK(clk));
DFFX1 gate95(.Q (g293), .QB (line95), .D(g6511), .CK(clk));
DFFX1 gate96(.Q (g690), .QB (line96), .D(key_out_93), .CK(clk));
DFFX1 gate97(.Q (g445), .QB (line97), .D(g4845), .CK(clk));
DFFX1 gate98(.Q (g374), .QB (line98), .D(g5694), .CK(clk));
DFFX1 gate99(.Q (g6), .QB (line99), .D(g6722), .CK(clk));
DFFX1 gate100(.Q (g687), .QB (line100), .D(g4139), .CK(clk));
DFFX1 gate101(.Q (g357), .QB (line101), .D(g5480), .CK(clk));
DFFX1 gate102(.Q (g386), .QB (line102), .D(g5697), .CK(clk));
DFFX1 gate103(.Q (g504), .QB (line103), .D(g6498), .CK(clk));
DFFX1 gate104(.Q (g665), .QB (line104), .D(g4126), .CK(clk));
DFFX1 gate105(.Q (g166), .QB (line105), .D(g5471), .CK(clk));
DFFX1 gate106(.Q (g541), .QB (line106), .D(g6505), .CK(clk));
DFFX1 gate107(.Q (g74), .QB (line107), .D(g6588), .CK(clk));
DFFX1 gate108(.Q (g338), .QB (line108), .D(g5475), .CK(clk));
DFFX1 gate109(.Q (g696), .QB (line109), .D(key_out_96), .CK(clk));
DFFX1 gate110(.Q (g516), .QB (line110), .D(g6501), .CK(clk));
DFFX1 gate111(.Q (g536), .QB (line111), .D(g6506), .CK(clk));
DFFX1 gate112(.Q (g683), .QB (line112), .D(g4135), .CK(clk));
DFFX1 gate113(.Q (g353), .QB (line113), .D(g5479), .CK(clk));
DFFX1 gate114(.Q (g545), .QB (line114), .D(g6824), .CK(clk));
DFFX1 gate115(.Q (g254), .QB (line115), .D(g3240), .CK(clk));
DFFX1 gate116(.Q (g341), .QB (line116), .D(g5476), .CK(clk));
DFFX1 gate117(.Q (g290), .QB (line117), .D(g3230), .CK(clk));
DFFX1 gate118(.Q (g2), .QB (line118), .D(g6721), .CK(clk));
DFFX1 gate119(.Q (g287), .QB (line119), .D(g3227), .CK(clk));
DFFX1 gate120(.Q (g336), .QB (line120), .D(g6925), .CK(clk));
DFFX1 gate121(.Q (g345), .QB (line121), .D(g5477), .CK(clk));
DFFX1 gate122(.Q (g628), .QB (line122), .D(g5489), .CK(clk));
DFFX1 gate123(.Q (g679), .QB (line123), .D(g4131), .CK(clk));
DFFX1 gate124(.Q (g28), .QB (line124), .D(g6727), .CK(clk));
DFFX1 gate125(.Q (g688), .QB (line125), .D(g4140), .CK(clk));
DFFX1 gate126(.Q (g283), .QB (line126), .D(g6842), .CK(clk));
DFFX1 gate127(.Q (g613), .QB (line127), .D(g4423), .CK(clk));
DFFX1 gate128(.Q (g10), .QB (line128), .D(g6723), .CK(clk));
DFFX1 gate129(.Q (g14), .QB (line129), .D(g6724), .CK(clk));
DFFX1 gate130(.Q (g680), .QB (line130), .D(g4132), .CK(clk));
DFFX1 gate131(.Q (g143), .QB (line131), .D(g6401), .CK(clk));
DFFX1 gate132(.Q (g672), .QB (line132), .D(g5491), .CK(clk));
DFFX1 gate133(.Q (g667), .QB (line133), .D(key_out_30), .CK(clk));
DFFX1 gate134(.Q (g366), .QB (line134), .D(g6278), .CK(clk));
DFFX1 gate135(.Q (g279), .QB (line135), .D(g6106), .CK(clk));
DFFX1 gate136(.Q (g492), .QB (line136), .D(g6744), .CK(clk));
DFFX1 gate137(.Q (g170), .QB (line137), .D(g6404), .CK(clk));
DFFX1 gate138(.Q (g686), .QB (line138), .D(g4138), .CK(clk));
DFFX1 gate139(.Q (g288), .QB (line139), .D(g3228), .CK(clk));
DFFX1 gate140(.Q (g638), .QB (line140), .D(key_out_103), .CK(clk));
DFFX1 gate141(.Q (g602), .QB (line141), .D(g4123), .CK(clk));
DFFX1 gate142(.Q (g642), .QB (line142), .D(g4658), .CK(clk));
DFFX1 gate143(.Q (g280), .QB (line143), .D(g5878), .CK(clk));
DFFX1 gate144(.Q (g663), .QB (line144), .D(g4125), .CK(clk));
DFFX1 gate145(.Q (g610), .QB (line145), .D(g4124), .CK(clk));
DFFX1 gate146(.Q (g148), .QB (line146), .D(g5874), .CK(clk));
DFFX1 gate147(.Q (g209), .QB (line147), .D(g6103), .CK(clk));
DFFX1 gate148(.Q (g675), .QB (line148), .D(key_out_39), .CK(clk));
DFFX1 gate149(.Q (g478), .QB (line149), .D(g1292), .CK(clk));
DFFX1 gate150(.Q (g122), .QB (line150), .D(g4115), .CK(clk));
DFFX1 gate151(.Q (g54), .QB (line151), .D(g6584), .CK(clk));
DFFX1 gate152(.Q (g594), .QB (line152), .D(g6596), .CK(clk));
DFFX1 gate153(.Q (g286), .QB (line153), .D(g3226), .CK(clk));
DFFX1 gate154(.Q (g489), .QB (line154), .D(g2587), .CK(clk));
DFFX1 gate155(.Q (g616), .QB (line155), .D(g4657), .CK(clk));
DFFX1 gate156(.Q (g79), .QB (line156), .D(g6589), .CK(clk));
DFFX1 gate157(.Q (g218), .QB (line157), .D(g3234), .CK(clk));
DFFX1 gate158(.Q (g242), .QB (line158), .D(g3238), .CK(clk));
DFFX1 gate159(.Q (g578), .QB (line159), .D(g6592), .CK(clk));
DFFX1 gate160(.Q (g184), .QB (line160), .D(g5473), .CK(clk));
DFFX1 gate161(.Q (g119), .QB (line161), .D(g4114), .CK(clk));
DFFX1 gate162(.Q (g668), .QB (line162), .D(g6800), .CK(clk));
DFFX1 gate163(.Q (g139), .QB (line163), .D(g5141), .CK(clk));
DFFX1 gate164(.Q (g422), .QB (line164), .D(g4854), .CK(clk));
DFFX1 gate165(.Q (g210), .QB (line165), .D(g6839), .CK(clk));
DFFX1 gate166(.Q (g394), .QB (line166), .D(g5699), .CK(clk));
DFFX1 gate167(.Q (g230), .QB (line167), .D(g3236), .CK(clk));
DFFX1 gate168(.Q (g25), .QB (line168), .D(g6601), .CK(clk));
DFFX1 gate169(.Q (g204), .QB (line169), .D(g5875), .CK(clk));
DFFX1 gate170(.Q (g658), .QB (line170), .D(g4425), .CK(clk));
DFFX1 gate171(.Q (g650), .QB (line171), .D(g5329), .CK(clk));
DFFX1 gate172(.Q (g378), .QB (line172), .D(g5695), .CK(clk));
DFFX1 gate173(.Q (g508), .QB (line173), .D(g6499), .CK(clk));
DFFX1 gate174(.Q (g548), .QB (line174), .D(g6825), .CK(clk));
DFFX1 gate175(.Q (g370), .QB (line175), .D(g5693), .CK(clk));
DFFX1 gate176(.Q (g406), .QB (line176), .D(g4850), .CK(clk));
DFFX1 gate177(.Q (g236), .QB (line177), .D(g3237), .CK(clk));
DFFX1 gate178(.Q (g500), .QB (line178), .D(g6497), .CK(clk));
DFFX1 gate179(.Q (g205), .QB (line179), .D(g6100), .CK(clk));
DFFX1 gate180(.Q (g197), .QB (line180), .D(g6509), .CK(clk));
DFFX1 gate181(.Q (g666), .QB (line181), .D(g4128), .CK(clk));
DFFX1 gate182(.Q (g114), .QB (line182), .D(g4116), .CK(clk));
DFFX1 gate183(.Q (g524), .QB (line183), .D(g6503), .CK(clk));
DFFX1 gate184(.Q (g260), .QB (line184), .D(g3241), .CK(clk));
DFFX1 gate185(.Q (g111), .QB (line185), .D(g6277), .CK(clk));
DFFX1 gate186(.Q (g131), .QB (line186), .D(g5139), .CK(clk));
DFFX1 gate187(.Q (g7), .QB (line187), .D(g6598), .CK(clk));
DFFX1 gate188(.Q (g19), .QB (line188), .D(g6600), .CK(clk));
DFFX1 gate189(.Q (g677), .QB (line189), .D(g4129), .CK(clk));
DFFX1 gate190(.Q (g582), .QB (line190), .D(g6593), .CK(clk));
DFFX1 gate191(.Q (g485), .QB (line191), .D(g6801), .CK(clk));
DFFX1 gate192(.Q (g699), .QB (line192), .D(key_out_102), .CK(clk));
DFFX1 gate193(.Q (g193), .QB (line193), .D(g5474), .CK(clk));
DFFX1 gate194(.Q (g135), .QB (line194), .D(g5140), .CK(clk));
DFFX1 gate195(.Q (g382), .QB (line195), .D(g5696), .CK(clk));
DFFX1 gate196(.Q (g414), .QB (line196), .D(g4852), .CK(clk));
DFFX1 gate197(.Q (g434), .QB (line197), .D(g4848), .CK(clk));
DFFX1 gate198(.Q (g266), .QB (line198), .D(g4659), .CK(clk));
DFFX1 gate199(.Q (g49), .QB (line199), .D(g6583), .CK(clk));
DFFX1 gate200(.Q (g152), .QB (line200), .D(g6402), .CK(clk));
DFFX1 gate201(.Q (g692), .QB (line201), .D(key_out_98), .CK(clk));
DFFX1 gate202(.Q (g277), .QB (line202), .D(g6104), .CK(clk));
DFFX1 gate203(.Q (g127), .QB (line203), .D(g6941), .CK(clk));
DFFX1 gate204(.Q (g161), .QB (line204), .D(g6403), .CK(clk));
DFFX1 gate205(.Q (g512), .QB (line205), .D(g6500), .CK(clk));
DFFX1 gate206(.Q (g532), .QB (line206), .D(g6508), .CK(clk));
DFFX1 gate207(.Q (g64), .QB (line207), .D(g6586), .CK(clk));
DFFX1 gate208(.Q (g694), .QB (line208), .D(key_out_99), .CK(clk));
DFFX1 gate209(.Q (g691), .QB (line209), .D(key_out_95), .CK(clk));
DFFX1 gate210(.Q (g1), .QB (line210), .D(g6720), .CK(clk));
DFFX1 gate211(.Q (g59), .QB (line211), .D(g6585), .CK(clk));
INVX1 gate212(.O (I8854), .I (g6696));
INVX1 gate213(.O (g1289), .I (I2272));
INVX1 gate214(.O (I9125), .I (g6855));
INVX1 gate215(.O (I6783), .I (g4822));
INVX1 gate216(.O (I4424), .I (g2097));
INVX1 gate217(.O (g6895), .I (I9152));
INVX1 gate218(.O (g1835), .I (I2919));
INVX1 gate219(.O (I3040), .I (g1770));
INVX1 gate220(.O (g6837), .I (g6822));
INVX1 gate221(.O (I7466), .I (g5624));
INVX1 gate222(.O (I4809), .I (g2974));
INVX1 gate223(.O (g3537), .I (I4757));
INVX1 gate224(.O (g5457), .I (g5304));
INVX1 gate225(.O (g6062), .I (g5824));
INVX1 gate226(.O (g4040), .I (I5343));
INVX1 gate227(.O (I6001), .I (g4162));
INVX1 gate228(.O (g5549), .I (g5331));
INVX1 gate229(.O (I4477), .I (g3063));
INVX1 gate230(.O (g3612), .I (I4809));
INVX1 gate231(.O (I7055), .I (g5318));
INVX1 gate232(.O (g2892), .I (g1982));
INVX1 gate233(.O (I5264), .I (g3638));
INVX1 gate234(.O (I2225), .I (g696));
INVX1 gate235(.O (g4123), .I (I5451));
INVX1 gate236(.O (g4323), .I (g4086));
INVX1 gate237(.O (g908), .I (I1932));
INVX1 gate238(.O (I5933), .I (g4346));
INVX1 gate239(.O (I8252), .I (g6294));
INVX1 gate240(.O (I2473), .I (g971));
INVX1 gate241(.O (I7333), .I (g5386));
INVX1 gate242(.O (I8812), .I (g6688));
INVX1 gate243(.O (g1674), .I (g985));
INVX1 gate244(.O (I3528), .I (g1422));
INVX1 gate245(.O (I8958), .I (g6774));
INVX1 gate246(.O (I5050), .I (g3246));
INVX1 gate247(.O (g3234), .I (I4501));
INVX1 gate248(.O (I2324), .I (key_out_128));
INVX1 gate249(.O (g2945), .I (I4133));
INVX1 gate250(.O (g5121), .I (I6775));
INVX1 gate251(.O (g1997), .I (g1398));
INVX1 gate252(.O (g3128), .I (I4375));
INVX1 gate253(.O (I8005), .I (g6110));
INVX1 gate254(.O (g1541), .I (g1094));
INVX1 gate255(.O (g5670), .I (g5527));
INVX1 gate256(.O (g2738), .I (g2327));
INVX1 gate257(.O (g6842), .I (I9047));
INVX1 gate258(.O (g4528), .I (I6096));
INVX1 gate259(.O (g2244), .I (I3379));
INVX1 gate260(.O (g6192), .I (g5946));
INVX1 gate261(.O (g2709), .I (I3864));
INVX1 gate262(.O (g1332), .I (I2349));
INVX1 gate263(.O (g4530), .I (I6102));
INVX1 gate264(.O (g1680), .I (g1011));
INVX1 gate265(.O (g2078), .I (g1345));
INVX1 gate266(.O (g1209), .I (I2215));
INVX1 gate267(.O (I3010), .I (g1504));
INVX1 gate268(.O (g5813), .I (I7612));
INVX1 gate269(.O (I7509), .I (g5587));
INVX1 gate270(.O (I5379), .I (g3940));
INVX1 gate271(.O (g3800), .I (g3388));
INVX1 gate272(.O (g2907), .I (g1914));
INVX1 gate273(.O (g6854), .I (I9085));
INVX1 gate274(.O (g2035), .I (I3144));
INVX1 gate275(.O (g2959), .I (g1861));
INVX1 gate276(.O (g6941), .I (I9236));
INVX1 gate277(.O (g4010), .I (g3601));
INVX1 gate278(.O (I2287), .I (g927));
INVX1 gate279(.O (I4273), .I (g2197));
INVX1 gate280(.O (I8270), .I (g6300));
INVX1 gate281(.O (g5740), .I (I7501));
INVX1 gate282(.O (I5777), .I (g3807));
INVX1 gate283(.O (g2876), .I (g1943));
INVX1 gate284(.O (g873), .I (g306));
INVX1 gate285(.O (g4839), .I (I6525));
INVX1 gate286(.O (I5882), .I (g3871));
INVX1 gate287(.O (g2656), .I (I3800));
INVX1 gate288(.O (I8473), .I (g6485));
INVX1 gate289(.O (I2199), .I (g33));
INVX1 gate290(.O (g900), .I (I1927));
INVX1 gate291(.O (g6708), .I (I8834));
INVX1 gate292(.O (I2399), .I (g729));
INVX1 gate293(.O (I3278), .I (g1695));
INVX1 gate294(.O (g6520), .I (I8476));
INVX1 gate295(.O (g940), .I (g64));
INVX1 gate296(.O (I6677), .I (g4757));
INVX1 gate297(.O (g3902), .I (g3575));
INVX1 gate298(.O (g5687), .I (g5567));
INVX1 gate299(.O (g2915), .I (g1931));
INVX1 gate300(.O (g847), .I (g590));
INVX1 gate301(.O (I3235), .I (g1807));
INVX1 gate302(.O (I3343), .I (g1623));
INVX1 gate303(.O (g6431), .I (I8295));
INVX1 gate304(.O (g709), .I (g114));
INVX1 gate305(.O (g6812), .I (I8984));
INVX1 gate306(.O (I6576), .I (g4700));
INVX1 gate307(.O (g749), .I (I1847));
INVX1 gate308(.O (g3090), .I (I4331));
INVX1 gate309(.O (I9107), .I (g6855));
INVX1 gate310(.O (g2214), .I (I3349));
INVX1 gate311(.O (g4618), .I (g4246));
INVX1 gate312(.O (g6376), .I (g6267));
INVX1 gate313(.O (g4143), .I (I5511));
INVX1 gate314(.O (I6349), .I (g4569));
INVX1 gate315(.O (g4343), .I (g4011));
INVX1 gate316(.O (I5674), .I (g4003));
INVX1 gate317(.O (I8177), .I (g6173));
INVX1 gate318(.O (g2110), .I (g1381));
INVX1 gate319(.O (I3134), .I (g1336));
INVX1 gate320(.O (g6405), .I (I8229));
INVX1 gate321(.O (I3334), .I (g1330));
INVX1 gate322(.O (I7197), .I (g5431));
INVX1 gate323(.O (g4566), .I (g4198));
INVX1 gate324(.O (I7397), .I (g5561));
INVX1 gate325(.O (I4534), .I (g2858));
INVX1 gate326(.O (g1714), .I (g1110));
INVX1 gate327(.O (I4961), .I (g3597));
INVX1 gate328(.O (g2663), .I (g2308));
INVX1 gate329(.O (g3456), .I (g2640));
INVX1 gate330(.O (g5141), .I (I6801));
INVX1 gate331(.O (g922), .I (I1947));
INVX1 gate332(.O (g4693), .I (I6283));
INVX1 gate333(.O (g4134), .I (I5484));
INVX1 gate334(.O (g5570), .I (g5392));
INVX1 gate335(.O (g5860), .I (g5634));
INVX1 gate336(.O (g4334), .I (g3733));
INVX1 gate337(.O (I3804), .I (g2575));
INVX1 gate338(.O (I2207), .I (g7));
INVX1 gate339(.O (I5153), .I (g3330));
INVX1 gate340(.O (g3355), .I (g3100));
INVX1 gate341(.O (g5645), .I (g5537));
INVX1 gate342(.O (g6733), .I (I8891));
INVX1 gate343(.O (g5691), .I (g5568));
INVX1 gate344(.O (g4804), .I (g4473));
INVX1 gate345(.O (I9047), .I (g6838));
INVX1 gate346(.O (I4414), .I (g2090));
INVX1 gate347(.O (g6610), .I (I8696));
INVX1 gate348(.O (g2877), .I (g2434));
INVX1 gate349(.O (I4903), .I (g3223));
INVX1 gate350(.O (g6796), .I (I8958));
INVX1 gate351(.O (g3063), .I (I4288));
INVX1 gate352(.O (I3313), .I (g1337));
INVX1 gate353(.O (g5879), .I (g5770));
INVX1 gate354(.O (g3463), .I (g2682));
INVX1 gate355(.O (I4513), .I (g2765));
INVX1 gate356(.O (g1623), .I (I2578));
INVX1 gate357(.O (g5358), .I (I7012));
INVX1 gate358(.O (I3202), .I (g1812));
INVX1 gate359(.O (I2215), .I (g695));
INVX1 gate360(.O (g4113), .I (I5421));
INVX1 gate361(.O (g1076), .I (I2115));
INVX1 gate362(.O (g6069), .I (g5791));
INVX1 gate363(.O (I7817), .I (g5924));
INVX1 gate364(.O (g6540), .I (g6474));
INVX1 gate365(.O (I6352), .I (g4564));
INVX1 gate366(.O (I1865), .I (g279));
INVX1 gate367(.O (g4202), .I (I5622));
INVX1 gate368(.O (I6867), .I (g5082));
INVX1 gate369(.O (I5511), .I (g3876));
INVX1 gate370(.O (g5587), .I (I7349));
INVX1 gate371(.O (I8144), .I (g6182));
INVX1 gate372(.O (g1175), .I (g42));
INVX1 gate373(.O (g1375), .I (I2411));
INVX1 gate374(.O (g3118), .I (I4366));
INVX1 gate375(.O (g3318), .I (I4593));
INVX1 gate376(.O (g2464), .I (I3596));
INVX1 gate377(.O (g3872), .I (g3312));
INVX1 gate378(.O (g4494), .I (I6004));
INVX1 gate379(.O (I2870), .I (key_out_126));
INVX1 gate380(.O (g4518), .I (I6066));
INVX1 gate381(.O (I4288), .I (g2215));
INVX1 gate382(.O (g5615), .I (I7372));
INVX1 gate383(.O (g4567), .I (I6139));
INVX1 gate384(.O (I4382), .I (g2265));
INVX1 gate385(.O (I3776), .I (g2044));
INVX1 gate386(.O (g3057), .I (I4282));
INVX1 gate387(.O (I5600), .I (g3821));
INVX1 gate388(.O (I3593), .I (g1295));
INVX1 gate389(.O (I2825), .I (key_out_123));
INVX1 gate390(.O (g1285), .I (g852));
INVX1 gate391(.O (g3457), .I (g2653));
INVX1 gate392(.O (g5174), .I (g5099));
INVX1 gate393(.O (I6386), .I (g4462));
INVX1 gate394(.O (I3965), .I (g2268));
INVX1 gate395(.O (I8488), .I (g6426));
INVX1 gate396(.O (g6849), .I (I9074));
INVX1 gate397(.O (I6599), .I (g4823));
INVX1 gate398(.O (I2408), .I (g719));
INVX1 gate399(.O (g3834), .I (I5027));
INVX1 gate400(.O (g2295), .I (g1578));
INVX1 gate401(.O (g1384), .I (I2420));
INVX1 gate402(.O (g1339), .I (I2370));
INVX1 gate403(.O (g5545), .I (g5331));
INVX1 gate404(.O (I6170), .I (g4343));
INVX1 gate405(.O (I9128), .I (g6864));
INVX1 gate406(.O (g6898), .I (I9161));
INVX1 gate407(.O (g1838), .I (g1595));
INVX1 gate408(.O (g6900), .I (I9167));
INVX1 gate409(.O (g2194), .I (I3331));
INVX1 gate410(.O (g6797), .I (I8961));
INVX1 gate411(.O (g2394), .I (I3537));
INVX1 gate412(.O (I3050), .I (g1439));
INVX1 gate413(.O (I3641), .I (g1491));
INVX1 gate414(.O (I2943), .I (g1715));
INVX1 gate415(.O (I5736), .I (g4022));
INVX1 gate416(.O (g6510), .I (I8450));
INVX1 gate417(.O (I6280), .I (g4430));
INVX1 gate418(.O (g4933), .I (I6625));
INVX1 gate419(.O (g5420), .I (I7086));
INVX1 gate420(.O (g4521), .I (I6075));
INVX1 gate421(.O (g1672), .I (g1094));
INVX1 gate422(.O (I7058), .I (g5281));
INVX1 gate423(.O (I2887), .I (key_out_122));
INVX1 gate424(.O (I2122), .I (g689));
INVX1 gate425(.O (g1477), .I (g952));
INVX1 gate426(.O (g3232), .I (I4495));
INVX1 gate427(.O (I2228), .I (g15));
INVX1 gate428(.O (g5794), .I (I7593));
INVX1 gate429(.O (g1643), .I (I2608));
INVX1 gate430(.O (I4495), .I (g3022));
INVX1 gate431(.O (I4437), .I (g2108));
INVX1 gate432(.O (g2705), .I (I3858));
INVX1 gate433(.O (g3813), .I (g3258));
INVX1 gate434(.O (I8650), .I (g6529));
INVX1 gate435(.O (I3379), .I (g1647));
INVX1 gate436(.O (g2242), .I (I3373));
INVX1 gate437(.O (g1205), .I (g45));
INVX1 gate438(.O (I2033), .I (g678));
INVX1 gate439(.O (I5871), .I (g3744));
INVX1 gate440(.O (g774), .I (I1859));
INVX1 gate441(.O (g6819), .I (I8994));
INVX1 gate442(.O (g6694), .I (I8800));
INVX1 gate443(.O (g4379), .I (I5848));
INVX1 gate444(.O (g5905), .I (g5852));
INVX1 gate445(.O (g3519), .I (g2740));
INVX1 gate446(.O (I7856), .I (g5994));
INVX1 gate447(.O (g921), .I (g111));
INVX1 gate448(.O (g1551), .I (g1011));
INVX1 gate449(.O (g1742), .I (I2756));
INVX1 gate450(.O (I4752), .I (g2859));
INVX1 gate451(.O (g6488), .I (g6367));
INVX1 gate452(.O (g2254), .I (I3391));
INVX1 gate453(.O (I8594), .I (g6446));
INVX1 gate454(.O (g2814), .I (I4023));
INVX1 gate455(.O (g4289), .I (I5746));
INVX1 gate456(.O (g4658), .I (I6247));
INVX1 gate457(.O (I6756), .I (g4775));
INVX1 gate458(.O (g6701), .I (I8821));
INVX1 gate459(.O (I8972), .I (g6795));
INVX1 gate460(.O (I3271), .I (g1748));
INVX1 gate461(.O (I2845), .I (key_out_127));
INVX1 gate462(.O (g5300), .I (I6952));
INVX1 gate463(.O (g2350), .I (I3502));
INVX1 gate464(.O (I8806), .I (g6686));
INVX1 gate465(.O (I3611), .I (g1771));
INVX1 gate466(.O (I2137), .I (g1));
INVX1 gate467(.O (I8943), .I (g6774));
INVX1 gate468(.O (I2337), .I (key_out_128));
INVX1 gate469(.O (I2913), .I (g1792));
INVX1 gate470(.O (g1754), .I (I2773));
INVX1 gate471(.O (g6886), .I (I9125));
INVX1 gate472(.O (g2409), .I (g1815));
INVX1 gate473(.O (g894), .I (I1917));
INVX1 gate474(.O (g1273), .I (key_out_31));
INVX1 gate475(.O (I5424), .I (g3725));
INVX1 gate476(.O (I6403), .I (g4492));
INVX1 gate477(.O (g6314), .I (I8044));
INVX1 gate478(.O (g4799), .I (g4485));
INVX1 gate479(.O (I9155), .I (g6882));
INVX1 gate480(.O (g2836), .I (g2509));
INVX1 gate481(.O (g2212), .I (I3343));
INVX1 gate482(.O (I6763), .I (g4780));
INVX1 gate483(.O (g3860), .I (I5081));
INVX1 gate484(.O (g2967), .I (I4166));
INVX1 gate485(.O (g6825), .I (I9008));
INVX1 gate486(.O (g5440), .I (g5266));
INVX1 gate487(.O (g3710), .I (g3029));
INVX1 gate488(.O (I5523), .I (g3840));
INVX1 gate489(.O (g843), .I (g574));
INVX1 gate490(.O (g1543), .I (g1006));
INVX1 gate491(.O (g4132), .I (I5478));
INVX1 gate492(.O (g6408), .I (g6283));
INVX1 gate493(.O (g4153), .I (I5545));
INVX1 gate494(.O (I6359), .I (g4566));
INVX1 gate495(.O (g6136), .I (I7856));
INVX1 gate496(.O (g2822), .I (I4031));
INVX1 gate497(.O (I8891), .I (g6706));
INVX1 gate498(.O (I8913), .I (g6743));
INVX1 gate499(.O (I2692), .I (g1037));
INVX1 gate500(.O (g6594), .I (I8650));
INVX1 gate501(.O (g946), .I (g361));
INVX1 gate502(.O (g1729), .I (I2731));
INVX1 gate503(.O (I5551), .I (g4059));
INVX1 gate504(.O (g4802), .I (I6470));
INVX1 gate505(.O (g3962), .I (I5214));
INVX1 gate506(.O (I2154), .I (g14));
INVX1 gate507(.O (I4189), .I (g2159));
INVX1 gate508(.O (I5499), .I (g3847));
INVX1 gate509(.O (g5151), .I (I6819));
INVX1 gate510(.O (g3158), .I (I4398));
INVX1 gate511(.O (g6806), .I (I8978));
INVX1 gate512(.O (I4706), .I (g2877));
INVX1 gate513(.O (g5875), .I (I7637));
INVX1 gate514(.O (g5530), .I (I7270));
INVX1 gate515(.O (I9167), .I (g6878));
INVX1 gate516(.O (I5926), .I (g4153));
INVX1 gate517(.O (g2921), .I (g1950));
INVX1 gate518(.O (g6065), .I (g5784));
INVX1 gate519(.O (I6315), .I (g4446));
INVX1 gate520(.O (I4371), .I (g2555));
INVX1 gate521(.O (g6887), .I (I9128));
INVX1 gate522(.O (I4429), .I (g2102));
INVX1 gate523(.O (g6122), .I (I7838));
INVX1 gate524(.O (g6465), .I (I8329));
INVX1 gate525(.O (g6322), .I (I8056));
INVX1 gate526(.O (g1660), .I (g985));
INVX1 gate527(.O (g1946), .I (I3053));
INVX1 gate528(.O (g6230), .I (g6040));
INVX1 gate529(.O (g5010), .I (I6646));
INVX1 gate530(.O (g4511), .I (I6045));
INVX1 gate531(.O (I6874), .I (g4861));
INVX1 gate532(.O (g2895), .I (g1894));
INVX1 gate533(.O (g6033), .I (g5824));
INVX1 gate534(.O (g2837), .I (g2512));
INVX1 gate535(.O (I2979), .I (g1263));
INVX1 gate536(.O (I3864), .I (g2044));
INVX1 gate537(.O (g5884), .I (g5864));
INVX1 gate538(.O (I8342), .I (g6314));
INVX1 gate539(.O (I2218), .I (g11));
INVX1 gate540(.O (g1513), .I (g878));
INVX1 gate541(.O (I2312), .I (g897));
INVX1 gate542(.O (I3714), .I (g1852));
INVX1 gate543(.O (I4297), .I (g2555));
INVX1 gate544(.O (I8255), .I (g6292));
INVX1 gate545(.O (I8815), .I (g6689));
INVX1 gate546(.O (g4492), .I (I5998));
INVX1 gate547(.O (I1868), .I (g280));
INVX1 gate548(.O (I7608), .I (g5605));
INVX1 gate549(.O (I5862), .I (g3863));
INVX1 gate550(.O (g1679), .I (g985));
INVX1 gate551(.O (g1378), .I (I2414));
INVX1 gate552(.O (g4714), .I (I6324));
INVX1 gate553(.O (I2293), .I (g971));
INVX1 gate554(.O (g5278), .I (I6937));
INVX1 gate555(.O (g3284), .I (g3019));
INVX1 gate556(.O (I4684), .I (g2687));
INVX1 gate557(.O (I8497), .I (g6481));
INVX1 gate558(.O (g3239), .I (I4516));
INVX1 gate559(.O (I6537), .I (g4711));
INVX1 gate560(.O (g3545), .I (g3085));
INVX1 gate561(.O (g2788), .I (I3983));
INVX1 gate562(.O (g6137), .I (I7859));
INVX1 gate563(.O (g5667), .I (g5524));
INVX1 gate564(.O (g6891), .I (I9140));
INVX1 gate565(.O (g1831), .I (I2907));
INVX1 gate566(.O (g1335), .I (I2358));
INVX1 gate567(.O (g3380), .I (g2831));
INVX1 gate568(.O (I4791), .I (g2814));
INVX1 gate569(.O (g6337), .I (I8089));
INVX1 gate570(.O (I4309), .I (g2525));
INVX1 gate571(.O (I2828), .I (key_out_127));
INVX1 gate572(.O (g3832), .I (I5023));
INVX1 gate573(.O (g1288), .I (I2269));
INVX1 gate574(.O (g5566), .I (I7318));
INVX1 gate575(.O (g3853), .I (I5068));
INVX1 gate576(.O (I3736), .I (g2460));
INVX1 gate577(.O (I6612), .I (g4660));
INVX1 gate578(.O (I7161), .I (g5465));
INVX1 gate579(.O (I7361), .I (g5566));
INVX1 gate580(.O (g2842), .I (I4050));
INVX1 gate581(.O (g1805), .I (I2854));
INVX1 gate582(.O (I6417), .I (g4617));
INVX1 gate583(.O (I3623), .I (g1491));
INVX1 gate584(.O (g4262), .I (I5713));
INVX1 gate585(.O (I7051), .I (g5219));
INVX1 gate586(.O (I2221), .I (g43));
INVX1 gate587(.O (g3559), .I (g2603));
INVX1 gate588(.O (g4736), .I (I6366));
INVX1 gate589(.O (g2485), .I (I3614));
INVX1 gate590(.O (I7451), .I (g5597));
INVX1 gate591(.O (I2703), .I (g1189));
INVX1 gate592(.O (I8267), .I (g6297));
INVX1 gate593(.O (g4623), .I (g4262));
INVX1 gate594(.O (g1947), .I (I3056));
INVX1 gate595(.O (I5885), .I (g3746));
INVX1 gate596(.O (I7999), .I (g6137));
INVX1 gate597(.O (g878), .I (g639));
INVX1 gate598(.O (I7146), .I (g5231));
INVX1 gate599(.O (I6330), .I (g4560));
INVX1 gate600(.O (I7346), .I (g5531));
INVX1 gate601(.O (I3871), .I (g2145));
INVX1 gate602(.O (I8329), .I (g6305));
INVX1 gate603(.O (g4375), .I (I5840));
INVX1 gate604(.O (g4871), .I (I6599));
INVX1 gate605(.O (I8761), .I (g6563));
INVX1 gate606(.O (g3204), .I (I4441));
INVX1 gate607(.O (g4722), .I (I6346));
INVX1 gate608(.O (g710), .I (g128));
INVX1 gate609(.O (I4498), .I (g2686));
INVX1 gate610(.O (g829), .I (g323));
INVX1 gate611(.O (g5113), .I (I6753));
INVX1 gate612(.O (g1632), .I (g760));
INVX1 gate613(.O (g1037), .I (I2067));
INVX1 gate614(.O (g3100), .I (I4347));
INVX1 gate615(.O (I8828), .I (g6661));
INVX1 gate616(.O (g6726), .I (I8872));
INVX1 gate617(.O (g6497), .I (I8411));
INVX1 gate618(.O (g1653), .I (I2630));
INVX1 gate619(.O (g2640), .I (I3782));
INVX1 gate620(.O (I8727), .I (g6536));
INVX1 gate621(.O (g2031), .I (I3140));
INVX1 gate622(.O (I5436), .I (g3729));
INVX1 gate623(.O (g2252), .I (I3385));
INVX1 gate624(.O (g5908), .I (g5753));
INVX1 gate625(.O (g2958), .I (g1861));
INVX1 gate626(.O (I7472), .I (g5626));
INVX1 gate627(.O (g2176), .I (I3319));
INVX1 gate628(.O (I2716), .I (g1115));
INVX1 gate629(.O (I5831), .I (g3842));
INVX1 gate630(.O (I2349), .I (g1160));
INVX1 gate631(.O (g4139), .I (I5499));
INVX1 gate632(.O (I5182), .I (key_out_5));
INVX1 gate633(.O (g5518), .I (I7258));
INVX1 gate634(.O (g5567), .I (g5418));
INVX1 gate635(.O (I5382), .I (g3952));
INVX1 gate636(.O (g2405), .I (I3543));
INVX1 gate637(.O (I2848), .I (key_out_127));
INVX1 gate638(.O (g1917), .I (I3016));
INVX1 gate639(.O (g2829), .I (g2491));
INVX1 gate640(.O (g2765), .I (I3946));
INVX1 gate641(.O (I7116), .I (g5299));
INVX1 gate642(.O (I4019), .I (g1841));
INVX1 gate643(.O (g4424), .I (I5923));
INVX1 gate644(.O (I6090), .I (g4393));
INVX1 gate645(.O (I4362), .I (g2555));
INVX1 gate646(.O (I3672), .I (g1656));
INVX1 gate647(.O (g3040), .I (I4255));
INVX1 gate648(.O (I3077), .I (g1439));
INVX1 gate649(.O (g4809), .I (I6485));
INVX1 gate650(.O (g5593), .I (I7355));
INVX1 gate651(.O (g3440), .I (I4678));
INVX1 gate652(.O (g3969), .I (I5233));
INVX1 gate653(.O (g6312), .I (I8040));
INVX1 gate654(.O (I6366), .I (g4569));
INVX1 gate655(.O (I4452), .I (g2117));
INVX1 gate656(.O (g2974), .I (I4173));
INVX1 gate657(.O (g6401), .I (I8217));
INVX1 gate658(.O (g895), .I (g139));
INVX1 gate659(.O (I6456), .I (g4633));
INVX1 gate660(.O (g4523), .I (I6081));
INVX1 gate661(.O (g1233), .I (I2231));
INVX1 gate662(.O (I6649), .I (g4693));
INVX1 gate663(.O (g4643), .I (g4293));
INVX1 gate664(.O (g5264), .I (g4943));
INVX1 gate665(.O (I9158), .I (g6887));
INVX1 gate666(.O (g1054), .I (g485));
INVX1 gate667(.O (g5160), .I (g5099));
INVX1 gate668(.O (g2796), .I (I3999));
INVX1 gate669(.O (I6355), .I (g4569));
INVX1 gate670(.O (g2473), .I (I3605));
INVX1 gate671(.O (I3099), .I (g1519));
INVX1 gate672(.O (I8576), .I (g6436));
INVX1 gate673(.O (g1770), .I (I2805));
INVX1 gate674(.O (I8866), .I (g6701));
INVX1 gate675(.O (I3304), .I (g1740));
INVX1 gate676(.O (I4486), .I (g3093));
INVX1 gate677(.O (g5521), .I (I7261));
INVX1 gate678(.O (I3499), .I (g1450));
INVX1 gate679(.O (I8716), .I (g6518));
INVX1 gate680(.O (g1725), .I (g1113));
INVX1 gate681(.O (I7596), .I (g5605));
INVX1 gate682(.O (g6727), .I (I8875));
INVX1 gate683(.O (g3875), .I (I5106));
INVX1 gate684(.O (g2324), .I (I3478));
INVX1 gate685(.O (I4504), .I (g2726));
INVX1 gate686(.O (I2119), .I (g688));
INVX1 gate687(.O (g5450), .I (g5292));
INVX1 gate688(.O (I5037), .I (g3705));
INVX1 gate689(.O (g5996), .I (g5824));
INVX1 gate690(.O (g4104), .I (I5394));
INVX1 gate691(.O (g6592), .I (I8644));
INVX1 gate692(.O (g4099), .I (I5379));
INVX1 gate693(.O (g4499), .I (I6015));
INVX1 gate694(.O (I2352), .I (key_out_126));
INVX1 gate695(.O (I6063), .I (g4381));
INVX1 gate696(.O (g6746), .I (I8916));
INVX1 gate697(.O (I2867), .I (key_out_123));
INVX1 gate698(.O (I8699), .I (g6573));
INVX1 gate699(.O (g2177), .I (I3322));
INVX1 gate700(.O (g5179), .I (g5099));
INVX1 gate701(.O (g5379), .I (I7035));
INVX1 gate702(.O (I2893), .I (key_out_120));
INVX1 gate703(.O (g5878), .I (I7646));
INVX1 gate704(.O (I3044), .I (g1257));
INVX1 gate705(.O (g1189), .I (I2196));
INVX1 gate706(.O (g3839), .I (I5040));
INVX1 gate707(.O (g6932), .I (I9217));
INVX1 gate708(.O (g4273), .I (I5728));
INVX1 gate709(.O (g5658), .I (g5512));
INVX1 gate710(.O (g6624), .I (I8730));
INVX1 gate711(.O (I6118), .I (g4406));
INVX1 gate712(.O (I6318), .I (g4447));
INVX1 gate713(.O (I3983), .I (g2276));
INVX1 gate714(.O (g2849), .I (g2577));
INVX1 gate715(.O (I3572), .I (g1295));
INVX1 gate716(.O (g1787), .I (I2835));
INVX1 gate717(.O (I5442), .I (g3731));
INVX1 gate718(.O (I4678), .I (g2670));
INVX1 gate719(.O (I6057), .I (g4379));
INVX1 gate720(.O (I8524), .I (g6496));
INVX1 gate721(.O (I4331), .I (g2555));
INVX1 gate722(.O (I8644), .I (g6526));
INVX1 gate723(.O (I3543), .I (g1461));
INVX1 gate724(.O (I6989), .I (g5307));
INVX1 gate725(.O (I2614), .I (key_out_122));
INVX1 gate726(.O (g1675), .I (g1101));
INVX1 gate727(.O (I2370), .I (key_out_122));
INVX1 gate728(.O (I2125), .I (g698));
INVX1 gate729(.O (g3235), .I (I4504));
INVX1 gate730(.O (g3343), .I (g3090));
INVX1 gate731(.O (I5233), .I (key_out_4));
INVX1 gate732(.O (I2821), .I (g1221));
INVX1 gate733(.O (g4712), .I (I6318));
INVX1 gate734(.O (g985), .I (g638));
INVX1 gate735(.O (g6576), .I (g6487));
INVX1 gate736(.O (I6549), .I (g4699));
INVX1 gate737(.O (I8258), .I (g6293));
INVX1 gate738(.O (I8818), .I (g6690));
INVX1 gate739(.O (I3534), .I (g1295));
INVX1 gate740(.O (g2245), .I (I3382));
INVX1 gate741(.O (I3729), .I (g2436));
INVX1 gate742(.O (I3961), .I (g1835));
INVX1 gate743(.O (I5454), .I (g3874));
INVX1 gate744(.O (g2291), .I (I3434));
INVX1 gate745(.O (g5997), .I (g5854));
INVX1 gate746(.O (g4534), .I (I6114));
INVX1 gate747(.O (I3927), .I (g2245));
INVX1 gate748(.O (I5532), .I (g3861));
INVX1 gate749(.O (g1684), .I (I2668));
INVX1 gate750(.O (g6699), .I (I8815));
INVX1 gate751(.O (g1639), .I (g815));
INVX1 gate752(.O (g1338), .I (I2367));
INVX1 gate753(.O (g1963), .I (I3074));
INVX1 gate754(.O (I8186), .I (g6179));
INVX1 gate755(.O (I6321), .I (g4559));
INVX1 gate756(.O (I4226), .I (g2525));
INVX1 gate757(.O (g1109), .I (I2137));
INVX1 gate758(.O (g1791), .I (I2845));
INVX1 gate759(.O (I8975), .I (g6791));
INVX1 gate760(.O (I3946), .I (g2256));
INVX1 gate761(.O (g889), .I (g310));
INVX1 gate762(.O (I2306), .I (g896));
INVX1 gate763(.O (g3792), .I (g3388));
INVX1 gate764(.O (I6625), .I (g4745));
INVX1 gate765(.O (g2819), .I (g2467));
INVX1 gate766(.O (g4014), .I (I5316));
INVX1 gate767(.O (I8426), .I (g6424));
INVX1 gate768(.O (I5412), .I (g4034));
INVX1 gate769(.O (g4660), .I (I6253));
INVX1 gate770(.O (I6253), .I (g4608));
INVX1 gate771(.O (g2088), .I (I3202));
INVX1 gate772(.O (g2923), .I (g1969));
INVX1 gate773(.O (I4173), .I (g2408));
INVX1 gate774(.O (I8614), .I (g6537));
INVX1 gate775(.O (I3513), .I (g1450));
INVX1 gate776(.O (g2488), .I (I3617));
INVX1 gate777(.O (g1759), .I (I2782));
INVX1 gate778(.O (I2756), .I (g1175));
INVX1 gate779(.O (g2701), .I (I3855));
INVX1 gate780(.O (I7190), .I (g5432));
INVX1 gate781(.O (I8821), .I (g6691));
INVX1 gate782(.O (g6524), .I (I8488));
INVX1 gate783(.O (I6740), .I (g4781));
INVX1 gate784(.O (g4513), .I (I6051));
INVX1 gate785(.O (I8984), .I (g6794));
INVX1 gate786(.O (I7501), .I (g5596));
INVX1 gate787(.O (g1957), .I (I3068));
INVX1 gate788(.O (g2215), .I (I3352));
INVX1 gate789(.O (g6119), .I (I7829));
INVX1 gate790(.O (I2904), .I (g1256));
INVX1 gate791(.O (g6319), .I (I8051));
INVX1 gate792(.O (g1049), .I (g266));
INVX1 gate793(.O (g5901), .I (g5753));
INVX1 gate794(.O (g2886), .I (g1966));
INVX1 gate795(.O (I6552), .I (g4702));
INVX1 gate796(.O (I4059), .I (g1878));
INVX1 gate797(.O (g4036), .I (I5337));
INVX1 gate798(.O (g3094), .I (I4337));
INVX1 gate799(.O (I4459), .I (g2134));
INVX1 gate800(.O (I8544), .I (g6453));
INVX1 gate801(.O (g4679), .I (I6269));
INVX1 gate802(.O (g6352), .I (I8110));
INVX1 gate803(.O (g6818), .I (I8991));
INVX1 gate804(.O (g6577), .I (g6488));
INVX1 gate805(.O (I1847), .I (g209));
INVX1 gate806(.O (I3288), .I (g1710));
INVX1 gate807(.O (g3567), .I (g3074));
INVX1 gate808(.O (I3382), .I (g1284));
INVX1 gate809(.O (g1715), .I (I2716));
INVX1 gate810(.O (g4135), .I (I5487));
INVX1 gate811(.O (I7704), .I (g5723));
INVX1 gate812(.O (g848), .I (g594));
INVX1 gate813(.O (g5092), .I (g4753));
INVX1 gate814(.O (g1498), .I (I2479));
INVX1 gate815(.O (I2763), .I (key_out_120));
INVX1 gate816(.O (g2870), .I (g2296));
INVX1 gate817(.O (I3022), .I (g1426));
INVX1 gate818(.O (I4261), .I (g1857));
INVX1 gate819(.O (I2391), .I (g774));
INVX1 gate820(.O (g4382), .I (I5857));
INVX1 gate821(.O (g3776), .I (g3466));
INVX1 gate822(.O (g6893), .I (I9146));
INVX1 gate823(.O (g1833), .I (I2913));
INVX1 gate824(.O (I3422), .I (g1641));
INVX1 gate825(.O (g5574), .I (g5407));
INVX1 gate826(.O (I3749), .I (g2484));
INVX1 gate827(.O (g3593), .I (g2997));
INVX1 gate828(.O (g6211), .I (g5992));
INVX1 gate829(.O (g2650), .I (I3794));
INVX1 gate830(.O (g5714), .I (I7475));
INVX1 gate831(.O (g932), .I (g337));
INVX1 gate832(.O (I8061), .I (g6113));
INVX1 gate833(.O (g4805), .I (g4473));
INVX1 gate834(.O (g4022), .I (I5328));
INVX1 gate835(.O (g1584), .I (g743));
INVX1 gate836(.O (g4422), .I (g4111));
INVX1 gate837(.O (g6599), .I (I8665));
INVX1 gate838(.O (g1539), .I (g878));
INVX1 gate839(.O (I5109), .I (g3710));
INVX1 gate840(.O (g2408), .I (I3546));
INVX1 gate841(.O (I2159), .I (g465));
INVX1 gate842(.O (I6570), .I (g4719));
INVX1 gate843(.O (g2136), .I (g1395));
INVX1 gate844(.O (I4664), .I (g2924));
INVX1 gate845(.O (I8027), .I (g6237));
INVX1 gate846(.O (I4246), .I (g2194));
INVX1 gate847(.O (g2336), .I (I3488));
INVX1 gate848(.O (g5580), .I (I7336));
INVX1 gate849(.O (g716), .I (I1832));
INVX1 gate850(.O (I3560), .I (g1673));
INVX1 gate851(.O (g736), .I (I1841));
INVX1 gate852(.O (I6525), .I (g4770));
INVX1 gate853(.O (g2768), .I (g2367));
INVX1 gate854(.O (g6370), .I (I8174));
INVX1 gate855(.O (g2594), .I (I3723));
INVX1 gate856(.O (g4798), .I (I6464));
INVX1 gate857(.O (g6325), .I (I8061));
INVX1 gate858(.O (g6821), .I (g6785));
INVX1 gate859(.O (g4560), .I (g4188));
INVX1 gate860(.O (g2806), .I (g2446));
INVX1 gate861(.O (I3632), .I (g1295));
INVX1 gate862(.O (g3450), .I (I4688));
INVX1 gate863(.O (I3037), .I (g1769));
INVX1 gate864(.O (g6939), .I (I9230));
INVX1 gate865(.O (g1052), .I (g668));
INVX1 gate866(.O (I3653), .I (g1305));
INVX1 gate867(.O (I3102), .I (g1426));
INVX1 gate868(.O (I2115), .I (g687));
INVX1 gate869(.O (I2315), .I (key_out_124));
INVX1 gate870(.O (I2811), .I (key_out_128));
INVX1 gate871(.O (g6083), .I (g5809));
INVX1 gate872(.O (g2887), .I (g1858));
INVX1 gate873(.O (I2047), .I (g682));
INVX1 gate874(.O (g6544), .I (I8544));
INVX1 gate875(.O (I6607), .I (g4745));
INVX1 gate876(.O (g4632), .I (g4281));
INVX1 gate877(.O (g5889), .I (g5742));
INVX1 gate878(.O (g5476), .I (I7164));
INVX1 gate879(.O (g2934), .I (g2004));
INVX1 gate880(.O (g2230), .I (I3355));
INVX1 gate881(.O (g4437), .I (I5948));
INVX1 gate882(.O (g4102), .I (I5388));
INVX1 gate883(.O (g4302), .I (g4068));
INVX1 gate884(.O (I5865), .I (g3743));
INVX1 gate885(.O (g6106), .I (I7814));
INVX1 gate886(.O (g4579), .I (g4206));
INVX1 gate887(.O (g4869), .I (g4662));
INVX1 gate888(.O (g6306), .I (I8030));
INVX1 gate889(.O (I3752), .I (g2044));
INVX1 gate890(.O (g5375), .I (I7029));
INVX1 gate891(.O (I8107), .I (g6136));
INVX1 gate892(.O (g4719), .I (I6337));
INVX1 gate893(.O (g1730), .I (g1114));
INVX1 gate894(.O (g3289), .I (g3034));
INVX1 gate895(.O (g1504), .I (I2485));
INVX1 gate896(.O (g3777), .I (g3388));
INVX1 gate897(.O (I6587), .I (g4803));
INVX1 gate898(.O (I8159), .I (g6167));
INVX1 gate899(.O (I6111), .I (g4404));
INVX1 gate900(.O (g3835), .I (I5030));
INVX1 gate901(.O (I6311), .I (g4444));
INVX1 gate902(.O (I8223), .I (g6325));
INVX1 gate903(.O (g2096), .I (I3212));
INVX1 gate904(.O (I9143), .I (g6886));
INVX1 gate905(.O (g3882), .I (I5119));
INVX1 gate906(.O (g1070), .I (g94));
INVX1 gate907(.O (g2550), .I (I3665));
INVX1 gate908(.O (I6615), .I (g4745));
INVX1 gate909(.O (g3271), .I (g3042));
INVX1 gate910(.O (I4671), .I (g2928));
INVX1 gate911(.O (I2880), .I (key_out_123));
INVX1 gate912(.O (g2845), .I (g2565));
INVX1 gate913(.O (g1897), .I (I2992));
INVX1 gate914(.O (g6622), .I (I8724));
INVX1 gate915(.O (I2537), .I (g971));
INVX1 gate916(.O (I5896), .I (g3879));
INVX1 gate917(.O (g2195), .I (I3334));
INVX1 gate918(.O (g4265), .I (I5716));
INVX1 gate919(.O (g2891), .I (g1884));
INVX1 gate920(.O (g2913), .I (g1925));
INVX1 gate921(.O (g5139), .I (I6795));
INVX1 gate922(.O (I3364), .I (g1648));
INVX1 gate923(.O (g5384), .I (g5220));
INVX1 gate924(.O (I9134), .I (g6864));
INVX1 gate925(.O (I2272), .I (g908));
INVX1 gate926(.O (g6904), .I (I9179));
INVX1 gate927(.O (g4786), .I (I6448));
INVX1 gate928(.O (g3799), .I (g3388));
INVX1 gate929(.O (g6514), .I (I8462));
INVX1 gate930(.O (g4364), .I (I5825));
INVX1 gate931(.O (I8447), .I (g6410));
INVX1 gate932(.O (I3770), .I (g2145));
INVX1 gate933(.O (I5019), .I (g3318));
INVX1 gate934(.O (I2417), .I (g774));
INVX1 gate935(.O (g6403), .I (I8223));
INVX1 gate936(.O (g5809), .I (I7608));
INVX1 gate937(.O (I7683), .I (g5702));
INVX1 gate938(.O (g6841), .I (I9044));
INVX1 gate939(.O (g3541), .I (g2643));
INVX1 gate940(.O (I2982), .I (g1426));
INVX1 gate941(.O (g1678), .I (I2658));
INVX1 gate942(.O (g4770), .I (I6414));
INVX1 gate943(.O (g1006), .I (I2047));
INVX1 gate944(.O (I2234), .I (g697));
INVX1 gate945(.O (g1331), .I (I2346));
INVX1 gate946(.O (g4296), .I (I5753));
INVX1 gate947(.O (I2128), .I (g18));
INVX1 gate948(.O (g3238), .I (I4513));
INVX1 gate949(.O (I3553), .I (g1305));
INVX1 gate950(.O (I6020), .I (g4176));
INVX1 gate951(.O (g3332), .I (g3079));
INVX1 gate952(.O (g5477), .I (I7167));
INVX1 gate953(.O (I6420), .I (g4618));
INVX1 gate954(.O (g6695), .I (I8803));
INVX1 gate955(.O (I2330), .I (g1122));
INVX1 gate956(.O (g3209), .I (I4452));
INVX1 gate957(.O (I6507), .I (g4644));
INVX1 gate958(.O (g4532), .I (I6108));
INVX1 gate959(.O (g1682), .I (g829));
INVX1 gate960(.O (g6107), .I (I7817));
INVX1 gate961(.O (I9113), .I (g6855));
INVX1 gate962(.O (I1856), .I (g204));
INVX1 gate963(.O (g1305), .I (I2293));
INVX1 gate964(.O (g6536), .I (I8524));
INVX1 gate965(.O (g3802), .I (g3388));
INVX1 gate966(.O (I5728), .I (g4022));
INVX1 gate967(.O (g2481), .I (I3608));
INVX1 gate968(.O (I7475), .I (g5627));
INVX1 gate969(.O (g931), .I (g54));
INVX1 gate970(.O (g1748), .I (I2763));
INVX1 gate971(.O (g2692), .I (I3840));
INVX1 gate972(.O (I4217), .I (g2163));
INVX1 gate973(.O (g2097), .I (I3215));
INVX1 gate974(.O (I4066), .I (g2582));
INVX1 gate975(.O (g5551), .I (I7295));
INVX1 gate976(.O (g5742), .I (g5686));
INVX1 gate977(.O (g2726), .I (I3886));
INVX1 gate978(.O (g5099), .I (I6737));
INVX1 gate979(.O (g2497), .I (I3626));
INVX1 gate980(.O (I5385), .I (g3962));
INVX1 gate981(.O (g5304), .I (I6956));
INVX1 gate982(.O (g2154), .I (I3271));
INVX1 gate983(.O (g1755), .I (I2776));
INVX1 gate984(.O (g4189), .I (I5597));
INVX1 gate985(.O (I8978), .I (g6792));
INVX1 gate986(.O (g4706), .I (I6308));
INVX1 gate987(.O (g6416), .I (I8258));
INVX1 gate988(.O (I8243), .I (g6286));
INVX1 gate989(.O (I8417), .I (g6420));
INVX1 gate990(.O (g3901), .I (g3575));
INVX1 gate991(.O (I6630), .I (g4745));
INVX1 gate992(.O (I7646), .I (g5774));
INVX1 gate993(.O (I3675), .I (g1491));
INVX1 gate994(.O (g6522), .I (I8482));
INVX1 gate995(.O (g6115), .I (g5879));
INVX1 gate996(.O (g1045), .I (g699));
INVX1 gate997(.O (I3281), .I (g1761));
INVX1 gate998(.O (I7039), .I (g5309));
INVX1 gate999(.O (I7484), .I (g5630));
INVX1 gate1000(.O (g1173), .I (I2185));
INVX1 gate1001(.O (I4455), .I (g2118));
INVX1 gate1002(.O (I8629), .I (g6544));
INVX1 gate1003(.O (g5273), .I (I6930));
INVX1 gate1004(.O (I4133), .I (g2040));
INVX1 gate1005(.O (g1491), .I (I2476));
INVX1 gate1006(.O (g760), .I (I1853));
INVX1 gate1007(.O (g2783), .I (I3979));
INVX1 gate1008(.O (g4281), .I (I5736));
INVX1 gate1009(.O (g3600), .I (I4791));
INVX1 gate1010(.O (g2112), .I (I3240));
INVX1 gate1011(.O (g1283), .I (g853));
INVX1 gate1012(.O (g2312), .I (I3462));
INVX1 gate1013(.O (g1369), .I (I2405));
INVX1 gate1014(.O (I6750), .I (g4771));
INVX1 gate1015(.O (g6654), .I (I8758));
INVX1 gate1016(.O (g3714), .I (g3041));
INVX1 gate1017(.O (I7583), .I (g5605));
INVX1 gate1018(.O (I3684), .I (g1733));
INVX1 gate1019(.O (I5006), .I (g3604));
INVX1 gate1020(.O (I8800), .I (g6684));
INVX1 gate1021(.O (g1059), .I (key_out_40));
INVX1 gate1022(.O (g1578), .I (I2552));
INVX1 gate1023(.O (g2001), .I (I3112));
INVX1 gate1024(.O (I5406), .I (g3976));
INVX1 gate1025(.O (g5572), .I (g5399));
INVX1 gate1026(.O (I3109), .I (g1504));
INVX1 gate1027(.O (I3791), .I (g2044));
INVX1 gate1028(.O (g2293), .I (g1567));
INVX1 gate1029(.O (g6880), .I (I9107));
INVX1 gate1030(.O (g6595), .I (I8653));
INVX1 gate1031(.O (g4138), .I (I5496));
INVX1 gate1032(.O (g1535), .I (g1088));
INVX1 gate1033(.O (g4639), .I (g4289));
INVX1 gate1034(.O (g6537), .I (I8527));
INVX1 gate1035(.O (g5543), .I (g5331));
INVX1 gate1036(.O (I3808), .I (g2125));
INVX1 gate1037(.O (I7276), .I (g5375));
INVX1 gate1038(.O (I5487), .I (g3881));
INVX1 gate1039(.O (I2355), .I (key_out_125));
INVX1 gate1040(.O (g4109), .I (I5409));
INVX1 gate1041(.O (g4309), .I (g4074));
INVX1 gate1042(.O (g2828), .I (g2488));
INVX1 gate1043(.O (g2830), .I (g2494));
INVX1 gate1044(.O (g2727), .I (g2324));
INVX1 gate1045(.O (g4808), .I (g4473));
INVX1 gate1046(.O (I2964), .I (g1257));
INVX1 gate1047(.O (g821), .I (I1880));
INVX1 gate1048(.O (g6612), .I (I8702));
INVX1 gate1049(.O (g5534), .I (I7276));
INVX1 gate1050(.O (g5729), .I (I7494));
INVX1 gate1051(.O (I6666), .I (g4740));
INVX1 gate1052(.O (I9179), .I (g6875));
INVX1 gate1053(.O (g1415), .I (g1246));
INVX1 gate1054(.O (g4707), .I (I6311));
INVX1 gate1055(.O (g6417), .I (I8261));
INVX1 gate1056(.O (I7404), .I (g5541));
INVX1 gate1057(.O (g3076), .I (I4309));
INVX1 gate1058(.O (I8512), .I (g6441));
INVX1 gate1059(.O (g3889), .I (g3575));
INVX1 gate1060(.O (I6528), .I (g4815));
INVX1 gate1061(.O (g1664), .I (I2643));
INVX1 gate1062(.O (g1246), .I (I2237));
INVX1 gate1063(.O (g6234), .I (g6057));
INVX1 gate1064(.O (I3575), .I (g1305));
INVX1 gate1065(.O (g5885), .I (g5865));
INVX1 gate1066(.O (g6328), .I (I8066));
INVX1 gate1067(.O (g1203), .I (I2207));
INVX1 gate1068(.O (I5445), .I (g4040));
INVX1 gate1069(.O (g5946), .I (g5729));
INVX1 gate1070(.O (g6542), .I (I8538));
INVX1 gate1071(.O (g6330), .I (I8070));
INVX1 gate1072(.O (g1721), .I (I2721));
INVX1 gate1073(.O (I5091), .I (g3242));
INVX1 gate1074(.O (I8056), .I (g6109));
INVX1 gate1075(.O (g2932), .I (g1998));
INVX1 gate1076(.O (I8456), .I (g6417));
INVX1 gate1077(.O (g5903), .I (g5753));
INVX1 gate1078(.O (I3833), .I (g2266));
INVX1 gate1079(.O (I2318), .I (key_out_120));
INVX1 gate1080(.O (g4715), .I (I6327));
INVX1 gate1081(.O (I2367), .I (key_out_126));
INVX1 gate1082(.O (I1924), .I (g663));
INVX1 gate1083(.O (g6800), .I (I8966));
INVX1 gate1084(.O (I5169), .I (key_out_6));
INVX1 gate1085(.O (I6410), .I (g4473));
INVX1 gate1086(.O (g4098), .I (I5376));
INVX1 gate1087(.O (g3500), .I (g2647));
INVX1 gate1088(.O (g4498), .I (I6012));
INVX1 gate1089(.O (I2057), .I (g685));
INVX1 gate1090(.O (g1502), .I (g709));
INVX1 gate1091(.O (I5059), .I (g3259));
INVX1 gate1092(.O (I5920), .I (g4228));
INVX1 gate1093(.O (I2457), .I (g1253));
INVX1 gate1094(.O (I3584), .I (g1678));
INVX1 gate1095(.O (I5868), .I (g3864));
INVX1 gate1096(.O (I2989), .I (g1519));
INVX1 gate1097(.O (I2193), .I (g693));
INVX1 gate1098(.O (g5436), .I (I7116));
INVX1 gate1099(.O (g3384), .I (g2834));
INVX1 gate1100(.O (g1940), .I (I3047));
INVX1 gate1101(.O (g2576), .I (I3687));
INVX1 gate1102(.O (g2866), .I (g1905));
INVX1 gate1103(.O (g5135), .I (I6783));
INVX1 gate1104(.O (g2716), .I (I3871));
INVX1 gate1105(.O (g3838), .I (I5037));
INVX1 gate1106(.O (I7906), .I (g5912));
INVX1 gate1107(.O (I3268), .I (g1656));
INVX1 gate1108(.O (I3019), .I (g1755));
INVX1 gate1109(.O (g3424), .I (I4671));
INVX1 gate1110(.O (g5382), .I (I7042));
INVX1 gate1111(.O (I5793), .I (g3803));
INVX1 gate1112(.O (I3419), .I (g1287));
INVX1 gate1113(.O (g6902), .I (I9173));
INVX1 gate1114(.O (I6143), .I (g4237));
INVX1 gate1115(.O (I6343), .I (g4458));
INVX1 gate1116(.O (g846), .I (g586));
INVX1 gate1117(.O (g1671), .I (g985));
INVX1 gate1118(.O (g5805), .I (I7604));
INVX1 gate1119(.O (I5415), .I (g3723));
INVX1 gate1120(.O (g6512), .I (I8456));
INVX1 gate1121(.O (I3452), .I (g1450));
INVX1 gate1122(.O (g4162), .I (I5562));
INVX1 gate1123(.O (g5022), .I (I6666));
INVX1 gate1124(.O (g1030), .I (I2057));
INVX1 gate1125(.O (I8279), .I (g6307));
INVX1 gate1126(.O (g3231), .I (I4492));
INVX1 gate1127(.O (g6490), .I (g6371));
INVX1 gate1128(.O (I2321), .I (g898));
INVX1 gate1129(.O (g6823), .I (I9002));
INVX1 gate1130(.O (g3477), .I (g2692));
INVX1 gate1131(.O (g6166), .I (I7892));
INVX1 gate1132(.O (g6366), .I (I8162));
INVX1 gate1133(.O (I6334), .I (g4454));
INVX1 gate1134(.O (I8872), .I (g6695));
INVX1 gate1135(.O (g2241), .I (I3370));
INVX1 gate1136(.O (g1564), .I (g1030));
INVX1 gate1137(.O (I7892), .I (g5916));
INVX1 gate1138(.O (I3086), .I (g1439));
INVX1 gate1139(.O (g6529), .I (I8503));
INVX1 gate1140(.O (I8843), .I (g6658));
INVX1 gate1141(.O (g6649), .I (I8745));
INVX1 gate1142(.O (I6555), .I (g4703));
INVX1 gate1143(.O (g1741), .I (I2753));
INVX1 gate1144(.O (I6792), .I (g5097));
INVX1 gate1145(.O (g3104), .I (I4351));
INVX1 gate1146(.O (I3385), .I (g1318));
INVX1 gate1147(.O (g2524), .I (I3647));
INVX1 gate1148(.O (g2644), .I (I3788));
INVX1 gate1149(.O (I8834), .I (g6661));
INVX1 gate1150(.O (g6698), .I (I8812));
INVX1 gate1151(.O (g1638), .I (g754));
INVX1 gate1152(.O (g839), .I (key_out_32));
INVX1 gate1153(.O (I6621), .I (g4745));
INVX1 gate1154(.O (g2119), .I (g1391));
INVX1 gate1155(.O (I5502), .I (g3853));
INVX1 gate1156(.O (g1108), .I (I2134));
INVX1 gate1157(.O (I3025), .I (g1439));
INVX1 gate1158(.O (I2552), .I (g971));
INVX1 gate1159(.O (g5437), .I (I7119));
INVX1 gate1160(.O (g4385), .I (I5862));
INVX1 gate1161(.O (I3425), .I (g1274));
INVX1 gate1162(.O (I9092), .I (g6855));
INVX1 gate1163(.O (I4441), .I (g2109));
INVX1 gate1164(.O (g2818), .I (g2464));
INVX1 gate1165(.O (g2867), .I (g1908));
INVX1 gate1166(.O (g1883), .I (g1797));
INVX1 gate1167(.O (g5579), .I (I7333));
INVX1 gate1168(.O (I7478), .I (g5628));
INVX1 gate1169(.O (g4425), .I (I5926));
INVX1 gate1170(.O (I7035), .I (g5150));
INVX1 gate1171(.O (I5388), .I (g3969));
INVX1 gate1172(.O (I7517), .I (g5593));
INVX1 gate1173(.O (g2893), .I (g1985));
INVX1 gate1174(.O (g5752), .I (I7509));
INVX1 gate1175(.O (I8232), .I (g6332));
INVX1 gate1176(.O (g5917), .I (I7683));
INVX1 gate1177(.O (I6567), .I (g4715));
INVX1 gate1178(.O (g6720), .I (I8854));
INVX1 gate1179(.O (I3678), .I (g1690));
INVX1 gate1180(.O (g2975), .I (I4176));
INVX1 gate1181(.O (I5030), .I (g3242));
INVX1 gate1182(.O (I3331), .I (g1631));
INVX1 gate1183(.O (g1861), .I (I2967));
INVX1 gate1184(.O (g6367), .I (I8165));
INVX1 gate1185(.O (g1048), .I (g492));
INVX1 gate1186(.O (I5430), .I (g3727));
INVX1 gate1187(.O (g2599), .I (I3729));
INVX1 gate1188(.O (g5042), .I (I6672));
INVX1 gate1189(.O (g1711), .I (I2712));
INVX1 gate1190(.O (I3635), .I (g1305));
INVX1 gate1191(.O (g6652), .I (I8752));
INVX1 gate1192(.O (g5442), .I (g5270));
INVX1 gate1193(.O (g1055), .I (g269));
INVX1 gate1194(.O (I2570), .I (key_out_124));
INVX1 gate1195(.O (I2860), .I (key_out_125));
INVX1 gate1196(.O (g6057), .I (g5824));
INVX1 gate1197(.O (g4131), .I (I5475));
INVX1 gate1198(.O (I4743), .I (g2594));
INVX1 gate1199(.O (I3105), .I (g1439));
INVX1 gate1200(.O (g2170), .I (I3301));
INVX1 gate1201(.O (g2370), .I (I3522));
INVX1 gate1202(.O (g4406), .I (I5913));
INVX1 gate1203(.O (g6193), .I (g5957));
INVX1 gate1204(.O (g1333), .I (I2352));
INVX1 gate1205(.O (g2125), .I (I3255));
INVX1 gate1206(.O (I8552), .I (g6455));
INVX1 gate1207(.O (g1774), .I (I2817));
INVX1 gate1208(.O (g4766), .I (I6406));
INVX1 gate1209(.O (g4105), .I (I5397));
INVX1 gate1210(.O (g1846), .I (I2940));
INVX1 gate1211(.O (g5054), .I (g4816));
INVX1 gate1212(.O (g4801), .I (g4487));
INVX1 gate1213(.O (g6834), .I (g6821));
INVX1 gate1214(.O (g4487), .I (I5991));
INVX1 gate1215(.O (I7110), .I (g5291));
INVX1 gate1216(.O (g3534), .I (I4752));
INVX1 gate1217(.O (I5910), .I (g3750));
INVX1 gate1218(.O (g5770), .I (g5645));
INVX1 gate1219(.O (I3755), .I (g2125));
INVX1 gate1220(.O (g5296), .I (I6946));
INVX1 gate1221(.O (I8687), .I (g6568));
INVX1 gate1222(.O (I6933), .I (g5124));
INVX1 gate1223(.O (g2544), .I (I3662));
INVX1 gate1224(.O (g6598), .I (I8662));
INVX1 gate1225(.O (I5609), .I (g3893));
INVX1 gate1226(.O (I4474), .I (g3052));
INVX1 gate1227(.O (I2358), .I (g1176));
INVX1 gate1228(.O (g3014), .I (I4217));
INVX1 gate1229(.O (g6121), .I (I7835));
INVX1 gate1230(.O (I7002), .I (g5308));
INVX1 gate1231(.O (g766), .I (I1856));
INVX1 gate1232(.O (g3885), .I (I5124));
INVX1 gate1233(.O (g4226), .I (g4050));
INVX1 gate1234(.O (g2106), .I (g1378));
INVX1 gate1235(.O (g2306), .I (g1743));
INVX1 gate1236(.O (I3373), .I (g1320));
INVX1 gate1237(.O (g2790), .I (g2413));
INVX1 gate1238(.O (g6232), .I (g6048));
INVX1 gate1239(.O (I5217), .I (key_out_11));
INVX1 gate1240(.O (I8570), .I (g6433));
INVX1 gate1241(.O (I8860), .I (g6699));
INVX1 gate1242(.O (I4480), .I (g3073));
INVX1 gate1243(.O (g1994), .I (I3105));
INVX1 gate1244(.O (g1290), .I (I2275));
INVX1 gate1245(.O (I2275), .I (g909));
INVX1 gate1246(.O (g6938), .I (I9227));
INVX1 gate1247(.O (I5466), .I (g3787));
INVX1 gate1248(.O (g4173), .I (I5577));
INVX1 gate1249(.O (I8710), .I (g6517));
INVX1 gate1250(.O (g2461), .I (I3593));
INVX1 gate1251(.O (I7590), .I (g5605));
INVX1 gate1252(.O (I3602), .I (g1491));
INVX1 gate1253(.O (I3007), .I (g1439));
INVX1 gate1254(.O (g2756), .I (g2353));
INVX1 gate1255(.O (g2622), .I (I3764));
INVX1 gate1256(.O (I3059), .I (g1519));
INVX1 gate1257(.O (I3578), .I (g1484));
INVX1 gate1258(.O (I3868), .I (g2125));
INVX1 gate1259(.O (g5888), .I (g5731));
INVX1 gate1260(.O (g1256), .I (g838));
INVX1 gate1261(.O (g6519), .I (I8473));
INVX1 gate1262(.O (I6289), .I (g4433));
INVX1 gate1263(.O (I9024), .I (g6803));
INVX1 gate1264(.O (I5448), .I (g3960));
INVX1 gate1265(.O (I3767), .I (g2125));
INVX1 gate1266(.O (g5787), .I (g5685));
INVX1 gate1267(.O (g2904), .I (g1991));
INVX1 gate1268(.O (g6552), .I (I8552));
INVX1 gate1269(.O (g6606), .I (I8684));
INVX1 gate1270(.O (g2446), .I (I3581));
INVX1 gate1271(.O (I5333), .I (key_out_10));
INVX1 gate1272(.O (I2284), .I (g922));
INVX1 gate1273(.O (g1381), .I (I2417));
INVX1 gate1274(.O (g4718), .I (I6334));
INVX1 gate1275(.O (g4767), .I (g4601));
INVX1 gate1276(.O (I3261), .I (g1783));
INVX1 gate1277(.O (g1847), .I (I2943));
INVX1 gate1278(.O (I4688), .I (g3207));
INVX1 gate1279(.O (I5774), .I (g3807));
INVX1 gate1280(.O (I9077), .I (g6845));
INVX1 gate1281(.O (I8659), .I (g6523));
INVX1 gate1282(.O (g4535), .I (g4173));
INVX1 gate1283(.O (I4976), .I (g3575));
INVX1 gate1284(.O (g1685), .I (I2671));
INVX1 gate1285(.O (g2145), .I (I3268));
INVX1 gate1286(.O (I8506), .I (g6483));
INVX1 gate1287(.O (g2841), .I (g2541));
INVX1 gate1288(.O (g4582), .I (g4210));
INVX1 gate1289(.O (g3022), .I (I4229));
INVX1 gate1290(.O (g2391), .I (I3534));
INVX1 gate1291(.O (g6586), .I (I8626));
INVX1 gate1292(.O (g952), .I (I2029));
INVX1 gate1293(.O (g1263), .I (g846));
INVX1 gate1294(.O (g964), .I (g357));
INVX1 gate1295(.O (I2420), .I (g791));
INVX1 gate1296(.O (g2695), .I (I3843));
INVX1 gate1297(.O (g2637), .I (I3779));
INVX1 gate1298(.O (g1950), .I (I3059));
INVX1 gate1299(.O (g5138), .I (I6792));
INVX1 gate1300(.O (g4227), .I (g4059));
INVX1 gate1301(.O (I7295), .I (g5439));
INVX1 gate1302(.O (g5791), .I (I7590));
INVX1 gate1303(.O (g3798), .I (g3388));
INVX1 gate1304(.O (I9104), .I (g6864));
INVX1 gate1305(.O (g5309), .I (g5063));
INVX1 gate1306(.O (g2159), .I (I3284));
INVX1 gate1307(.O (g6570), .I (I8594));
INVX1 gate1308(.O (g4246), .I (I5692));
INVX1 gate1309(.O (I6132), .I (g4219));
INVX1 gate1310(.O (I8174), .I (g6173));
INVX1 gate1311(.O (g6525), .I (I8491));
INVX1 gate1312(.O (g6710), .I (I8840));
INVX1 gate1313(.O (I5418), .I (g4036));
INVX1 gate1314(.O (I6680), .I (g4713));
INVX1 gate1315(.O (g4721), .I (I6343));
INVX1 gate1316(.O (g1631), .I (I2588));
INVX1 gate1317(.O (g2416), .I (I3556));
INVX1 gate1318(.O (g3095), .I (I4340));
INVX1 gate1319(.O (g3037), .I (I4252));
INVX1 gate1320(.O (I3502), .I (g1295));
INVX1 gate1321(.O (g1257), .I (g845));
INVX1 gate1322(.O (g1101), .I (I2125));
INVX1 gate1323(.O (I2204), .I (g694));
INVX1 gate1324(.O (I2630), .I (key_out_123));
INVX1 gate1325(.O (I5493), .I (g3834));
INVX1 gate1326(.O (I8180), .I (g6176));
INVX1 gate1327(.O (I4220), .I (g2164));
INVX1 gate1328(.O (I7966), .I (g6166));
INVX1 gate1329(.O (I8591), .I (g6448));
INVX1 gate1330(.O (g2315), .I (I3465));
INVX1 gate1331(.O (g5957), .I (g5866));
INVX1 gate1332(.O (g6879), .I (I9104));
INVX1 gate1333(.O (g6607), .I (I8687));
INVX1 gate1334(.O (I6558), .I (g4705));
INVX1 gate1335(.O (g4502), .I (I6020));
INVX1 gate1336(.O (g5049), .I (I6685));
INVX1 gate1337(.O (I9044), .I (g6836));
INVX1 gate1338(.O (g927), .I (I1958));
INVX1 gate1339(.O (I1942), .I (g664));
INVX1 gate1340(.O (I4023), .I (g2315));
INVX1 gate1341(.O (g3719), .I (g3053));
INVX1 gate1342(.O (g6506), .I (I8438));
INVX1 gate1343(.O (g5575), .I (g5411));
INVX1 gate1344(.O (I8420), .I (g6422));
INVX1 gate1345(.O (I3388), .I (g1324));
INVX1 gate1346(.O (g2874), .I (g1849));
INVX1 gate1347(.O (g3752), .I (I4935));
INVX1 gate1348(.O (I5397), .I (g3932));
INVX1 gate1349(.O (I3028), .I (g1504));
INVX1 gate1350(.O (g4188), .I (I5594));
INVX1 gate1351(.O (g6587), .I (I8629));
INVX1 gate1352(.O (g4388), .I (I5871));
INVX1 gate1353(.O (I5421), .I (g3724));
INVX1 gate1354(.O (I3428), .I (g1825));
INVX1 gate1355(.O (I2973), .I (g1687));
INVX1 gate1356(.O (I7254), .I (g5458));
INVX1 gate1357(.O (I7814), .I (g5922));
INVX1 gate1358(.O (I3247), .I (g1791));
INVX1 gate1359(.O (g3042), .I (I4261));
INVX1 gate1360(.O (g6615), .I (I8707));
INVX1 gate1361(.O (I7150), .I (g5355));
INVX1 gate1362(.O (I4327), .I (g2525));
INVX1 gate1363(.O (g4428), .I (I5933));
INVX1 gate1364(.O (g3786), .I (g3388));
INVX1 gate1365(.O (g5584), .I (I7346));
INVX1 gate1366(.O (g5539), .I (g5331));
INVX1 gate1367(.O (g5896), .I (g5753));
INVX1 gate1368(.O (g1673), .I (I2653));
INVX1 gate1369(.O (g6374), .I (I8186));
INVX1 gate1370(.O (I3826), .I (g2145));
INVX1 gate1371(.O (g3364), .I (g3114));
INVX1 gate1372(.O (g3233), .I (I4498));
INVX1 gate1373(.O (I8515), .I (g6492));
INVX1 gate1374(.O (g4564), .I (g4192));
INVX1 gate1375(.O (g3054), .I (I4279));
INVX1 gate1376(.O (I5562), .I (g4002));
INVX1 gate1377(.O (I4303), .I (g1897));
INVX1 gate1378(.O (g2612), .I (I3752));
INVX1 gate1379(.O (I8300), .I (g6299));
INVX1 gate1380(.O (g6284), .I (I8002));
INVX1 gate1381(.O (g2243), .I (I3376));
INVX1 gate1382(.O (g3770), .I (I4961));
INVX1 gate1383(.O (I9014), .I (g6820));
INVX1 gate1384(.O (I3638), .I (g1484));
INVX1 gate1385(.O (g1772), .I (I2811));
INVX1 gate1386(.O (I5723), .I (g3942));
INVX1 gate1387(.O (g4741), .I (I6371));
INVX1 gate1388(.O (g6591), .I (I8641));
INVX1 gate1389(.O (g5052), .I (I6692));
INVX1 gate1390(.O (g6832), .I (I9021));
INVX1 gate1391(.O (g4910), .I (I6612));
INVX1 gate1392(.O (I2648), .I (g980));
INVX1 gate1393(.O (g2234), .I (I3367));
INVX1 gate1394(.O (g6853), .I (I9082));
INVX1 gate1395(.O (g1890), .I (g1359));
INVX1 gate1396(.O (I3883), .I (g2574));
INVX1 gate1397(.O (g6420), .I (I8270));
INVX1 gate1398(.O (I4240), .I (g2165));
INVX1 gate1399(.O (g2330), .I (g1777));
INVX1 gate1400(.O (g4108), .I (I5406));
INVX1 gate1401(.O (g4609), .I (I6182));
INVX1 gate1402(.O (g6507), .I (I8441));
INVX1 gate1403(.O (g4308), .I (I5777));
INVX1 gate1404(.O (g1011), .I (I2050));
INVX1 gate1405(.O (g1734), .I (g952));
INVX1 gate1406(.O (I3758), .I (g2041));
INVX1 gate1407(.O (g5086), .I (g4732));
INVX1 gate1408(.O (g897), .I (g41));
INVX1 gate1409(.O (I8040), .I (g6142));
INVX1 gate1410(.O (g951), .I (g84));
INVX1 gate1411(.O (I8969), .I (g6797));
INVX1 gate1412(.O (g2800), .I (g2430));
INVX1 gate1413(.O (g5730), .I (I7497));
INVX1 gate1414(.O (g2554), .I (I3669));
INVX1 gate1415(.O (g4758), .I (I6382));
INVX1 gate1416(.O (I2839), .I (key_out_122));
INVX1 gate1417(.O (I3861), .I (g1834));
INVX1 gate1418(.O (g6905), .I (I9182));
INVX1 gate1419(.O (g3029), .I (I4240));
INVX1 gate1420(.O (I3711), .I (g1848));
INVX1 gate1421(.O (I9182), .I (g6879));
INVX1 gate1422(.O (g3787), .I (I4986));
INVX1 gate1423(.O (g2213), .I (I3346));
INVX1 gate1424(.O (g5897), .I (g5731));
INVX1 gate1425(.O (g5025), .I (g4814));
INVX1 gate1426(.O (g6515), .I (g6408));
INVX1 gate1427(.O (g4861), .I (I6587));
INVX1 gate1428(.O (g5425), .I (I7091));
INVX1 gate1429(.O (I4347), .I (g2555));
INVX1 gate1430(.O (I2172), .I (g691));
INVX1 gate1431(.O (I2278), .I (g917));
INVX1 gate1432(.O (g4711), .I (I6315));
INVX1 gate1433(.O (g6100), .I (I7796));
INVX1 gate1434(.O (I4681), .I (g2947));
INVX1 gate1435(.O (g1480), .I (g985));
INVX1 gate1436(.O (g2902), .I (g1899));
INVX1 gate1437(.O (I8875), .I (g6697));
INVX1 gate1438(.O (I2143), .I (g2));
INVX1 gate1439(.O (I2343), .I (key_out_125));
INVX1 gate1440(.O (I6139), .I (g4222));
INVX1 gate1441(.O (g4133), .I (I5481));
INVX1 gate1442(.O (g3297), .I (g3046));
INVX1 gate1443(.O (g2512), .I (I3638));
INVX1 gate1444(.O (g2090), .I (I3206));
INVX1 gate1445(.O (g4846), .I (I6546));
INVX1 gate1446(.O (I2134), .I (g705));
INVX1 gate1447(.O (I6795), .I (g5022));
INVX1 gate1448(.O (I6737), .I (g4662));
INVX1 gate1449(.O (I2334), .I (key_out_127));
INVX1 gate1450(.O (I6809), .I (g5051));
INVX1 gate1451(.O (I5743), .I (g4022));
INVX1 gate1452(.O (g5331), .I (I6995));
INVX1 gate1453(.O (I5890), .I (g3878));
INVX1 gate1454(.O (I3509), .I (g1461));
INVX1 gate1455(.O (g3963), .I (I5217));
INVX1 gate1456(.O (g3791), .I (g3388));
INVX1 gate1457(.O (I8884), .I (g6704));
INVX1 gate1458(.O (I5505), .I (g3860));
INVX1 gate1459(.O (g1688), .I (I2688));
INVX1 gate1460(.O (I6672), .I (g4752));
INVX1 gate1461(.O (g4780), .I (I6434));
INVX1 gate1462(.O (g6040), .I (g5824));
INVX1 gate1463(.O (g1857), .I (I2961));
INVX1 gate1464(.O (I6231), .I (g4350));
INVX1 gate1465(.O (I3662), .I (g1688));
INVX1 gate1466(.O (g4509), .I (I6039));
INVX1 gate1467(.O (g5087), .I (g4736));
INVX1 gate1468(.O (I9095), .I (g6855));
INVX1 gate1469(.O (g5801), .I (I7600));
INVX1 gate1470(.O (g2155), .I (I3274));
INVX1 gate1471(.O (I9208), .I (g6922));
INVX1 gate1472(.O (g4662), .I (g4640));
INVX1 gate1473(.O (I3093), .I (g1426));
INVX1 gate1474(.O (g965), .I (I2033));
INVX1 gate1475(.O (I3493), .I (g1461));
INVX1 gate1476(.O (I3816), .I (g2580));
INVX1 gate1477(.O (g1326), .I (g894));
INVX1 gate1478(.O (I8235), .I (g6312));
INVX1 gate1479(.O (I6099), .I (g4398));
INVX1 gate1480(.O (I8282), .I (g6309));
INVX1 gate1481(.O (g3049), .I (I4270));
INVX1 gate1482(.O (g6528), .I (I8500));
INVX1 gate1483(.O (g1760), .I (I2785));
INVX1 gate1484(.O (g4493), .I (I6001));
INVX1 gate1485(.O (g6351), .I (I8107));
INVX1 gate1486(.O (I1850), .I (g210));
INVX1 gate1487(.O (g6875), .I (I9092));
INVX1 gate1488(.O (g834), .I (g341));
INVX1 gate1489(.O (I8988), .I (g6787));
INVX1 gate1490(.O (g6530), .I (I8506));
INVX1 gate1491(.O (g3575), .I (I4777));
INVX1 gate1492(.O (g5045), .I (I6677));
INVX1 gate1493(.O (I8693), .I (g6570));
INVX1 gate1494(.O (g6655), .I (I8761));
INVX1 gate1495(.O (g5445), .I (g5274));
INVX1 gate1496(.O (I5713), .I (g4022));
INVX1 gate1497(.O (g3604), .I (I4799));
INVX1 gate1498(.O (I8548), .I (g6454));
INVX1 gate1499(.O (g5491), .I (I7193));
INVX1 gate1500(.O (g3498), .I (g2634));
INVX1 gate1501(.O (g4381), .I (I5854));
INVX1 gate1502(.O (g4847), .I (I6549));
INVX1 gate1503(.O (g2118), .I (I3247));
INVX1 gate1504(.O (g2619), .I (I3761));
INVX1 gate1505(.O (I8555), .I (g6456));
INVX1 gate1506(.O (g2367), .I (I3519));
INVX1 gate1507(.O (g2872), .I (g1922));
INVX1 gate1508(.O (g1608), .I (I2570));
INVX1 gate1509(.O (g1220), .I (I2221));
INVX1 gate1510(.O (g4700), .I (I6292));
INVX1 gate1511(.O (g6410), .I (I8240));
INVX1 gate1512(.O (I9164), .I (g6885));
INVX1 gate1513(.O (g4397), .I (I5890));
INVX1 gate1514(.O (I9233), .I (g6938));
INVX1 gate1515(.O (I2776), .I (g1192));
INVX1 gate1516(.O (I7640), .I (g5773));
INVX1 gate1517(.O (g5407), .I (I7073));
INVX1 gate1518(.O (g6884), .I (I9119));
INVX1 gate1519(.O (I2593), .I (key_out_125));
INVX1 gate1520(.O (g5059), .I (I6697));
INVX1 gate1521(.O (g5920), .I (I7692));
INVX1 gate1522(.O (g6839), .I (I9038));
INVX1 gate1523(.O (g2457), .I (I3587));
INVX1 gate1524(.O (g5578), .I (g5425));
INVX1 gate1525(.O (I6444), .I (g4503));
INVX1 gate1526(.O (I6269), .I (g4655));
INVX1 gate1527(.O (g1423), .I (I2442));
INVX1 gate1528(.O (g923), .I (g332));
INVX1 gate1529(.O (I5857), .I (g3740));
INVX1 gate1530(.O (I7176), .I (g5437));
INVX1 gate1531(.O (g1588), .I (g798));
INVX1 gate1532(.O (I8113), .I (g6147));
INVX1 gate1533(.O (g5582), .I (I7342));
INVX1 gate1534(.O (g1161), .I (I2182));
INVX1 gate1535(.O (g6278), .I (I7966));
INVX1 gate1536(.O (g2686), .I (I3830));
INVX1 gate1537(.O (g6372), .I (I8180));
INVX1 gate1538(.O (g3162), .I (I4402));
INVX1 gate1539(.O (g5261), .I (I6918));
INVX1 gate1540(.O (g3019), .I (I4226));
INVX1 gate1541(.O (I4294), .I (g2525));
INVX1 gate1542(.O (I6543), .I (g4718));
INVX1 gate1543(.O (g6618), .I (I8716));
INVX1 gate1544(.O (g1665), .I (g985));
INVX1 gate1545(.O (I7829), .I (g5926));
INVX1 gate1546(.O (I3723), .I (g2158));
INVX1 gate1547(.O (g6143), .I (I7865));
INVX1 gate1548(.O (g4562), .I (I6132));
INVX1 gate1549(.O (g6235), .I (g6062));
INVX1 gate1550(.O (g2598), .I (I3726));
INVX1 gate1551(.O (g3052), .I (I4273));
INVX1 gate1552(.O (g1327), .I (I2334));
INVX1 gate1553(.O (I2521), .I (g1063));
INVX1 gate1554(.O (I3301), .I (g1730));
INVX1 gate1555(.O (g5415), .I (I7081));
INVX1 gate1556(.O (g3452), .I (g2625));
INVX1 gate1557(.O (g6282), .I (I7996));
INVX1 gate1558(.O (I2050), .I (g683));
INVX1 gate1559(.O (I5400), .I (g3963));
INVX1 gate1560(.O (g6566), .I (I8582));
INVX1 gate1561(.O (I8494), .I (g6428));
INVX1 gate1562(.O (I4501), .I (g2705));
INVX1 gate1563(.O (I6534), .I (g4706));
INVX1 gate1564(.O (I8518), .I (g6494));
INVX1 gate1565(.O (I3605), .I (g1681));
INVX1 gate1566(.O (g4723), .I (I6349));
INVX1 gate1567(.O (I8567), .I (g6432));
INVX1 gate1568(.O (g4101), .I (I5385));
INVX1 gate1569(.O (g6134), .I (I7852));
INVX1 gate1570(.O (g5664), .I (g5521));
INVX1 gate1571(.O (g2625), .I (I3767));
INVX1 gate1572(.O (I7270), .I (g5352));
INVX1 gate1573(.O (g2232), .I (I3361));
INVX1 gate1574(.O (g6548), .I (I8548));
INVX1 gate1575(.O (I6927), .I (g5124));
INVX1 gate1576(.O (g3086), .I (I4327));
INVX1 gate1577(.O (I2724), .I (g1220));
INVX1 gate1578(.O (g2253), .I (I3388));
INVX1 gate1579(.O (I2179), .I (g293));
INVX1 gate1580(.O (g3486), .I (g2869));
INVX1 gate1581(.O (g2813), .I (g2457));
INVX1 gate1582(.O (I2379), .I (key_out_122));
INVX1 gate1583(.O (g1696), .I (I2700));
INVX1 gate1584(.O (I7073), .I (g5281));
INVX1 gate1585(.O (I7796), .I (g5917));
INVX1 gate1586(.O (I6885), .I (g4872));
INVX1 gate1587(.O (I6414), .I (g4497));
INVX1 gate1588(.O (g3504), .I (g2675));
INVX1 gate1589(.O (I6946), .I (g5124));
INVX1 gate1590(.O (g1732), .I (I2738));
INVX1 gate1591(.O (g3881), .I (I5116));
INVX1 gate1592(.O (g2740), .I (I3909));
INVX1 gate1593(.O (I2658), .I (g1001));
INVX1 gate1594(.O (I3441), .I (g1502));
INVX1 gate1595(.O (I7069), .I (g5281));
INVX1 gate1596(.O (g3070), .I (I4297));
INVX1 gate1597(.O (I8264), .I (g6296));
INVX1 gate1598(.O (g6621), .I (I8721));
INVX1 gate1599(.O (I2835), .I (key_out_128));
INVX1 gate1600(.O (I7469), .I (g5625));
INVX1 gate1601(.O (g3897), .I (g3251));
INVX1 gate1602(.O (I5023), .I (g3263));
INVX1 gate1603(.O (g1472), .I (g952));
INVX1 gate1604(.O (g1043), .I (g486));
INVX1 gate1605(.O (I5977), .I (g4319));
INVX1 gate1606(.O (I8521), .I (g6495));
INVX1 gate1607(.O (I6036), .I (g4370));
INVX1 gate1608(.O (I8641), .I (g6524));
INVX1 gate1609(.O (I2611), .I (key_out_128));
INVX1 gate1610(.O (g893), .I (g23));
INVX1 gate1611(.O (g2687), .I (I3833));
INVX1 gate1612(.O (I8450), .I (g6412));
INVX1 gate1613(.O (I3669), .I (g1739));
INVX1 gate1614(.O (g1116), .I (I2154));
INVX1 gate1615(.O (g2586), .I (I3711));
INVX1 gate1616(.O (I3531), .I (g1593));
INVX1 gate1617(.O (I5451), .I (g3967));
INVX1 gate1618(.O (I6182), .I (g4249));
INVX1 gate1619(.O (g6518), .I (I8470));
INVX1 gate1620(.O (g6567), .I (I8585));
INVX1 gate1621(.O (I8724), .I (g6533));
INVX1 gate1622(.O (I6382), .I (g4460));
INVX1 gate1623(.O (g996), .I (I2041));
INVX1 gate1624(.O (g3331), .I (g3076));
INVX1 gate1625(.O (I3890), .I (g2145));
INVX1 gate1626(.O (g4772), .I (I6420));
INVX1 gate1627(.O (g5247), .I (g4900));
INVX1 gate1628(.O (g4531), .I (I6105));
INVX1 gate1629(.O (I5633), .I (g3768));
INVX1 gate1630(.O (I8878), .I (g6710));
INVX1 gate1631(.O (g1681), .I (I2663));
INVX1 gate1632(.O (I3505), .I (g1305));
INVX1 gate1633(.O (g6593), .I (I8647));
INVX1 gate1634(.O (g3766), .I (I4955));
INVX1 gate1635(.O (g1533), .I (g878));
INVX1 gate1636(.O (g5564), .I (g5382));
INVX1 gate1637(.O (I5103), .I (g3440));
INVX1 gate1638(.O (g2525), .I (I3650));
INVX1 gate1639(.O (g3801), .I (g3388));
INVX1 gate1640(.O (g3487), .I (g2622));
INVX1 gate1641(.O (g1914), .I (I3013));
INVX1 gate1642(.O (I5696), .I (g3942));
INVX1 gate1643(.O (g2691), .I (g2317));
INVX1 gate1644(.O (g4011), .I (g3486));
INVX1 gate1645(.O (I6798), .I (g5042));
INVX1 gate1646(.O (g4856), .I (I6576));
INVX1 gate1647(.O (g5741), .I (g5602));
INVX1 gate1648(.O (I2802), .I (g1204));
INVX1 gate1649(.O (I3074), .I (g1426));
INVX1 gate1650(.O (I3474), .I (g1450));
INVX1 gate1651(.O (I5753), .I (g4022));
INVX1 gate1652(.O (g5638), .I (I7397));
INVX1 gate1653(.O (g6160), .I (g5926));
INVX1 gate1654(.O (g3226), .I (I4477));
INVX1 gate1655(.O (I5508), .I (g3867));
INVX1 gate1656(.O (g6360), .I (I8144));
INVX1 gate1657(.O (g6933), .I (I9220));
INVX1 gate1658(.O (I5944), .I (g4356));
INVX1 gate1659(.O (g2962), .I (g2008));
INVX1 gate1660(.O (g6521), .I (I8479));
INVX1 gate1661(.O (I9098), .I (g6864));
INVX1 gate1662(.O (g2158), .I (I3281));
INVX1 gate1663(.O (I5472), .I (g3846));
INVX1 gate1664(.O (I8981), .I (g6793));
INVX1 gate1665(.O (g2506), .I (I3632));
INVX1 gate1666(.O (I3080), .I (g1519));
INVX1 gate1667(.O (I8674), .I (g6521));
INVX1 gate1668(.O (g1820), .I (I2880));
INVX1 gate1669(.O (I5043), .I (g3247));
INVX1 gate1670(.O (I6495), .I (g4607));
INVX1 gate1671(.O (g1936), .I (g1756));
INVX1 gate1672(.O (I6437), .I (g4501));
INVX1 gate1673(.O (g3173), .I (I4410));
INVX1 gate1674(.O (I6102), .I (g4399));
INVX1 gate1675(.O (I6302), .I (g4440));
INVX1 gate1676(.O (I8997), .I (g6790));
INVX1 gate1677(.O (g1117), .I (g32));
INVX1 gate1678(.O (I8541), .I (g6452));
INVX1 gate1679(.O (g1317), .I (I2306));
INVX1 gate1680(.O (g3491), .I (g2608));
INVX1 gate1681(.O (g2587), .I (I3714));
INVX1 gate1682(.O (I6579), .I (g4798));
INVX1 gate1683(.O (I5116), .I (g3259));
INVX1 gate1684(.O (I7852), .I (g5993));
INVX1 gate1685(.O (I5316), .I (g3557));
INVX1 gate1686(.O (g6724), .I (I8866));
INVX1 gate1687(.O (I3569), .I (g1789));
INVX1 gate1688(.O (g2111), .I (g1384));
INVX1 gate1689(.O (g2275), .I (I3422));
INVX1 gate1690(.O (g5466), .I (I7146));
INVX1 gate1691(.O (I8332), .I (g6306));
INVX1 gate1692(.O (g4713), .I (I6321));
INVX1 gate1693(.O (I7701), .I (g5720));
INVX1 gate1694(.O (g3369), .I (I4646));
INVX1 gate1695(.O (I8153), .I (g6185));
INVX1 gate1696(.O (g3007), .I (g2197));
INVX1 gate1697(.O (g2615), .I (I3755));
INVX1 gate1698(.O (g6878), .I (I9101));
INVX1 gate1699(.O (I2864), .I (key_out_125));
INVX1 gate1700(.O (g4569), .I (I6143));
INVX1 gate1701(.O (g5571), .I (g5395));
INVX1 gate1702(.O (g5861), .I (g5636));
INVX1 gate1703(.O (g3868), .I (key_out_10));
INVX1 gate1704(.O (g2174), .I (I3313));
INVX1 gate1705(.O (g3459), .I (g2664));
INVX1 gate1706(.O (g815), .I (I1877));
INVX1 gate1707(.O (g1775), .I (g952));
INVX1 gate1708(.O (g5448), .I (g5278));
INVX1 gate1709(.O (g1922), .I (I3025));
INVX1 gate1710(.O (g835), .I (g345));
INVX1 gate1711(.O (g5711), .I (I7472));
INVX1 gate1712(.O (g6835), .I (I9028));
INVX1 gate1713(.O (g1581), .I (g910));
INVX1 gate1714(.O (g6882), .I (I9113));
INVX1 gate1715(.O (I6042), .I (g4374));
INVX1 gate1716(.O (g1060), .I (g107));
INVX1 gate1717(.O (g2284), .I (I3431));
INVX1 gate1718(.O (I6786), .I (g4824));
INVX1 gate1719(.O (g1460), .I (I2457));
INVX1 gate1720(.O (g5774), .I (I7517));
INVX1 gate1721(.O (g4857), .I (I6579));
INVX1 gate1722(.O (g3793), .I (key_out_10));
INVX1 gate1723(.O (g6611), .I (I8699));
INVX1 gate1724(.O (g2591), .I (I3720));
INVX1 gate1725(.O (g3015), .I (I4220));
INVX1 gate1726(.O (g3227), .I (I4480));
INVX1 gate1727(.O (g1739), .I (I2749));
INVX1 gate1728(.O (I6054), .I (g4194));
INVX1 gate1729(.O (g5538), .I (g5331));
INVX1 gate1730(.O (I6296), .I (g4436));
INVX1 gate1731(.O (I4646), .I (g2602));
INVX1 gate1732(.O (I2623), .I (key_out_126));
INVX1 gate1733(.O (g4126), .I (I5460));
INVX1 gate1734(.O (g5509), .I (I7251));
INVX1 gate1735(.O (g4400), .I (I5899));
INVX1 gate1736(.O (g1937), .I (I3044));
INVX1 gate1737(.O (g6541), .I (I8535));
INVX1 gate1738(.O (I9185), .I (g6877));
INVX1 gate1739(.O (I2476), .I (g971));
INVX1 gate1740(.O (I7336), .I (g5534));
INVX1 gate1741(.O (I8600), .I (g6451));
INVX1 gate1742(.O (g2931), .I (g1988));
INVX1 gate1743(.O (g4760), .I (I6386));
INVX1 gate1744(.O (g1294), .I (I2287));
INVX1 gate1745(.O (I1877), .I (g283));
INVX1 gate1746(.O (g6332), .I (I8074));
INVX1 gate1747(.O (g5067), .I (g4801));
INVX1 gate1748(.O (g1190), .I (I2199));
INVX1 gate1749(.O (I2175), .I (g25));
INVX1 gate1750(.O (g6353), .I (I8113));
INVX1 gate1751(.O (g5994), .I (g5873));
INVX1 gate1752(.O (I3608), .I (g1461));
INVX1 gate1753(.O (g2905), .I (g1994));
INVX1 gate1754(.O (I6012), .I (g4167));
INVX1 gate1755(.O (g6744), .I (I8910));
INVX1 gate1756(.O (I3779), .I (g2125));
INVX1 gate1757(.O (g6802), .I (I8972));
INVX1 gate1758(.O (g2628), .I (I3770));
INVX1 gate1759(.O (g1156), .I (I2175));
INVX1 gate1760(.O (g2515), .I (I3641));
INVX1 gate1761(.O (g5493), .I (I7197));
INVX1 gate1762(.O (I7065), .I (g5281));
INVX1 gate1763(.O (g5256), .I (g5077));
INVX1 gate1764(.O (I6706), .I (g4731));
INVX1 gate1765(.O (g4220), .I (I5644));
INVX1 gate1766(.O (g3940), .I (I5177));
INVX1 gate1767(.O (I6371), .I (g4569));
INVX1 gate1768(.O (I4276), .I (g2170));
INVX1 gate1769(.O (g4423), .I (I5920));
INVX1 gate1770(.O (I3161), .I (g1270));
INVX1 gate1771(.O (I3361), .I (g1331));
INVX1 gate1772(.O (g5381), .I (I7039));
INVX1 gate1773(.O (g3388), .I (I4667));
INVX1 gate1774(.O (I9131), .I (g6855));
INVX1 gate1775(.O (I6956), .I (g5124));
INVX1 gate1776(.O (g6901), .I (I9170));
INVX1 gate1777(.O (I5460), .I (g3771));
INVX1 gate1778(.O (I5597), .I (g3821));
INVX1 gate1779(.O (I8623), .I (g6542));
INVX1 gate1780(.O (g3216), .I (I4459));
INVX1 gate1781(.O (I3665), .I (g1824));
INVX1 gate1782(.O (g5685), .I (g5552));
INVX1 gate1783(.O (g6511), .I (I8453));
INVX1 gate1784(.O (I8476), .I (g6457));
INVX1 gate1785(.O (I2424), .I (g719));
INVX1 gate1786(.O (g743), .I (I1844));
INVX1 gate1787(.O (g862), .I (g319));
INVX1 gate1788(.O (g2973), .I (I4170));
INVX1 gate1789(.O (g1954), .I (I3065));
INVX1 gate1790(.O (g3030), .I (I4243));
INVX1 gate1791(.O (g1250), .I (g123));
INVX1 gate1792(.O (I5739), .I (g3942));
INVX1 gate1793(.O (g1363), .I (I2399));
INVX1 gate1794(.O (I4986), .I (g3638));
INVX1 gate1795(.O (I3999), .I (g1837));
INVX1 gate1796(.O (g3247), .I (g2973));
INVX1 gate1797(.O (g4127), .I (I5463));
INVX1 gate1798(.O (I3346), .I (g1327));
INVX1 gate1799(.O (g5950), .I (g5730));
INVX1 gate1800(.O (g1053), .I (g197));
INVX1 gate1801(.O (g2040), .I (g1738));
INVX1 gate1802(.O (g6600), .I (I8668));
INVX1 gate1803(.O (g6574), .I (g6484));
INVX1 gate1804(.O (I2231), .I (g465));
INVX1 gate1805(.O (I1844), .I (g208));
INVX1 gate1806(.O (g2440), .I (I3575));
INVX1 gate1807(.O (g3564), .I (g2618));
INVX1 gate1808(.O (g6714), .I (g6670));
INVX1 gate1809(.O (I2643), .I (g965));
INVX1 gate1810(.O (g4146), .I (I5520));
INVX1 gate1811(.O (I5668), .I (g3828));
INVX1 gate1812(.O (g4633), .I (g4284));
INVX1 gate1813(.O (I8285), .I (g6310));
INVX1 gate1814(.O (I5840), .I (g3732));
INVX1 gate1815(.O (I8500), .I (g6431));
INVX1 gate1816(.O (g791), .I (I1865));
INVX1 gate1817(.O (g4103), .I (I5391));
INVX1 gate1818(.O (g6580), .I (g6491));
INVX1 gate1819(.O (I7859), .I (g6032));
INVX1 gate1820(.O (g5631), .I (g5536));
INVX1 gate1821(.O (g3638), .I (g3108));
INVX1 gate1822(.O (g5723), .I (I7484));
INVX1 gate1823(.O (I9173), .I (g6876));
INVX1 gate1824(.O (I3240), .I (g1460));
INVX1 gate1825(.O (g4732), .I (I6362));
INVX1 gate1826(.O (g3108), .I (I4354));
INVX1 gate1827(.O (g3308), .I (g3060));
INVX1 gate1828(.O (I6759), .I (g4778));
INVX1 gate1829(.O (g2875), .I (g1940));
INVX1 gate1830(.O (g4753), .I (I6377));
INVX1 gate1831(.O (g4508), .I (I6036));
INVX1 gate1832(.O (g917), .I (I1942));
INVX1 gate1833(.O (I8809), .I (g6687));
INVX1 gate1834(.O (I7342), .I (g5579));
INVX1 gate1835(.O (g6623), .I (I8727));
INVX1 gate1836(.O (g6076), .I (g5797));
INVX1 gate1837(.O (I7081), .I (g5281));
INVX1 gate1838(.O (g6889), .I (I9134));
INVX1 gate1839(.O (g5751), .I (I7506));
INVX1 gate1840(.O (I3316), .I (g1344));
INVX1 gate1841(.O (g3589), .I (g3094));
INVX1 gate1842(.O (I7481), .I (g5629));
INVX1 gate1843(.O (I3034), .I (g1519));
INVX1 gate1844(.O (g3466), .I (I4706));
INVX1 gate1845(.O (g2410), .I (I3550));
INVX1 gate1846(.O (I7692), .I (g5711));
INVX1 gate1847(.O (I3434), .I (g1627));
INVX1 gate1848(.O (I4516), .I (g2777));
INVX1 gate1849(.O (I7497), .I (g5687));
INVX1 gate1850(.O (g4116), .I (I5430));
INVX1 gate1851(.O (g6375), .I (I8189));
INVX1 gate1852(.O (g2884), .I (g1957));
INVX1 gate1853(.O (I2044), .I (g681));
INVX1 gate1854(.O (g3571), .I (g3084));
INVX1 gate1855(.O (g2839), .I (g2535));
INVX1 gate1856(.O (g3861), .I (I5084));
INVX1 gate1857(.O (g6722), .I (I8860));
INVX1 gate1858(.O (g4034), .I (I5333));
INVX1 gate1859(.O (I7960), .I (g5925));
INVX1 gate1860(.O (g852), .I (g634));
INVX1 gate1861(.O (I2269), .I (g899));
INVX1 gate1862(.O (g6651), .I (I8749));
INVX1 gate1863(.O (g3448), .I (I4684));
INVX1 gate1864(.O (g4565), .I (g4195));
INVX1 gate1865(.O (I3681), .I (g1821));
INVX1 gate1866(.O (I5053), .I (g3710));
INVX1 gate1867(.O (g3455), .I (g2637));
INVX1 gate1868(.O (g6285), .I (I8005));
INVX1 gate1869(.O (g4147), .I (I5523));
INVX1 gate1870(.O (g6500), .I (I8420));
INVX1 gate1871(.O (g2172), .I (I3307));
INVX1 gate1872(.O (I2712), .I (g1203));
INVX1 gate1873(.O (I9227), .I (g6937));
INVX1 gate1874(.O (I5568), .I (g3897));
INVX1 gate1875(.O (g4533), .I (I6111));
INVX1 gate1876(.O (g3846), .I (I5053));
INVX1 gate1877(.O (g2618), .I (I3758));
INVX1 gate1878(.O (I3596), .I (g1305));
INVX1 gate1879(.O (g2667), .I (I3811));
INVX1 gate1880(.O (g1683), .I (g1017));
INVX1 gate1881(.O (g2343), .I (I3493));
INVX1 gate1882(.O (g5168), .I (g5099));
INVX1 gate1883(.O (I3013), .I (g1519));
INVX1 gate1884(.O (g6339), .I (I8093));
INVX1 gate1885(.O (g3196), .I (I4433));
INVX1 gate1886(.O (g4914), .I (g4816));
INVX1 gate1887(.O (g3803), .I (I5002));
INVX1 gate1888(.O (g4210), .I (I5630));
INVX1 gate1889(.O (I7267), .I (g5458));
INVX1 gate1890(.O (g1894), .I (I2989));
INVX1 gate1891(.O (I5157), .I (g3454));
INVX1 gate1892(.O (g6838), .I (I9035));
INVX1 gate1893(.O (I9203), .I (g6921));
INVX1 gate1894(.O (I2961), .I (g1731));
INVX1 gate1895(.O (g6424), .I (I8282));
INVX1 gate1896(.O (g2134), .I (I3258));
INVX1 gate1897(.O (I6362), .I (g4569));
INVX1 gate1898(.O (g1735), .I (I2745));
INVX1 gate1899(.O (I8273), .I (g6301));
INVX1 gate1900(.O (g6809), .I (I8981));
INVX1 gate1901(.O (g5890), .I (g5753));
INVX1 gate1902(.O (g1782), .I (I2828));
INVX1 gate1903(.O (I4340), .I (g1935));
INVX1 gate1904(.O (I6452), .I (g4629));
INVX1 gate1905(.O (I5929), .I (g4152));
INVX1 gate1906(.O (g1661), .I (g1076));
INVX1 gate1907(.O (I8044), .I (g6252));
INVX1 gate1908(.O (g2555), .I (I3672));
INVX1 gate1909(.O (g6231), .I (g6044));
INVX1 gate1910(.O (g5011), .I (I6649));
INVX1 gate1911(.O (I8444), .I (g6421));
INVX1 gate1912(.O (g3067), .I (I4294));
INVX1 gate1913(.O (I2414), .I (g784));
INVX1 gate1914(.O (g729), .I (I1838));
INVX1 gate1915(.O (g5411), .I (I7077));
INVX1 gate1916(.O (g6523), .I (I8485));
INVX1 gate1917(.O (g861), .I (g179));
INVX1 gate1918(.O (I2946), .I (g1587));
INVX1 gate1919(.O (g2792), .I (g2416));
INVX1 gate1920(.O (g1627), .I (I2584));
INVX1 gate1921(.O (g4117), .I (I5433));
INVX1 gate1922(.O (g1292), .I (I2281));
INVX1 gate1923(.O (I5626), .I (g3914));
INVX1 gate1924(.O (g3093), .I (I4334));
INVX1 gate1925(.O (g898), .I (g47));
INVX1 gate1926(.O (g1998), .I (I3109));
INVX1 gate1927(.O (g1646), .I (I2617));
INVX1 gate1928(.O (g5992), .I (g5869));
INVX1 gate1929(.O (g4601), .I (g4191));
INVX1 gate1930(.O (g1084), .I (g98));
INVX1 gate1931(.O (g6104), .I (I7808));
INVX1 gate1932(.O (g854), .I (g646));
INVX1 gate1933(.O (g1039), .I (g662));
INVX1 gate1934(.O (g1484), .I (I2473));
INVX1 gate1935(.O (I3581), .I (g1491));
INVX1 gate1936(.O (g6499), .I (I8417));
INVX1 gate1937(.O (g1439), .I (I2449));
INVX1 gate1938(.O (I9028), .I (g6806));
INVX1 gate1939(.O (I8961), .I (g6778));
INVX1 gate1940(.O (g4775), .I (I6425));
INVX1 gate1941(.O (I6470), .I (g4473));
INVX1 gate1942(.O (g5573), .I (g5403));
INVX1 gate1943(.O (g3847), .I (I5056));
INVX1 gate1944(.O (g5480), .I (I7176));
INVX1 gate1945(.O (I6425), .I (g4619));
INVX1 gate1946(.O (I2831), .I (key_out_128));
INVX1 gate1947(.O (g2494), .I (I3623));
INVX1 gate1948(.O (I2182), .I (g692));
INVX1 gate1949(.O (g2518), .I (I3644));
INVX1 gate1950(.O (g1583), .I (g1001));
INVX1 gate1951(.O (g1702), .I (g1107));
INVX1 gate1952(.O (I2382), .I (g719));
INVX1 gate1953(.O (I8414), .I (g6418));
INVX1 gate1954(.O (g3263), .I (g3015));
INVX1 gate1955(.O (I8946), .I (g6778));
INVX1 gate1956(.O (g1919), .I (I3022));
INVX1 gate1957(.O (I2805), .I (g1205));
INVX1 gate1958(.O (I2916), .I (g1643));
INVX1 gate1959(.O (g2776), .I (g2378));
INVX1 gate1960(.O (I2749), .I (key_out_128));
INVX1 gate1961(.O (g4784), .I (I6444));
INVX1 gate1962(.O (g6044), .I (g5824));
INVX1 gate1963(.O (g1276), .I (g847));
INVX1 gate1964(.O (I4402), .I (g2283));
INVX1 gate1965(.O (I3294), .I (g1720));
INVX1 gate1966(.O (I3840), .I (g2125));
INVX1 gate1967(.O (I6406), .I (g4473));
INVX1 gate1968(.O (I5475), .I (g3852));
INVX1 gate1969(.O (g6572), .I (I8600));
INVX1 gate1970(.O (I4762), .I (g2862));
INVX1 gate1971(.O (I7349), .I (g5532));
INVX1 gate1972(.O (I6635), .I (g4745));
INVX1 gate1973(.O (g2264), .I (I3405));
INVX1 gate1974(.O (g6712), .I (g6676));
INVX1 gate1975(.O (g851), .I (g606));
INVX1 gate1976(.O (I6766), .I (g4783));
INVX1 gate1977(.O (I6087), .I (g4392));
INVX1 gate1978(.O (I6105), .I (g4400));
INVX1 gate1979(.O (g6543), .I (I8541));
INVX1 gate1980(.O (g4840), .I (I6528));
INVX1 gate1981(.O (I6305), .I (g4441));
INVX1 gate1982(.O (I6801), .I (g5045));
INVX1 gate1983(.O (g2360), .I (g1793));
INVX1 gate1984(.O (g2933), .I (I4123));
INVX1 gate1985(.O (g3723), .I (I4903));
INVX1 gate1986(.O (g1647), .I (I2620));
INVX1 gate1987(.O (g4190), .I (I5600));
INVX1 gate1988(.O (I5526), .I (g3848));
INVX1 gate1989(.O (I5998), .I (g4157));
INVX1 gate1990(.O (I8335), .I (g6308));
INVX1 gate1991(.O (I8831), .I (g6665));
INVX1 gate1992(.O (I9217), .I (g6931));
INVX1 gate1993(.O (g1546), .I (g1101));
INVX1 gate1994(.O (I2873), .I (key_out_126));
INVX1 gate1995(.O (I2037), .I (g679));
INVX1 gate1996(.O (g6534), .I (I8518));
INVX1 gate1997(.O (g6729), .I (I8881));
INVX1 gate1998(.O (g3605), .I (I4802));
INVX1 gate1999(.O (I5084), .I (key_out_6));
INVX1 gate2000(.O (I5603), .I (g3893));
INVX1 gate2001(.O (g2996), .I (I4189));
INVX1 gate2002(.O (I2653), .I (g996));
INVX1 gate2003(.O (I5484), .I (g3875));
INVX1 gate2004(.O (I3942), .I (g1833));
INVX1 gate2005(.O (g1503), .I (g878));
INVX1 gate2006(.O (I5439), .I (g3730));
INVX1 gate2007(.O (I8916), .I (g6742));
INVX1 gate2008(.O (g1925), .I (I3028));
INVX1 gate2009(.O (I8749), .I (g6560));
INVX1 gate2010(.O (g2179), .I (I3328));
INVX1 gate2011(.O (g6014), .I (g5824));
INVX1 gate2012(.O (g6885), .I (I9122));
INVX1 gate2013(.O (I6045), .I (g4375));
INVX1 gate2014(.O (g4704), .I (I6302));
INVX1 gate2015(.O (g6414), .I (I8252));
INVX1 gate2016(.O (I5702), .I (g3845));
INVX1 gate2017(.O (g1320), .I (I2315));
INVX1 gate2018(.O (g3041), .I (I4258));
INVX1 gate2019(.O (g5383), .I (I7045));
INVX1 gate2020(.O (g5924), .I (I7704));
INVX1 gate2021(.O (g5220), .I (g4903));
INVX1 gate2022(.O (I7119), .I (g5303));
INVX1 gate2023(.O (g6903), .I (I9176));
INVX1 gate2024(.O (g2777), .I (I3965));
INVX1 gate2025(.O (g3441), .I (I4681));
INVX1 gate2026(.O (g2835), .I (g2506));
INVX1 gate2027(.O (I3053), .I (g1407));
INVX1 gate2028(.O (I1958), .I (key_out_40));
INVX1 gate2029(.O (g4250), .I (I5702));
INVX1 gate2030(.O (g6513), .I (I8459));
INVX1 gate2031(.O (g913), .I (g658));
INVX1 gate2032(.O (I6283), .I (g4613));
INVX1 gate2033(.O (I7258), .I (g5458));
INVX1 gate2034(.O (I5952), .I (g4367));
INVX1 gate2035(.O (g4810), .I (I6488));
INVX1 gate2036(.O (g2882), .I (g1854));
INVX1 gate2037(.O (I7352), .I (g5533));
INVX1 gate2038(.O (g3673), .I (g3075));
INVX1 gate2039(.O (I2442), .I (g872));
INVX1 gate2040(.O (g1789), .I (I2839));
INVX1 gate2041(.O (g6036), .I (g5824));
INVX1 gate2042(.O (I8632), .I (g6548));
INVX1 gate2043(.O (I2364), .I (key_out_123));
INVX1 gate2044(.O (g980), .I (I2037));
INVX1 gate2045(.O (I8653), .I (g6531));
INVX1 gate2046(.O (g1771), .I (I2808));
INVX1 gate2047(.O (g3772), .I (g3466));
INVX1 gate2048(.O (I6582), .I (g4765));
INVX1 gate2049(.O (g5051), .I (I6689));
INVX1 gate2050(.O (g2981), .I (g2179));
INVX1 gate2051(.O (I8579), .I (g6438));
INVX1 gate2052(.O (I8869), .I (g6694));
INVX1 gate2053(.O (I4489), .I (g2975));
INVX1 gate2054(.O (g3458), .I (g2656));
INVX1 gate2055(.O (g865), .I (g188));
INVX1 gate2056(.O (I2296), .I (g893));
INVX1 gate2057(.O (g3890), .I (g3575));
INVX1 gate2058(.O (g2997), .I (I4192));
INVX1 gate2059(.O (I6015), .I (g4170));
INVX1 gate2060(.O (g2541), .I (I3659));
INVX1 gate2061(.O (I8752), .I (g6514));
INVX1 gate2062(.O (I4471), .I (g3040));
INVX1 gate2063(.O (I7170), .I (g5435));
INVX1 gate2064(.O (g6422), .I (I8276));
INVX1 gate2065(.O (g2353), .I (I3505));
INVX1 gate2066(.O (g4929), .I (I6621));
INVX1 gate2067(.O (I4955), .I (key_out_11));
INVX1 gate2068(.O (I3626), .I (g1684));
INVX1 gate2069(.O (g2744), .I (g2336));
INVX1 gate2070(.O (g909), .I (I1935));
INVX1 gate2071(.O (g1738), .I (g1108));
INVX1 gate2072(.O (g2802), .I (g2437));
INVX1 gate2073(.O (g3074), .I (I4303));
INVX1 gate2074(.O (g949), .I (g79));
INVX1 gate2075(.O (g1991), .I (I3102));
INVX1 gate2076(.O (g6560), .I (I8564));
INVX1 gate2077(.O (I5320), .I (key_out_9));
INVX1 gate2078(.O (g4626), .I (g4270));
INVX1 gate2079(.O (g1340), .I (I2373));
INVX1 gate2080(.O (I2029), .I (g677));
INVX1 gate2081(.O (I9021), .I (g6812));
INVX1 gate2082(.O (g3480), .I (g2986));
INVX1 gate2083(.O (g1690), .I (I2692));
INVX1 gate2084(.O (g6653), .I (I8755));
INVX1 gate2085(.O (g6102), .I (I7802));
INVX1 gate2086(.O (I2281), .I (g900));
INVX1 gate2087(.O (I7061), .I (g5281));
INVX1 gate2088(.O (I7187), .I (g5387));
INVX1 gate2089(.O (g6579), .I (g6490));
INVX1 gate2090(.O (g5116), .I (g4810));
INVX1 gate2091(.O (I5987), .I (g4224));
INVX1 gate2092(.O (g5316), .I (I6976));
INVX1 gate2093(.O (g1656), .I (I2635));
INVX1 gate2094(.O (I6689), .I (g4758));
INVX1 gate2095(.O (g5434), .I (I7110));
INVX1 gate2096(.O (g2574), .I (I3681));
INVX1 gate2097(.O (g2864), .I (g1887));
INVX1 gate2098(.O (g4778), .I (I6430));
INVX1 gate2099(.O (g855), .I (g650));
INVX1 gate2100(.O (g5147), .I (I6809));
INVX1 gate2101(.O (I3782), .I (g2145));
INVX1 gate2102(.O (g4894), .I (g4813));
INVX1 gate2103(.O (I2745), .I (g1249));
INVX1 gate2104(.O (I8189), .I (g6179));
INVX1 gate2105(.O (I4229), .I (g2284));
INVX1 gate2106(.O (I6430), .I (g4620));
INVX1 gate2107(.O (g3976), .I (I5252));
INVX1 gate2108(.O (I2791), .I (key_out_120));
INVX1 gate2109(.O (I6247), .I (g4609));
INVX1 gate2110(.O (I7514), .I (g5590));
INVX1 gate2111(.O (I2309), .I (key_out_120));
INVX1 gate2112(.O (I9101), .I (g6855));
INVX1 gate2113(.O (g1110), .I (I2140));
INVX1 gate2114(.O (I8888), .I (g6708));
INVX1 gate2115(.O (g2580), .I (I3691));
INVX1 gate2116(.O (g5210), .I (I6874));
INVX1 gate2117(.O (g6786), .I (I8946));
INVX1 gate2118(.O (I6564), .I (g4712));
INVX1 gate2119(.O (I8171), .I (g6170));
INVX1 gate2120(.O (I2808), .I (key_out_126));
INVX1 gate2121(.O (I8429), .I (g6425));
INVX1 gate2122(.O (g5596), .I (I7358));
INVX1 gate2123(.O (g6164), .I (g5926));
INVX1 gate2124(.O (g6364), .I (I8156));
INVX1 gate2125(.O (g6233), .I (g6052));
INVX1 gate2126(.O (I5991), .I (g4226));
INVX1 gate2127(.O (I2707), .I (g1190));
INVX1 gate2128(.O (g4292), .I (g4059));
INVX1 gate2129(.O (I7695), .I (g5714));
INVX1 gate2130(.O (I7637), .I (g5751));
INVX1 gate2131(.O (g2968), .I (g2179));
INVX1 gate2132(.O (I5078), .I (g3719));
INVX1 gate2133(.O (g1824), .I (I2890));
INVX1 gate2134(.O (g4526), .I (I6090));
INVX1 gate2135(.O (I5478), .I (g3859));
INVX1 gate2136(.O (g1236), .I (I2234));
INVX1 gate2137(.O (I7107), .I (g5277));
INVX1 gate2138(.O (I5907), .I (g3883));
INVX1 gate2139(.O (g6725), .I (I8869));
INVX1 gate2140(.O (g1762), .I (I2791));
INVX1 gate2141(.O (g2889), .I (g1975));
INVX1 gate2142(.O (I6108), .I (g4403));
INVX1 gate2143(.O (g4603), .I (I6170));
INVX1 gate2144(.O (g6532), .I (I8512));
INVX1 gate2145(.O (I6308), .I (g4443));
INVX1 gate2146(.O (I5517), .I (g3885));
INVX1 gate2147(.O (I9041), .I (g6835));
INVX1 gate2148(.O (I2449), .I (g971));
INVX1 gate2149(.O (g4439), .I (I5952));
INVX1 gate2150(.O (g5117), .I (I6763));
INVX1 gate2151(.O (g6553), .I (I8555));
INVX1 gate2152(.O (g4850), .I (I6558));
INVX1 gate2153(.O (I8684), .I (g6567));
INVX1 gate2154(.O (I5876), .I (g3870));
INVX1 gate2155(.O (I8745), .I (g6513));
INVX1 gate2156(.O (g2175), .I (I3316));
INVX1 gate2157(.O (g2871), .I (g1919));
INVX1 gate2158(.O (I2604), .I (key_out_124));
INVX1 gate2159(.O (g3183), .I (I4420));
INVX1 gate2160(.O (g2722), .I (I3883));
INVX1 gate2161(.O (I4462), .I (g2135));
INVX1 gate2162(.O (I8309), .I (g6304));
INVX1 gate2163(.O (g1556), .I (g878));
INVX1 gate2164(.O (I6066), .I (g4382));
INVX1 gate2165(.O (g3779), .I (g3466));
INVX1 gate2166(.O (g1222), .I (I2225));
INVX1 gate2167(.O (g4702), .I (I6296));
INVX1 gate2168(.O (g6412), .I (I8246));
INVX1 gate2169(.O (g896), .I (g22));
INVX1 gate2170(.O (g3023), .I (g2215));
INVX1 gate2171(.O (I7251), .I (g5458));
INVX1 gate2172(.O (g1928), .I (I3031));
INVX1 gate2173(.O (I7811), .I (g5921));
INVX1 gate2174(.O (g6706), .I (I8828));
INVX1 gate2175(.O (g5922), .I (I7698));
INVX1 gate2176(.O (I8707), .I (g6520));
INVX1 gate2177(.O (g1064), .I (g102));
INVX1 gate2178(.O (I2584), .I (key_out_31));
INVX1 gate2179(.O (I5214), .I (key_out_7));
INVX1 gate2180(.O (g6888), .I (I9131));
INVX1 gate2181(.O (g1899), .I (I2998));
INVX1 gate2182(.O (I6048), .I (g4376));
INVX1 gate2183(.O (g5581), .I (I7339));
INVX1 gate2184(.O (I6448), .I (g4626));
INVX1 gate2185(.O (g6371), .I (I8177));
INVX1 gate2186(.O (g4276), .I (I5731));
INVX1 gate2187(.O (I4249), .I (g2525));
INVX1 gate2188(.O (g5597), .I (I7361));
INVX1 gate2189(.O (I3004), .I (g1426));
INVX1 gate2190(.O (I1825), .I (g361));
INVX1 gate2191(.O (g4561), .I (g4189));
INVX1 gate2192(.O (g2838), .I (g2515));
INVX1 gate2193(.O (I3647), .I (g1747));
INVX1 gate2194(.O (g3451), .I (g2615));
INVX1 gate2195(.O (I2162), .I (g197));
INVX1 gate2196(.O (g1563), .I (g1006));
INVX1 gate2197(.O (I9011), .I (g6819));
INVX1 gate2198(.O (I4192), .I (g1847));
INVX1 gate2199(.O (g2809), .I (I4019));
INVX1 gate2200(.O (I3764), .I (g2044));
INVX1 gate2201(.O (g5784), .I (I7583));
INVX1 gate2202(.O (I3546), .I (g1586));
INVX1 gate2203(.O (I5002), .I (g3612));
INVX1 gate2204(.O (g4527), .I (I6093));
INVX1 gate2205(.O (g4404), .I (I5907));
INVX1 gate2206(.O (g1295), .I (I2290));
INVX1 gate2207(.O (g4647), .I (g4296));
INVX1 gate2208(.O (g3346), .I (I4623));
INVX1 gate2209(.O (I5236), .I (g3545));
INVX1 gate2210(.O (g2672), .I (I3816));
INVX1 gate2211(.O (g2231), .I (I3358));
INVX1 gate2212(.O (g4764), .I (I6400));
INVX1 gate2213(.O (g5995), .I (g5824));
INVX1 gate2214(.O (I9074), .I (g6844));
INVX1 gate2215(.O (g5479), .I (I7173));
INVX1 gate2216(.O (g2643), .I (I3785));
INVX1 gate2217(.O (I6780), .I (g4825));
INVX1 gate2218(.O (g6745), .I (I8913));
INVX1 gate2219(.O (g1394), .I (g1206));
INVX1 gate2220(.O (g4503), .I (I6023));
INVX1 gate2221(.O (I7612), .I (g5605));
INVX1 gate2222(.O (g1731), .I (I2735));
INVX1 gate2223(.O (I2728), .I (g1232));
INVX1 gate2224(.O (g1557), .I (g1017));
INVX1 gate2225(.O (g2634), .I (I3776));
INVX1 gate2226(.O (g1966), .I (I3077));
INVX1 gate2227(.O (g4224), .I (g4046));
INVX1 gate2228(.O (I5556), .I (g4059));
INVX1 gate2229(.O (I2185), .I (g29));
INVX1 gate2230(.O (g2104), .I (g1372));
INVX1 gate2231(.O (g2099), .I (g1366));
INVX1 gate2232(.O (g3240), .I (I4519));
INVX1 gate2233(.O (I2385), .I (g784));
INVX1 gate2234(.O (g6707), .I (I8831));
INVX1 gate2235(.O (g1471), .I (I2464));
INVX1 gate2236(.O (g4120), .I (I5442));
INVX1 gate2237(.O (I4031), .I (g1846));
INVX1 gate2238(.O (g4320), .I (g4011));
INVX1 gate2239(.O (I4252), .I (g2555));
INVX1 gate2240(.O (I3617), .I (g1305));
INVX1 gate2241(.O (I3906), .I (g2234));
INVX1 gate2242(.O (I6093), .I (g4394));
INVX1 gate2243(.O (I8162), .I (g6189));
INVX1 gate2244(.O (g3043), .I (I4264));
INVX1 gate2245(.O (g971), .I (g658));
INVX1 gate2246(.O (I5899), .I (g3748));
INVX1 gate2247(.O (I4176), .I (g2268));
INVX1 gate2248(.O (I6816), .I (g5111));
INVX1 gate2249(.O (I3516), .I (g1295));
INVX1 gate2250(.O (g2754), .I (g2347));
INVX1 gate2251(.O (g4617), .I (g4242));
INVX1 gate2252(.O (g3034), .I (I4249));
INVX1 gate2253(.O (g1254), .I (g152));
INVX1 gate2254(.O (g1814), .I (I2873));
INVX1 gate2255(.O (g6575), .I (g6486));
INVX1 gate2256(.O (g4516), .I (I6060));
INVX1 gate2257(.O (g6715), .I (g6673));
INVX1 gate2258(.O (g4771), .I (I6417));
INVX1 gate2259(.O (g2044), .I (I3161));
INVX1 gate2260(.O (I6685), .I (g4716));
INVX1 gate2261(.O (g5250), .I (g4929));
INVX1 gate2262(.O (g6604), .I (I8678));
INVX1 gate2263(.O (g1038), .I (g127));
INVX1 gate2264(.O (I6397), .I (g4473));
INVX1 gate2265(.O (g6498), .I (I8414));
INVX1 gate2266(.O (g1773), .I (I2814));
INVX1 gate2267(.O (I2131), .I (g24));
INVX1 gate2268(.O (g5432), .I (I7104));
INVX1 gate2269(.O (g4299), .I (I5756));
INVX1 gate2270(.O (g6833), .I (I9024));
INVX1 gate2271(.O (I8730), .I (g6535));
INVX1 gate2272(.O (g5453), .I (g5296));
INVX1 gate2273(.O (I4270), .I (g2555));
INVX1 gate2274(.O (g2862), .I (I4066));
INVX1 gate2275(.O (I2635), .I (g1055));
INVX1 gate2276(.O (g2712), .I (g2320));
INVX1 gate2277(.O (I8881), .I (g6711));
INVX1 gate2278(.O (I5394), .I (g4016));
INVX1 gate2279(.O (g1769), .I (I2802));
INVX1 gate2280(.O (g3914), .I (I5153));
INVX1 gate2281(.O (g6584), .I (I8620));
INVX1 gate2282(.O (I1859), .I (g277));
INVX1 gate2283(.O (g6539), .I (I8531));
INVX1 gate2284(.O (g6896), .I (I9155));
INVX1 gate2285(.O (g1836), .I (I2922));
INVX1 gate2286(.O (g5568), .I (g5423));
INVX1 gate2287(.O (I8070), .I (g6116));
INVX1 gate2288(.O (I5731), .I (g3942));
INVX1 gate2289(.O (I8470), .I (g6461));
INVX1 gate2290(.O (I8897), .I (g6707));
INVX1 gate2291(.O (g1918), .I (I3019));
INVX1 gate2292(.O (I3244), .I (g1772));
INVX1 gate2293(.O (I7490), .I (g5583));
INVX1 gate2294(.O (I4980), .I (key_out_3));
INVX1 gate2295(.O (g5912), .I (g5853));
INVX1 gate2296(.O (I4324), .I (g1918));
INVX1 gate2297(.O (I3140), .I (g1317));
INVX1 gate2298(.O (g2961), .I (g1861));
INVX1 gate2299(.O (I5071), .I (g3263));
INVX1 gate2300(.O (I3340), .I (g1282));
INVX1 gate2301(.O (I5705), .I (g3942));
INVX1 gate2302(.O (g6162), .I (g5926));
INVX1 gate2303(.O (I3478), .I (g1450));
INVX1 gate2304(.O (g6362), .I (I8150));
INVX1 gate2305(.O (g6419), .I (I8267));
INVX1 gate2306(.O (I6723), .I (g4761));
INVX1 gate2307(.O (g4140), .I (I5502));
INVX1 gate2308(.O (g6052), .I (g5824));
INVX1 gate2309(.O (g2927), .I (g1979));
INVX1 gate2310(.O (I5948), .I (g4360));
INVX1 gate2311(.O (I9220), .I (g6930));
INVX1 gate2312(.O (g2885), .I (g1963));
INVX1 gate2313(.O (I7355), .I (g5535));
INVX1 gate2314(.O (I8678), .I (g6565));
INVX1 gate2315(.O (I2445), .I (g971));
INVX1 gate2316(.O (g2660), .I (I3804));
INVX1 gate2317(.O (g2946), .I (g2296));
INVX1 gate2318(.O (g938), .I (g59));
INVX1 gate2319(.O (g4435), .I (I5944));
INVX1 gate2320(.O (I2373), .I (key_out_123));
INVX1 gate2321(.O (g4517), .I (I6063));
INVX1 gate2322(.O (I7698), .I (g5717));
INVX1 gate2323(.O (I3656), .I (g1484));
INVX1 gate2324(.O (g3601), .I (I4794));
INVX1 gate2325(.O (I2491), .I (g821));
INVX1 gate2326(.O (g2903), .I (g1902));
INVX1 gate2327(.O (I8635), .I (g6552));
INVX1 gate2328(.O (g6728), .I (I8878));
INVX1 gate2329(.O (g6486), .I (g6363));
INVX1 gate2330(.O (I2169), .I (g269));
INVX1 gate2331(.O (g942), .I (g69));
INVX1 gate2332(.O (g6730), .I (I8884));
INVX1 gate2333(.O (I9161), .I (g6880));
INVX1 gate2334(.O (g3775), .I (g3388));
INVX1 gate2335(.O (g6504), .I (I8432));
INVX1 gate2336(.O (g3922), .I (I5157));
INVX1 gate2337(.O (I7463), .I (g5622));
INVX1 gate2338(.O (I2578), .I (key_out_128));
INVX1 gate2339(.O (g6385), .I (g6271));
INVX1 gate2340(.O (g6881), .I (I9110));
INVX1 gate2341(.O (I5409), .I (g3980));
INVX1 gate2342(.O (g2036), .I (g1764));
INVX1 gate2343(.O (g706), .I (I1825));
INVX1 gate2344(.O (I6441), .I (g4624));
INVX1 gate2345(.O (g4915), .I (g4669));
INVX1 gate2346(.O (g2178), .I (I3325));
INVX1 gate2347(.O (g2436), .I (I3569));
INVX1 gate2348(.O (g2679), .I (I3823));
INVX1 gate2349(.O (g6070), .I (g5824));
INVX1 gate2350(.O (g2378), .I (I3525));
INVX1 gate2351(.O (g3060), .I (I4285));
INVX1 gate2352(.O (I3310), .I (g1640));
INVX1 gate2353(.O (g6897), .I (I9158));
INVX1 gate2354(.O (g1837), .I (I2925));
INVX1 gate2355(.O (I8755), .I (g6561));
INVX1 gate2356(.O (g3460), .I (g2667));
INVX1 gate2357(.O (I8226), .I (g6328));
INVX1 gate2358(.O (g6425), .I (I8285));
INVX1 gate2359(.O (g2135), .I (I3261));
INVX1 gate2360(.O (I4510), .I (g2753));
INVX1 gate2361(.O (I9146), .I (g6890));
INVX1 gate2362(.O (g4110), .I (I5412));
INVX1 gate2363(.O (I7167), .I (g5434));
INVX1 gate2364(.O (I7318), .I (g5452));
INVX1 gate2365(.O (I4291), .I (g2241));
INVX1 gate2366(.O (g5894), .I (g5731));
INVX1 gate2367(.O (g2805), .I (g2443));
INVX1 gate2368(.O (g910), .I (I1938));
INVX1 gate2369(.O (g1788), .I (g985));
INVX1 gate2370(.O (g2422), .I (I3560));
INVX1 gate2371(.O (I6772), .I (g4788));
INVX1 gate2372(.O (I7193), .I (g5466));
INVX1 gate2373(.O (I8491), .I (g6480));
INVX1 gate2374(.O (g3079), .I (I4312));
INVX1 gate2375(.O (I6531), .I (g4704));
INVX1 gate2376(.O (g4402), .I (g4017));
INVX1 gate2377(.O (g784), .I (I1862));
INVX1 gate2378(.O (g1249), .I (I2240));
INVX1 gate2379(.O (g4824), .I (g4615));
INVX1 gate2380(.O (g837), .I (g353));
INVX1 gate2381(.O (g5661), .I (g5518));
INVX1 gate2382(.O (g3840), .I (I5043));
INVX1 gate2383(.O (g719), .I (I1835));
INVX1 gate2384(.O (I3590), .I (g1781));
INVX1 gate2385(.O (g6406), .I (I8232));
INVX1 gate2386(.O (g5475), .I (I7161));
INVX1 gate2387(.O (I7686), .I (g5705));
INVX1 gate2388(.O (g1842), .I (g1612));
INVX1 gate2389(.O (I2721), .I (g1219));
INVX1 gate2390(.O (g1192), .I (g44));
INVX1 gate2391(.O (I8459), .I (g6427));
INVX1 gate2392(.O (g6105), .I (I7811));
INVX1 gate2393(.O (g6087), .I (g5813));
INVX1 gate2394(.O (g6801), .I (I8969));
INVX1 gate2395(.O (g6305), .I (I8027));
INVX1 gate2396(.O (g5292), .I (I6942));
INVX1 gate2397(.O (I8767), .I (g6619));
INVX1 gate2398(.O (g6487), .I (g6365));
INVX1 gate2399(.O (I3556), .I (g1484));
INVX1 gate2400(.O (g3501), .I (g2650));
INVX1 gate2401(.O (I3222), .I (g1790));
INVX1 gate2402(.O (I8535), .I (g6447));
INVX1 gate2403(.O (g4657), .I (I6244));
INVX1 gate2404(.O (I8582), .I (g6439));
INVX1 gate2405(.O (g1854), .I (I2958));
INVX1 gate2406(.O (I9116), .I (g6864));
INVX1 gate2407(.O (I8261), .I (g6298));
INVX1 gate2408(.O (g5084), .I (g4727));
INVX1 gate2409(.O (g4222), .I (I5654));
INVX1 gate2410(.O (g2437), .I (I3572));
INVX1 gate2411(.O (g2653), .I (I3797));
INVX1 gate2412(.O (I6992), .I (g5151));
INVX1 gate2413(.O (I1932), .I (g667));
INVX1 gate2414(.O (g2102), .I (I3222));
INVX1 gate2415(.O (g5439), .I (g5261));
INVX1 gate2416(.O (I3785), .I (g2346));
INVX1 gate2417(.O (I2940), .I (g1653));
INVX1 gate2418(.O (I5837), .I (g3850));
INVX1 gate2419(.O (g2869), .I (g2433));
INVX1 gate2420(.O (I2388), .I (g878));
INVX1 gate2421(.O (I6573), .I (g4721));
INVX1 gate2422(.O (I3563), .I (g1461));
INVX1 gate2423(.O (g5702), .I (I7463));
INVX1 gate2424(.O (I8246), .I (g6290));
INVX1 gate2425(.O (g1219), .I (I2218));
INVX1 gate2426(.O (g1640), .I (I2601));
INVX1 gate2427(.O (g2752), .I (g2343));
INVX1 gate2428(.O (g6373), .I (I8183));
INVX1 gate2429(.O (g3363), .I (g3110));
INVX1 gate2430(.O (g6491), .I (g6373));
INVX1 gate2431(.O (g5919), .I (I7689));
INVX1 gate2432(.O (I2671), .I (g1017));
INVX1 gate2433(.O (g1812), .I (I2867));
INVX1 gate2434(.O (I8721), .I (g6534));
INVX1 gate2435(.O (I2428), .I (g774));
INVX1 gate2436(.O (g4563), .I (g4190));
INVX1 gate2437(.O (g3053), .I (I4276));
INVX1 gate2438(.O (g1176), .I (I2190));
INVX1 gate2439(.O (g2265), .I (I3408));
INVX1 gate2440(.O (g3453), .I (g2628));
INVX1 gate2441(.O (g6283), .I (I7999));
INVX1 gate2442(.O (g6369), .I (I8171));
INVX1 gate2443(.O (g2042), .I (I3155));
INVX1 gate2444(.O (g6602), .I (I8674));
INVX1 gate2445(.O (I5249), .I (key_out_8));
INVX1 gate2446(.O (g6407), .I (I8235));
INVX1 gate2447(.O (g6578), .I (g6489));
INVX1 gate2448(.O (g4844), .I (I6540));
INVX1 gate2449(.O (g2164), .I (I3291));
INVX1 gate2450(.O (g1286), .I (g854));
INVX1 gate2451(.O (g2364), .I (I3516));
INVX1 gate2452(.O (g2233), .I (I3364));
INVX1 gate2453(.O (g4194), .I (I5612));
INVX1 gate2454(.O (g1911), .I (I3010));
INVX1 gate2455(.O (g4394), .I (I5885));
INVX1 gate2456(.O (g6535), .I (I8521));
INVX1 gate2457(.O (I6976), .I (g5136));
INVX1 gate2458(.O (g3912), .I (g3505));
INVX1 gate2459(.O (I2741), .I (key_out_124));
INVX1 gate2460(.O (g5527), .I (I7267));
INVX1 gate2461(.O (g6582), .I (I8614));
INVX1 gate2462(.O (I8940), .I (g6783));
INVX1 gate2463(.O (g4731), .I (I6359));
INVX1 gate2464(.O (I2910), .I (g1645));
INVX1 gate2465(.O (I3071), .I (g1504));
INVX1 gate2466(.O (g5647), .I (g5509));
INVX1 gate2467(.O (I3705), .I (g2316));
INVX1 gate2468(.O (I3471), .I (g1450));
INVX1 gate2469(.O (g2296), .I (I3441));
INVX1 gate2470(.O (g1733), .I (I2741));
INVX1 gate2471(.O (I2638), .I (key_out_122));
INVX1 gate2472(.O (g1270), .I (g844));
INVX1 gate2473(.O (g5546), .I (g5388));
INVX1 gate2474(.O (I5854), .I (g3857));
INVX1 gate2475(.O (I4465), .I (g2945));
INVX1 gate2476(.O (g6015), .I (g5857));
INVX1 gate2477(.O (g4705), .I (I6305));
INVX1 gate2478(.O (g6415), .I (I8255));
INVX1 gate2479(.O (I6126), .I (g4240));
INVX1 gate2480(.O (I6400), .I (g4473));
INVX1 gate2481(.O (g4242), .I (I5686));
INVX1 gate2482(.O (I2883), .I (key_out_123));
INVX1 gate2483(.O (I8671), .I (g6519));
INVX1 gate2484(.O (g5925), .I (I7707));
INVX1 gate2485(.O (I8030), .I (g6239));
INVX1 gate2486(.O (I4433), .I (g2103));
INVX1 gate2487(.O (g1324), .I (I2327));
INVX1 gate2488(.O (I5708), .I (g3942));
INVX1 gate2489(.O (I5520), .I (g3835));
INVX1 gate2490(.O (g6721), .I (I8857));
INVX1 gate2491(.O (I5640), .I (g3770));
INVX1 gate2492(.O (g5120), .I (I6772));
INVX1 gate2493(.O (I8564), .I (g6429));
INVX1 gate2494(.O (g2706), .I (I3861));
INVX1 gate2495(.O (I5252), .I (key_out_3));
INVX1 gate2496(.O (I3773), .I (g2524));
INVX1 gate2497(.O (g1177), .I (I2193));
INVX1 gate2498(.O (g4150), .I (I5532));
INVX1 gate2499(.O (I2165), .I (g690));
INVX1 gate2500(.O (g1206), .I (I2212));
INVX1 gate2501(.O (g4350), .I (g4010));
INVX1 gate2502(.O (g2888), .I (g1972));
INVX1 gate2503(.O (I7358), .I (g5565));
INVX1 gate2504(.O (I4195), .I (g2173));
INVX1 gate2505(.O (g2029), .I (I3134));
INVX1 gate2506(.O (I7506), .I (g5584));
INVX1 gate2507(.O (I5376), .I (g4014));
INVX1 gate2508(.O (g2171), .I (I3304));
INVX1 gate2509(.O (I4337), .I (g1934));
INVX1 gate2510(.O (I8910), .I (g6730));
INVX1 gate2511(.O (g2787), .I (g2405));
INVX1 gate2512(.O (g6502), .I (I8426));
INVX1 gate2513(.O (g2956), .I (g1861));
INVX1 gate2514(.O (I6023), .I (g4151));
INVX1 gate2515(.O (I8638), .I (g6553));
INVX1 gate2516(.O (g1287), .I (g855));
INVX1 gate2517(.O (g2675), .I (I3819));
INVX1 gate2518(.O (I3836), .I (g1832));
INVX1 gate2519(.O (I3212), .I (g1806));
INVX1 gate2520(.O (I7587), .I (g5605));
INVX1 gate2521(.O (g6940), .I (I9233));
INVX1 gate2522(.O (g4769), .I (g4606));
INVX1 gate2523(.O (g1849), .I (I2949));
INVX1 gate2524(.O (g3778), .I (g3388));
INVX1 gate2525(.O (g6188), .I (g5950));
INVX1 gate2526(.O (I2196), .I (g3));
INVX1 gate2527(.O (g5299), .I (I6949));
INVX1 gate2528(.O (g1781), .I (I2825));
INVX1 gate2529(.O (I6051), .I (g4185));
INVX1 gate2530(.O (g1898), .I (I2995));
INVX1 gate2531(.O (g3782), .I (g3388));
INVX1 gate2532(.O (I8217), .I (g6319));
INVX1 gate2533(.O (I8758), .I (g6562));
INVX1 gate2534(.O (I8066), .I (g6114));
INVX1 gate2535(.O (g5892), .I (g5742));
INVX1 gate2536(.O (I6327), .I (g4451));
INVX1 gate2537(.O (g6428), .I (I8290));
INVX1 gate2538(.O (g3075), .I (I4306));
INVX1 gate2539(.O (g4229), .I (g4059));
INVX1 gate2540(.O (g2109), .I (I3235));
INVX1 gate2541(.O (I7284), .I (g5383));
INVX1 gate2542(.O (I4255), .I (g2179));
INVX1 gate2543(.O (I6346), .I (g4563));
INVX1 gate2544(.O (I8165), .I (g6189));
INVX1 gate2545(.O (g4822), .I (g4614));
INVX1 gate2546(.O (g1291), .I (I2278));
INVX1 gate2547(.O (I5124), .I (g3719));
INVX1 gate2548(.O (I2067), .I (g686));
INVX1 gate2549(.O (g6564), .I (I8576));
INVX1 gate2550(.O (I5324), .I (g3466));
INVX1 gate2551(.O (I7832), .I (g5943));
INVX1 gate2552(.O (g6826), .I (I9011));
INVX1 gate2553(.O (I5469), .I (g3838));
INVX1 gate2554(.O (I2290), .I (g971));
INVX1 gate2555(.O (g1344), .I (I2379));
INVX1 gate2556(.O (I4354), .I (g1953));
INVX1 gate2557(.O (g5140), .I (I6798));
INVX1 gate2558(.O (I5177), .I (key_out_2));
INVX1 gate2559(.O (g3084), .I (I4321));
INVX1 gate2560(.O (g5478), .I (I7170));
INVX1 gate2561(.O (g1819), .I (I2877));
INVX1 gate2562(.O (I6753), .I (g4772));
INVX1 gate2563(.O (g2957), .I (g1861));
INVX1 gate2564(.O (I8803), .I (g6685));
INVX1 gate2565(.O (g1088), .I (I2119));
INVX1 gate2566(.O (g1852), .I (I2952));
INVX1 gate2567(.O (I6072), .I (g4385));
INVX1 gate2568(.O (g6609), .I (I8693));
INVX1 gate2569(.O (g5435), .I (I7113));
INVX1 gate2570(.O (g6308), .I (I8034));
INVX1 gate2571(.O (I3062), .I (g1776));
INVX1 gate2572(.O (g5082), .I (g4723));
INVX1 gate2573(.O (g2449), .I (I3584));
INVX1 gate2574(.O (I3620), .I (g1484));
INVX1 gate2575(.O (I3462), .I (g1450));
INVX1 gate2576(.O (I8538), .I (g6450));
INVX1 gate2577(.O (g2575), .I (I3684));
INVX1 gate2578(.O (g2865), .I (g2296));
INVX1 gate2579(.O (g6883), .I (I9116));
INVX1 gate2580(.O (g5876), .I (I7640));
INVX1 gate2581(.O (g4837), .I (g4473));
INVX1 gate2582(.O (I8509), .I (g6437));
INVX1 gate2583(.O (I2700), .I (g1173));
INVX1 gate2584(.O (g2604), .I (I3736));
INVX1 gate2585(.O (I4267), .I (g2525));
INVX1 gate2586(.O (g2098), .I (g1363));
INVX1 gate2587(.O (I4312), .I (g2555));
INVX1 gate2588(.O (g4620), .I (g4251));
INVX1 gate2589(.O (g4462), .I (I5977));
INVX1 gate2590(.O (g6589), .I (I8635));
INVX1 gate2591(.O (g945), .I (g536));
INVX1 gate2592(.O (I8662), .I (g6525));
INVX1 gate2593(.O (I3788), .I (g2554));
INVX1 gate2594(.O (g6466), .I (I8332));
INVX1 gate2595(.O (g5915), .I (I7679));
INVX1 gate2596(.O (g3952), .I (I5182));
INVX1 gate2597(.O (I6434), .I (g4622));
INVX1 gate2598(.O (I8467), .I (g6457));
INVX1 gate2599(.O (I8994), .I (g6789));
INVX1 gate2600(.O (I8290), .I (g6291));
INVX1 gate2601(.O (g1114), .I (I2150));
INVX1 gate2602(.O (g6165), .I (g5926));
INVX1 gate2603(.O (g6571), .I (I8597));
INVX1 gate2604(.O (g6365), .I (I8159));
INVX1 gate2605(.O (g2584), .I (I3705));
INVX1 gate2606(.O (g4788), .I (I6452));
INVX1 gate2607(.O (g6048), .I (g5824));
INVX1 gate2608(.O (I1841), .I (g207));
INVX1 gate2609(.O (g6711), .I (I8843));
INVX1 gate2610(.O (I8093), .I (g6122));
INVX1 gate2611(.O (g5110), .I (I6740));
INVX1 gate2612(.O (g4249), .I (I5699));
INVX1 gate2613(.O (g5310), .I (g5067));
INVX1 gate2614(.O (I3298), .I (g1725));
INVX1 gate2615(.O (g1825), .I (I2893));
INVX1 gate2616(.O (g6827), .I (I9014));
INVX1 gate2617(.O (g1650), .I (I2627));
INVX1 gate2618(.O (I3485), .I (g1450));
INVX1 gate2619(.O (g3527), .I (I4743));
INVX1 gate2620(.O (g809), .I (I1874));
INVX1 gate2621(.O (I6697), .I (g4722));
INVX1 gate2622(.O (g4842), .I (I6534));
INVX1 gate2623(.O (g849), .I (g598));
INVX1 gate2624(.O (g2268), .I (I3419));
INVX1 gate2625(.O (g4192), .I (I5606));
INVX1 gate2626(.O (g4392), .I (I5879));
INVX1 gate2627(.O (g3546), .I (g3095));
INVX1 gate2628(.O (g4485), .I (I5987));
INVX1 gate2629(.O (I2817), .I (key_out_124));
INVX1 gate2630(.O (g5824), .I (g5631));
INVX1 gate2631(.O (g1336), .I (I2361));
INVX1 gate2632(.O (g6803), .I (I8975));
INVX1 gate2633(.O (g3970), .I (I5236));
INVX1 gate2634(.O (g1594), .I (key_out_123));
INVX1 gate2635(.O (g4854), .I (I6570));
INVX1 gate2636(.O (g6538), .I (g6469));
INVX1 gate2637(.O (g1972), .I (I3083));
INVX1 gate2638(.O (I5923), .I (g4299));
INVX1 gate2639(.O (g6509), .I (I8447));
INVX1 gate2640(.O (g1806), .I (I2857));
INVX1 gate2641(.O (g5877), .I (I7643));
INVX1 gate2642(.O (g5590), .I (I7352));
INVX1 gate2643(.O (g1943), .I (I3050));
INVX1 gate2644(.O (I3708), .I (g1946));
INVX1 gate2645(.O (g3224), .I (I4471));
INVX1 gate2646(.O (g2086), .I (I3198));
INVX1 gate2647(.O (g2728), .I (I3890));
INVX1 gate2648(.O (I3031), .I (g1504));
INVX1 gate2649(.O (I4468), .I (g2583));
INVX1 gate2650(.O (g3320), .I (g3067));
INVX1 gate2651(.O (g6067), .I (g5788));
INVX1 gate2652(.O (g1887), .I (I2982));
INVX1 gate2653(.O (I3431), .I (g1275));
INVX1 gate2654(.O (g1122), .I (I2162));
INVX1 gate2655(.O (g6418), .I (I8264));
INVX1 gate2656(.O (g6467), .I (I8335));
INVX1 gate2657(.O (g1322), .I (I2321));
INVX1 gate2658(.O (g4520), .I (I6072));
INVX1 gate2659(.O (g1934), .I (I3037));
INVX1 gate2660(.O (I2041), .I (g680));
INVX1 gate2661(.O (I3376), .I (g1328));
INVX1 gate2662(.O (g4431), .I (I5938));
INVX1 gate2663(.O (g4252), .I (I5708));
INVX1 gate2664(.O (I1874), .I (g282));
INVX1 gate2665(.O (I3405), .I (g1321));
INVX1 gate2666(.O (g3906), .I (g3575));
INVX1 gate2667(.O (g2470), .I (I3602));
INVX1 gate2668(.O (g3789), .I (g3388));
INVX1 gate2669(.O (g5064), .I (I6706));
INVX1 gate2670(.O (g2025), .I (g1276));
INVX1 gate2671(.O (g6493), .I (g6375));
INVX1 gate2672(.O (g5899), .I (g5753));
INVX1 gate2673(.O (I6775), .I (g4790));
INVX1 gate2674(.O (g4376), .I (I5843));
INVX1 gate2675(.O (g4405), .I (I5910));
INVX1 gate2676(.O (g3771), .I (I4964));
INVX1 gate2677(.O (I5825), .I (g3914));
INVX1 gate2678(.O (g872), .I (g143));
INVX1 gate2679(.O (g1550), .I (g996));
INVX1 gate2680(.O (I6060), .I (g4380));
INVX1 gate2681(.O (g4286), .I (I5743));
INVX1 gate2682(.O (g4765), .I (I6403));
INVX1 gate2683(.O (I1880), .I (g276));
INVX1 gate2684(.O (I4198), .I (g2276));
INVX1 gate2685(.O (g3299), .I (g3049));
INVX1 gate2686(.O (g5563), .I (g5381));
INVX1 gate2687(.O (I4398), .I (g2086));
INVX1 gate2688(.O (g4911), .I (I6615));
INVX1 gate2689(.O (I3733), .I (g2031));
INVX1 gate2690(.O (g6700), .I (I8818));
INVX1 gate2691(.O (g1395), .I (I2428));
INVX1 gate2692(.O (g1891), .I (I2986));
INVX1 gate2693(.O (g1337), .I (I2364));
INVX1 gate2694(.O (g5237), .I (g5083));
INVX1 gate2695(.O (g3892), .I (g3575));
INVX1 gate2696(.O (g2678), .I (g2312));
INVX1 gate2697(.O (I3225), .I (g1813));
INVX1 gate2698(.O (g6421), .I (I8273));
INVX1 gate2699(.O (I2890), .I (key_out_122));
INVX1 gate2700(.O (I8585), .I (g6442));
INVX1 gate2701(.O (I5594), .I (g3821));
INVX1 gate2702(.O (g4270), .I (I5723));
INVX1 gate2703(.O (I7372), .I (g5493));
INVX1 gate2704(.O (g1807), .I (I2860));
INVX1 gate2705(.O (g4225), .I (g4059));
INVX1 gate2706(.O (g2682), .I (I3826));
INVX1 gate2707(.O (g2766), .I (g2361));
INVX1 gate2708(.O (I6995), .I (g5220));
INVX1 gate2709(.O (I1935), .I (g666));
INVX1 gate2710(.O (g2087), .I (g1352));
INVX1 gate2711(.O (g2105), .I (g1375));
INVX1 gate2712(.O (I6937), .I (g5124));
INVX1 gate2713(.O (I7143), .I (g5323));
INVX1 gate2714(.O (I8441), .I (g6419));
INVX1 gate2715(.O (g2801), .I (I4003));
INVX1 gate2716(.O (I2411), .I (g736));
INVX1 gate2717(.O (g5089), .I (I6723));
INVX1 gate2718(.O (g5489), .I (I7187));
INVX1 gate2719(.O (I5065), .I (g3714));
INVX1 gate2720(.O (g4124), .I (I5454));
INVX1 gate2721(.O (g714), .I (g131));
INVX1 gate2722(.O (I3540), .I (g1670));
INVX1 gate2723(.O (g4980), .I (g4678));
INVX1 gate2724(.O (g2748), .I (I3923));
INVX1 gate2725(.O (g6562), .I (I8570));
INVX1 gate2726(.O (I3206), .I (g1823));
INVX1 gate2727(.O (g5705), .I (I7466));
INVX1 gate2728(.O (I2992), .I (g1741));
INVX1 gate2729(.O (g3478), .I (g2695));
INVX1 gate2730(.O (g1142), .I (I2169));
INVX1 gate2731(.O (g2755), .I (g2350));
INVX1 gate2732(.O (I4258), .I (g2169));
INVX1 gate2733(.O (g5242), .I (g5085));
INVX1 gate2734(.O (I8168), .I (g6170));
INVX1 gate2735(.O (g6723), .I (I8863));
INVX1 gate2736(.O (g1255), .I (g161));
INVX1 gate2737(.O (I5033), .I (g3527));
INVX1 gate2738(.O (g6101), .I (I7799));
INVX1 gate2739(.O (g6817), .I (I8988));
INVX1 gate2740(.O (I5433), .I (g3728));
INVX1 gate2741(.O (g4206), .I (I5626));
INVX1 gate2742(.O (g3082), .I (I4315));
INVX1 gate2743(.O (g3482), .I (g2713));
INVX1 gate2744(.O (I8531), .I (g6444));
INVX1 gate2745(.O (g1692), .I (I2696));
INVX1 gate2746(.O (g6605), .I (I8681));
INVX1 gate2747(.O (g1726), .I (I2728));
INVX1 gate2748(.O (g3876), .I (I5109));
INVX1 gate2749(.O (g2173), .I (I3310));
INVX1 gate2750(.O (I6942), .I (g5124));
INVX1 gate2751(.O (g2091), .I (g1355));
INVX1 gate2752(.O (I5496), .I (g3839));
INVX1 gate2753(.O (g1960), .I (I3071));
INVX1 gate2754(.O (g2491), .I (I3620));
INVX1 gate2755(.O (g5150), .I (I6816));
INVX1 gate2756(.O (g4849), .I (I6555));
INVX1 gate2757(.O (g2169), .I (I3298));
INVX1 gate2758(.O (g2283), .I (I3428));
INVX1 gate2759(.O (I7113), .I (g5295));
INVX1 gate2760(.O (I8411), .I (g6415));
INVX1 gate2761(.O (I5337), .I (key_out_1));
INVX1 gate2762(.O (I5913), .I (g3751));
INVX1 gate2763(.O (g2602), .I (g2061));
INVX1 gate2764(.O (g6585), .I (I8623));
INVX1 gate2765(.O (g2007), .I (g1411));
INVX1 gate2766(.O (g5773), .I (I7514));
INVX1 gate2767(.O (g4399), .I (I5896));
INVX1 gate2768(.O (I3797), .I (g2125));
INVX1 gate2769(.O (I6250), .I (g4514));
INVX1 gate2770(.O (g2059), .I (g1402));
INVX1 gate2771(.O (g2920), .I (g1947));
INVX1 gate2772(.O (I4170), .I (g2157));
INVX1 gate2773(.O (g4781), .I (I6437));
INVX1 gate2774(.O (g6441), .I (I8309));
INVX1 gate2775(.O (I8074), .I (g6118));
INVX1 gate2776(.O (g2767), .I (g2364));
INVX1 gate2777(.O (g4900), .I (I6607));
INVX1 gate2778(.O (g1783), .I (I2831));
INVX1 gate2779(.O (g3110), .I (I4358));
INVX1 gate2780(.O (I4821), .I (g2877));
INVX1 gate2781(.O (I2688), .I (g1030));
INVX1 gate2782(.O (I2857), .I (key_out_126));
INVX1 gate2783(.O (g2535), .I (I3653));
INVX1 gate2784(.O (I3291), .I (g1714));
INVX1 gate2785(.O (g1979), .I (I3090));
INVX1 gate2786(.O (g1112), .I (g336));
INVX1 gate2787(.O (g1267), .I (g843));
INVX1 gate2788(.O (I7494), .I (g5691));
INVX1 gate2789(.O (g4510), .I (I6042));
INVX1 gate2790(.O (I3144), .I (g1319));
INVX1 gate2791(.O (g5918), .I (I7686));
INVX1 gate2792(.O (g1001), .I (I2044));
INVX1 gate2793(.O (g3002), .I (g2215));
INVX1 gate2794(.O (I8573), .I (g6435));
INVX1 gate2795(.O (I8863), .I (g6700));
INVX1 gate2796(.O (I4483), .I (g3082));
INVX1 gate2797(.O (g1293), .I (I2284));
INVX1 gate2798(.O (g6368), .I (I8168));
INVX1 gate2799(.O (g4144), .I (I5514));
INVX1 gate2800(.O (I8713), .I (g6522));
INVX1 gate2801(.O (I7593), .I (g5605));
INVX1 gate2802(.O (I3819), .I (g2044));
INVX1 gate2803(.O (g3236), .I (I4507));
INVX1 gate2804(.O (g1329), .I (I2340));
INVX1 gate2805(.O (I3694), .I (g1811));
INVX1 gate2806(.O (g1761), .I (I2788));
INVX1 gate2807(.O (g857), .I (g170));
INVX1 gate2808(.O (g5993), .I (g5872));
INVX1 gate2809(.O (g6531), .I (I8509));
INVX1 gate2810(.O (I5081), .I (key_out_8));
INVX1 gate2811(.O (I3923), .I (g2581));
INVX1 gate2812(.O (I4306), .I (g1898));
INVX1 gate2813(.O (I2760), .I (key_out_127));
INVX1 gate2814(.O (g2664), .I (I3808));
INVX1 gate2815(.O (I5481), .I (g3866));
INVX1 gate2816(.O (I3488), .I (g1295));
INVX1 gate2817(.O (g6743), .I (I8907));
INVX1 gate2818(.O (g6890), .I (I9137));
INVX1 gate2819(.O (g1830), .I (I2904));
INVX1 gate2820(.O (I5692), .I (g3942));
INVX1 gate2821(.O (I7264), .I (g5458));
INVX1 gate2822(.O (g4852), .I (I6564));
INVX1 gate2823(.O (g6505), .I (I8435));
INVX1 gate2824(.O (I3215), .I (g1820));
INVX1 gate2825(.O (g1221), .I (g46));
INVX1 gate2826(.O (g6411), .I (I8243));
INVX1 gate2827(.O (g6734), .I (I8894));
INVX1 gate2828(.O (g3222), .I (I4465));
INVX1 gate2829(.O (I3886), .I (g2215));
INVX1 gate2830(.O (I8857), .I (g6698));
INVX1 gate2831(.O (g1703), .I (I2707));
INVX1 gate2832(.O (I2608), .I (key_out_123));
INVX1 gate2833(.O (g5921), .I (I7695));
INVX1 gate2834(.O (g4215), .I (I5637));
INVX1 gate2835(.O (I2779), .I (g1038));
INVX1 gate2836(.O (I7996), .I (g6137));
INVX1 gate2837(.O (g6074), .I (g5794));
INVX1 gate2838(.O (g3064), .I (I4291));
INVX1 gate2839(.O (g3785), .I (g3466));
INVX1 gate2840(.O (g1624), .I (I2581));
INVX1 gate2841(.O (g1953), .I (I3062));
INVX1 gate2842(.O (I4003), .I (g2284));
INVX1 gate2843(.O (g5895), .I (g5742));
INVX1 gate2844(.O (g4114), .I (I5424));
INVX1 gate2845(.O (g4314), .I (g4080));
INVX1 gate2846(.O (I2588), .I (key_out_127));
INVX1 gate2847(.O (I3650), .I (g1650));
INVX1 gate2848(.O (g6080), .I (g5805));
INVX1 gate2849(.O (I2361), .I (g1075));
INVX1 gate2850(.O (g6573), .I (I8603));
INVX1 gate2851(.O (I4391), .I (g2275));
INVX1 gate2852(.O (g6713), .I (g6679));
INVX1 gate2853(.O (I3408), .I (g1644));
INVX1 gate2854(.O (g3237), .I (I4510));
INVX1 gate2855(.O (I7835), .I (g5926));
INVX1 gate2856(.O (I2327), .I (key_out_124));
INVX1 gate2857(.O (g6569), .I (I8591));
INVX1 gate2858(.O (g2030), .I (I3137));
INVX1 gate2859(.O (g5788), .I (I7587));
INVX1 gate2860(.O (g2430), .I (I3563));
INVX1 gate2861(.O (I2346), .I (key_out_127));
INVX1 gate2862(.O (g4136), .I (I5490));
INVX1 gate2863(.O (I8183), .I (g6176));
INVX1 gate2864(.O (I4223), .I (g2176));
INVX1 gate2865(.O (I8220), .I (g6322));
INVX1 gate2866(.O (g4768), .I (I6410));
INVX1 gate2867(.O (g1848), .I (I2946));
INVX1 gate2868(.O (I9140), .I (g6888));
INVX1 gate2869(.O (g2826), .I (g2481));
INVX1 gate2870(.O (g1699), .I (I2703));
INVX1 gate2871(.O (g1747), .I (I2760));
INVX1 gate2872(.O (g838), .I (key_out_12));
INVX1 gate2873(.O (I6075), .I (g4386));
INVX1 gate2874(.O (I2696), .I (g1156));
INVX1 gate2875(.O (I4757), .I (g2861));
INVX1 gate2876(.O (I7799), .I (g5918));
INVX1 gate2877(.O (I3065), .I (g1426));
INVX1 gate2878(.O (g3557), .I (g2598));
INVX1 gate2879(.O (I5746), .I (g4022));
INVX1 gate2880(.O (g4806), .I (g4473));
INVX1 gate2881(.O (g5392), .I (I7058));
INVX1 gate2882(.O (I8423), .I (g6423));
INVX1 gate2883(.O (I9035), .I (g6812));
INVX1 gate2884(.O (I6949), .I (g5050));
INVX1 gate2885(.O (g4943), .I (I6635));
INVX1 gate2886(.O (I3465), .I (g1724));
INVX1 gate2887(.O (I3322), .I (g1333));
INVX1 gate2888(.O (I9082), .I (g6849));
INVX1 gate2889(.O (g3705), .I (g3014));
INVX1 gate2890(.O (I8588), .I (g6443));
INVX1 gate2891(.O (I4522), .I (g2801));
INVX1 gate2892(.O (I2753), .I (g1174));
INVX1 gate2893(.O (g842), .I (g571));
INVX1 gate2894(.O (I6292), .I (g4434));
INVX1 gate2895(.O (I4315), .I (g2245));
INVX1 gate2896(.O (g3242), .I (g3083));
INVX1 gate2897(.O (g4122), .I (I5448));
INVX1 gate2898(.O (g4228), .I (I5668));
INVX1 gate2899(.O (g4322), .I (I5793));
INVX1 gate2900(.O (I2240), .I (g19));
INVX1 gate2901(.O (I1938), .I (g332));
INVX1 gate2902(.O (g2108), .I (I3232));
INVX1 gate2903(.O (g2609), .I (I3749));
INVX1 gate2904(.O (I6646), .I (g4687));
INVX1 gate2905(.O (g2308), .I (I3452));
INVX1 gate2906(.O (I8665), .I (g6527));
INVX1 gate2907(.O (I8051), .I (g6108));
INVX1 gate2908(.O (I7153), .I (g5358));
INVX1 gate2909(.O (g2883), .I (g1954));
INVX1 gate2910(.O (I6084), .I (g4391));
INVX1 gate2911(.O (I6039), .I (g4182));
INVX1 gate2912(.O (I5068), .I (key_out_4));
INVX1 gate2913(.O (I3096), .I (g1439));
INVX1 gate2914(.O (g1644), .I (I2611));
INVX1 gate2915(.O (I3496), .I (g1326));
INVX1 gate2916(.O (g715), .I (g135));
INVX1 gate2917(.O (I3550), .I (g1295));
INVX1 gate2918(.O (I7802), .I (g5920));
INVX1 gate2919(.O (g5708), .I (I7469));
INVX1 gate2920(.O (g1119), .I (I2159));
INVX1 gate2921(.O (g1319), .I (I2312));
INVX1 gate2922(.O (g2066), .I (g1341));
INVX1 gate2923(.O (g3150), .I (I4391));
INVX1 gate2924(.O (g5219), .I (I6885));
INVX1 gate2925(.O (I3137), .I (g1315));
INVX1 gate2926(.O (I8103), .I (g6134));
INVX1 gate2927(.O (I3395), .I (g1286));
INVX1 gate2928(.O (I3337), .I (g1338));
INVX1 gate2929(.O (g4496), .I (I6008));
INVX1 gate2930(.O (g1352), .I (I2391));
INVX1 gate2931(.O (I9110), .I (g6864));
INVX1 gate2932(.O (g1577), .I (g1001));
INVX1 gate2933(.O (g4550), .I (I6126));
INVX1 gate2934(.O (g3773), .I (g3466));
INVX1 gate2935(.O (g4845), .I (I6543));
INVX1 gate2936(.O (I4537), .I (g2877));
INVX1 gate2937(.O (I8696), .I (g6569));
INVX1 gate2938(.O (g2165), .I (I3294));
INVX1 gate2939(.O (g5958), .I (g5818));
INVX1 gate2940(.O (I2147), .I (g6));
INVX1 gate2941(.O (g6608), .I (I8690));
INVX1 gate2942(.O (g4195), .I (I5615));
INVX1 gate2943(.O (g4137), .I (I5493));
INVX1 gate2944(.O (g830), .I (g338));
INVX1 gate2945(.O (I5716), .I (g3942));
INVX1 gate2946(.O (g3769), .I (g3622));
INVX1 gate2947(.O (I9002), .I (g6802));
INVX1 gate2948(.O (g2827), .I (g2485));
INVX1 gate2949(.O (I6952), .I (g5124));
INVX1 gate2950(.O (I5848), .I (g3856));
INVX1 gate2951(.O (g3836), .I (I5033));
INVX1 gate2952(.O (g3212), .I (I4455));
INVX1 gate2953(.O (g6423), .I (I8279));
INVX1 gate2954(.O (I4243), .I (g1853));
INVX1 gate2955(.O (g2333), .I (I3485));
INVX1 gate2956(.O (I8240), .I (g6287));
INVX1 gate2957(.O (g1975), .I (I3086));
INVX1 gate2958(.O (I5699), .I (g3844));
INVX1 gate2959(.O (g4807), .I (g4473));
INVX1 gate2960(.O (I9236), .I (g6939));
INVX1 gate2961(.O (g3967), .I (I5223));
INVX1 gate2962(.O (I6561), .I (g4707));
INVX1 gate2963(.O (g6588), .I (I8632));
INVX1 gate2964(.O (I4935), .I (g3369));
INVX1 gate2965(.O (I2596), .I (g985));
INVX1 gate2966(.O (g6161), .I (g5926));
INVX1 gate2967(.O (g1274), .I (g856));
INVX1 gate2968(.O (g6361), .I (I8147));
INVX1 gate2969(.O (g1426), .I (I2445));
INVX1 gate2970(.O (g2196), .I (I3337));
INVX1 gate2971(.O (I7600), .I (g5605));
INVX1 gate2972(.O (g2803), .I (g2440));
INVX1 gate2973(.O (I6004), .I (g4159));
INVX1 gate2974(.O (g3229), .I (I4486));
INVX1 gate2975(.O (I6986), .I (g5230));
INVX1 gate2976(.O (g6051), .I (g5824));
INVX1 gate2977(.O (g5270), .I (I6927));
INVX1 gate2978(.O (g804), .I (I1871));
INVX1 gate2979(.O (I3255), .I (g1650));
INVX1 gate2980(.O (g2538), .I (I3656));
INVX1 gate2981(.O (g1325), .I (I2330));
INVX1 gate2982(.O (g1821), .I (I2883));
INVX1 gate2983(.O (g844), .I (g578));
INVX1 gate2984(.O (I3481), .I (g1461));
INVX1 gate2985(.O (I8034), .I (g6242));
INVX1 gate2986(.O (g4142), .I (I5508));
INVX1 gate2987(.O (g4248), .I (I5696));
INVX1 gate2988(.O (g2509), .I (I3635));
INVX1 gate2989(.O (I6546), .I (g4692));
INVX1 gate2990(.O (I3726), .I (g2030));
INVX1 gate2991(.O (g4815), .I (I6495));
INVX1 gate2992(.O (I5644), .I (g4059));
INVX1 gate2993(.O (I8147), .I (g6182));
INVX1 gate2994(.O (g5124), .I (I6780));
INVX1 gate2995(.O (g6103), .I (I7805));
INVX1 gate2996(.O (I5119), .I (g3714));
INVX1 gate2997(.O (g4692), .I (I6280));
INVX1 gate2998(.O (g2467), .I (I3599));
INVX1 gate2999(.O (I8681), .I (g6566));
INVX1 gate3000(.O (g4726), .I (I6352));
INVX1 gate3001(.O (g5469), .I (I7153));
INVX1 gate3002(.O (g4154), .I (I5548));
INVX1 gate3003(.O (I2601), .I (key_out_126));
INVX1 gate3004(.O (g6696), .I (I8806));
INVX1 gate3005(.O (g1636), .I (I2593));
INVX1 gate3006(.O (g3921), .I (g3512));
INVX1 gate3007(.O (g5540), .I (I7284));
INVX1 gate3008(.O (I5577), .I (g4022));
INVX1 gate3009(.O (g1106), .I (I2128));
INVX1 gate3010(.O (g6732), .I (I8888));
INVX1 gate3011(.O (g853), .I (g642));
INVX1 gate3012(.O (g2256), .I (I3395));
INVX1 gate3013(.O (g1790), .I (I2842));
INVX1 gate3014(.O (I2922), .I (g1774));
INVX1 gate3015(.O (g6508), .I (I8444));
INVX1 gate3016(.O (I5893), .I (g3747));
INVX1 gate3017(.O (I3979), .I (g1836));
INVX1 gate3018(.O (I2581), .I (g946));
INVX1 gate3019(.O (I3112), .I (g1439));
INVX1 gate3020(.O (g1461), .I (I2460));
INVX1 gate3021(.O (g3462), .I (g2679));
INVX1 gate3022(.O (g1756), .I (I2779));
INVX1 gate3023(.O (g2381), .I (I3528));
INVX1 gate3024(.O (I6789), .I (g4871));
INVX1 gate3025(.O (g4783), .I (I6441));
INVX1 gate3026(.O (g6043), .I (g5824));
INVX1 gate3027(.O (I7871), .I (g6097));
INVX1 gate3028(.O (I2460), .I (g952));
INVX1 gate3029(.O (I3001), .I (g1267));
INVX1 gate3030(.O (g4112), .I (I5418));
INVX1 gate3031(.O (g4218), .I (I5640));
INVX1 gate3032(.O (g2197), .I (I3340));
INVX1 gate3033(.O (g4267), .I (I5720));
INVX1 gate3034(.O (I4166), .I (g2390));
INVX1 gate3035(.O (g2397), .I (I3540));
INVX1 gate3036(.O (I4366), .I (g2244));
INVX1 gate3037(.O (g5199), .I (I6867));
INVX1 gate3038(.O (g5399), .I (I7065));
INVX1 gate3039(.O (g1046), .I (g489));
INVX1 gate3040(.O (I3761), .I (g2505));
INVX1 gate3041(.O (g3788), .I (g3466));
INVX1 gate3042(.O (g6034), .I (g5824));
INVX1 gate3043(.O (g6434), .I (I8300));
INVX1 gate3044(.O (g6565), .I (I8579));
INVX1 gate3045(.O (I6299), .I (g4438));
INVX1 gate3046(.O (g4293), .I (I5750));
INVX1 gate3047(.O (g4129), .I (I5469));
INVX1 gate3048(.O (g5797), .I (I7596));
INVX1 gate3049(.O (I3830), .I (g2179));
INVX1 gate3050(.O (I2995), .I (g1742));
INVX1 gate3051(.O (g6147), .I (I7871));
INVX1 gate3052(.O (g1345), .I (I2382));
INVX1 gate3053(.O (g1841), .I (I2929));
INVX1 gate3054(.O (g6347), .I (I8103));
INVX1 gate3055(.O (I1832), .I (g143));
INVX1 gate3056(.O (I2479), .I (g1049));
INVX1 gate3057(.O (I7339), .I (g5540));
INVX1 gate3058(.O (g1191), .I (g38));
INVX1 gate3059(.O (I2668), .I (g1011));
INVX1 gate3060(.O (g1391), .I (I2424));
INVX1 gate3061(.O (I1853), .I (g211));
INVX1 gate3062(.O (g3192), .I (I4429));
INVX1 gate3063(.O (g6533), .I (I8515));
INVX1 gate3064(.O (g3085), .I (I4324));
INVX1 gate3065(.O (I3746), .I (g2035));
INVX1 gate3066(.O (I7838), .I (g5947));
INVX1 gate3067(.O (g4727), .I (I6355));
INVX1 gate3068(.O (I4964), .I (key_out_11));
INVX1 gate3069(.O (g3485), .I (g2986));
INVX1 gate3070(.O (I2190), .I (g297));
INVX1 gate3071(.O (g1695), .I (g1106));
INVX1 gate3072(.O (g6697), .I (I8809));
INVX1 gate3073(.O (g1637), .I (I2596));
INVX1 gate3074(.O (g1107), .I (I2131));
INVX1 gate3075(.O (g2631), .I (I3773));
INVX1 gate3076(.O (g6596), .I (I8656));
INVX1 gate3077(.O (g3854), .I (I5071));
INVX1 gate3078(.O (I5106), .I (g3247));
INVX1 gate3079(.O (I8597), .I (g6445));
INVX1 gate3080(.O (g2817), .I (g2461));
INVX1 gate3081(.O (I6244), .I (g4519));
INVX1 gate3082(.O (I7077), .I (g5281));
INVX1 gate3083(.O (g4703), .I (I6299));
INVX1 gate3084(.O (g6413), .I (I8249));
INVX1 gate3085(.O (I5790), .I (g3803));
INVX1 gate3086(.O (g1858), .I (I2964));
INVX1 gate3087(.O (I6078), .I (g4387));
INVX1 gate3088(.O (I6340), .I (g4561));
INVX1 gate3089(.O (I7643), .I (g5752));
INVX1 gate3090(.O (I3068), .I (g1439));
INVX1 gate3091(.O (g5923), .I (I7701));
INVX1 gate3092(.O (I9038), .I (g6833));
INVX1 gate3093(.O (I3468), .I (g1802));
INVX1 gate3094(.O (I4279), .I (g2230));
INVX1 gate3095(.O (I5756), .I (g3922));
INVX1 gate3096(.O (g6820), .I (I8997));
INVX1 gate3097(.O (g4624), .I (g4265));
INVX1 gate3098(.O (I6959), .I (g5089));
INVX1 gate3099(.O (I5622), .I (g3914));
INVX1 gate3100(.O (g3219), .I (I4462));
INVX1 gate3101(.O (I5027), .I (key_out_2));
INVX1 gate3102(.O (I4318), .I (g2171));
INVX1 gate3103(.O (I7634), .I (g5727));
INVX1 gate3104(.O (I5427), .I (g3726));
INVX1 gate3105(.O (g3031), .I (I4246));
INVX1 gate3106(.O (g1115), .I (g40));
INVX1 gate3107(.O (g6117), .I (g5880));
INVX1 gate3108(.O (g1315), .I (I2296));
INVX1 gate3109(.O (g1811), .I (I2864));
INVX1 gate3110(.O (g1642), .I (g809));
INVX1 gate3111(.O (I8479), .I (g6482));
INVX1 gate3112(.O (g2585), .I (I3708));
INVX1 gate3113(.O (I7104), .I (g5273));
INVX1 gate3114(.O (I5904), .I (g3749));
INVX1 gate3115(.O (I8668), .I (g6530));
INVX1 gate3116(.O (g5886), .I (g5753));
INVX1 gate3117(.O (I8840), .I (g6657));
INVX1 gate3118(.O (g2041), .I (I3152));
INVX1 gate3119(.O (g6601), .I (I8671));
INVX1 gate3120(.O (I5514), .I (g3882));
INVX1 gate3121(.O (I3349), .I (g1334));
INVX1 gate3122(.O (I2053), .I (g684));
INVX1 gate3123(.O (g5114), .I (I6756));
INVX1 gate3124(.O (I5403), .I (g3970));
INVX1 gate3125(.O (g5314), .I (I6972));
INVX1 gate3126(.O (I2453), .I (g952));
INVX1 gate3127(.O (g1654), .I (g878));
INVX1 gate3128(.O (g4716), .I (I6330));
INVX1 gate3129(.O (g4149), .I (I5529));
INVX1 gate3130(.O (g6922), .I (I9203));
INVX1 gate3131(.O (I8156), .I (g6167));
INVX1 gate3132(.O (I3198), .I (g1819));
INVX1 gate3133(.O (I3855), .I (g2550));
INVX1 gate3134(.O (I5391), .I (g3975));
INVX1 gate3135(.O (g3911), .I (I5148));
INVX1 gate3136(.O (g6581), .I (g6493));
INVX1 gate3137(.O (g4848), .I (I6552));
INVX1 gate3138(.O (I5637), .I (g3914));
INVX1 gate3139(.O (g1880), .I (g1603));
INVX1 gate3140(.O (g4198), .I (I5618));
INVX1 gate3141(.O (g4699), .I (I6289));
INVX1 gate3142(.O (g6597), .I (I8659));
INVX1 gate3143(.O (g4855), .I (I6573));
INVX1 gate3144(.O (g4398), .I (I5893));
INVX1 gate3145(.O (g2772), .I (I3961));
INVX1 gate3146(.O (I4321), .I (g1917));
INVX1 gate3147(.O (g5136), .I (I6786));
INVX1 gate3148(.O (g3225), .I (I4474));
INVX1 gate3149(.O (I5223), .I (g3537));
INVX1 gate3150(.O (g2743), .I (g2333));
INVX1 gate3151(.O (g6784), .I (I8940));
INVX1 gate3152(.O (g2890), .I (g1875));
INVX1 gate3153(.O (g3073), .I (I4300));
INVX1 gate3154(.O (g1978), .I (g1387));
INVX1 gate3155(.O (g3796), .I (g3388));
INVX1 gate3156(.O (g1017), .I (I2053));
INVX1 gate3157(.O (I2929), .I (g1659));
INVX1 gate3158(.O (g798), .I (I1868));
INVX1 gate3159(.O (g2505), .I (I3629));
INVX1 gate3160(.O (I3644), .I (g1685));
INVX1 gate3161(.O (g3124), .I (I4371));
INVX1 gate3162(.O (g1935), .I (I3040));
INVX1 gate3163(.O (g3980), .I (I5264));
INVX1 gate3164(.O (g2856), .I (g2010));
INVX1 gate3165(.O (g2734), .I (I3902));
INVX1 gate3166(.O (I8432), .I (g6411));
INVX1 gate3167(.O (I3319), .I (g1636));
INVX1 gate3168(.O (g1982), .I (I3093));
INVX1 gate3169(.O (g754), .I (I1850));
INVX1 gate3170(.O (g4524), .I (I6084));
INVX1 gate3171(.O (g836), .I (g349));
INVX1 gate3172(.O (I8453), .I (g6414));
INVX1 gate3173(.O (g6840), .I (I9041));
INVX1 gate3174(.O (I4519), .I (g2788));
INVX1 gate3175(.O (g4644), .I (I6231));
INVX1 gate3176(.O (I3152), .I (g1322));
INVX1 gate3177(.O (I3258), .I (g1760));
INVX1 gate3178(.O (g3540), .I (I4762));
INVX1 gate3179(.O (I3352), .I (g1285));
INVX1 gate3180(.O (g1328), .I (I2337));
INVX1 gate3181(.O (g5887), .I (g5742));
INVX1 gate3182(.O (g4119), .I (I5439));
INVX1 gate3183(.O (g5465), .I (I7143));
INVX1 gate3184(.O (g1542), .I (g878));
INVX1 gate3185(.O (g1330), .I (I2343));
INVX1 gate3186(.O (g3177), .I (I4414));
INVX1 gate3187(.O (I3717), .I (g2154));
INVX1 gate3188(.O (g5230), .I (I6895));
INVX1 gate3189(.O (g845), .I (g582));
INVX1 gate3190(.O (g4152), .I (I5542));
INVX1 gate3191(.O (g6501), .I (I8423));
INVX1 gate3192(.O (g4577), .I (g4202));
INVX1 gate3193(.O (g4717), .I (g4465));
INVX1 gate3194(.O (g5433), .I (I7107));
INVX1 gate3195(.O (I5654), .I (g3742));
INVX1 gate3196(.O (I6930), .I (g5017));
INVX1 gate3197(.O (g2863), .I (g2296));
INVX1 gate3198(.O (I6464), .I (g4562));
INVX1 gate3199(.O (I3599), .I (g1484));
INVX1 gate3200(.O (g2713), .I (I3868));
INVX1 gate3201(.O (I3274), .I (g1773));
INVX1 gate3202(.O (g4386), .I (I5865));
INVX1 gate3203(.O (g3199), .I (g1861));
INVX1 gate3204(.O (g5550), .I (g5331));
INVX1 gate3205(.O (I3614), .I (g1295));
INVX1 gate3206(.O (g3781), .I (I4976));
INVX1 gate3207(.O (I3370), .I (g1805));
INVX1 gate3208(.O (g5137), .I (I6789));
INVX1 gate3209(.O (g5395), .I (I7061));
INVX1 gate3210(.O (g5891), .I (g5731));
INVX1 gate3211(.O (g3898), .I (g3575));
INVX1 gate3212(.O (g3900), .I (g3575));
INVX1 gate3213(.O (I3325), .I (g1340));
INVX1 gate3214(.O (g4426), .I (I5929));
INVX1 gate3215(.O (I2735), .I (g1118));
INVX1 gate3216(.O (g3797), .I (g3388));
INVX1 gate3217(.O (I9085), .I (g6850));
INVX1 gate3218(.O (g1902), .I (I3001));
INVX1 gate3219(.O (g6163), .I (g5926));
INVX1 gate3220(.O (g4614), .I (g4308));
INVX1 gate3221(.O (I2782), .I (key_out_125));
INVX1 gate3222(.O (I7679), .I (g5726));
INVX1 gate3223(.O (g6363), .I (I8153));
INVX1 gate3224(.O (g4370), .I (I5831));
INVX1 gate3225(.O (I8626), .I (g6543));
INVX1 gate3226(.O (g3510), .I (g2709));
INVX1 gate3227(.O (I5612), .I (g3910));
INVX1 gate3228(.O (g6032), .I (g5770));
INVX1 gate3229(.O (g4125), .I (I5457));
INVX1 gate3230(.O (g2688), .I (I3836));
INVX1 gate3231(.O (g2857), .I (I4059));
INVX1 gate3232(.O (g3291), .I (g3037));
INVX1 gate3233(.O (I3083), .I (g1426));
INVX1 gate3234(.O (g2976), .I (g2197));
INVX1 gate3235(.O (g1823), .I (I2887));
INVX1 gate3236(.O (I2949), .I (g1263));
INVX1 gate3237(.O (g1366), .I (I2402));
INVX1 gate3238(.O (g5266), .I (I6923));
INVX1 gate3239(.O (I2627), .I (g1053));
INVX1 gate3240(.O (g1056), .I (g89));
INVX1 gate3241(.O (g6568), .I (I8588));
INVX1 gate3242(.O (I5328), .I (g3502));
INVX1 gate3243(.O (g1529), .I (g1076));
INVX1 gate3244(.O (I7805), .I (g5923));
INVX1 gate3245(.O (I5542), .I (g3984));
INVX1 gate3246(.O (I2998), .I (g1257));
INVX1 gate3247(.O (g1649), .I (g985));
INVX1 gate3248(.O (g1348), .I (I2385));
INVX1 gate3249(.O (g3259), .I (g2996));
INVX1 gate3250(.O (I4358), .I (g2525));
INVX1 gate3251(.O (g5248), .I (g4911));
INVX1 gate3252(.O (g4636), .I (g4286));
INVX1 gate3253(.O (g1355), .I (I2394));
INVX1 gate3254(.O (g4106), .I (I5400));
INVX1 gate3255(.O (g5255), .I (g4933));
INVX1 gate3256(.O (g3852), .I (I5065));
INVX1 gate3257(.O (I9031), .I (g6809));
INVX1 gate3258(.O (g2760), .I (I3942));
INVX1 gate3259(.O (g3488), .I (g2728));
INVX1 gate3260(.O (I8894), .I (g6709));
INVX1 gate3261(.O (g4790), .I (I6456));
INVX1 gate3262(.O (g5692), .I (I7451));
INVX1 gate3263(.O (I4587), .I (g2962));
INVX1 gate3264(.O (g5097), .I (I6733));
INVX1 gate3265(.O (g5726), .I (I7487));
INVX1 gate3266(.O (g4187), .I (I5591));
INVX1 gate3267(.O (I9176), .I (g6881));
INVX1 gate3268(.O (g4387), .I (I5868));
INVX1 gate3269(.O (I9005), .I (g6817));
INVX1 gate3270(.O (g1063), .I (g675));
INVX1 gate3271(.O (g3886), .I (g3346));
INVX1 gate3272(.O (g4622), .I (g4252));
INVX1 gate3273(.O (g2608), .I (I3746));
INVX1 gate3274(.O (I2919), .I (g1787));
INVX1 gate3275(.O (g2779), .I (g2394));
INVX1 gate3276(.O (g4904), .I (g4812));
INVX1 gate3277(.O (g3114), .I (I4362));
INVX1 gate3278(.O (I2952), .I (g1594));
INVX1 gate3279(.O (g1279), .I (g848));
INVX1 gate3280(.O (g4514), .I (I6054));
INVX1 gate3281(.O (g1720), .I (g1111));
INVX1 gate3282(.O (g4003), .I (g3441));
INVX1 gate3283(.O (g1118), .I (g36));
INVX1 gate3284(.O (I3391), .I (g1646));
INVX1 gate3285(.O (g1318), .I (I2309));
INVX1 gate3286(.O (g4403), .I (I5904));
INVX1 gate3287(.O (I5490), .I (g3832));
INVX1 gate3288(.O (g5112), .I (I6750));
INVX1 gate3289(.O (g2588), .I (I3717));
INVX1 gate3290(.O (g4145), .I (I5517));
INVX1 gate3291(.O (g4841), .I (I6531));
INVX1 gate3292(.O (I8603), .I (g6449));
INVX1 gate3293(.O (g2361), .I (I3513));
INVX1 gate3294(.O (I6769), .I (g4786));
INVX1 gate3295(.O (g4763), .I (I6397));
INVX1 gate3296(.O (g4191), .I (I5603));
INVX1 gate3297(.O (g4391), .I (I5876));
INVX1 gate3298(.O (I5056), .I (key_out_7));
INVX1 gate3299(.O (I2986), .I (g1504));
INVX1 gate3300(.O (I3307), .I (g1339));
INVX1 gate3301(.O (g1193), .I (I2204));
INVX1 gate3302(.O (I5529), .I (g3854));
INVX1 gate3303(.O (I4420), .I (g2096));
INVX1 gate3304(.O (I5148), .I (g3450));
INVX1 gate3305(.O (g3136), .I (I4382));
INVX1 gate3306(.O (g2327), .I (I3481));
INVX1 gate3307(.O (I6918), .I (g5124));
INVX1 gate3308(.O (I4507), .I (g2739));
INVX1 gate3309(.O (g5329), .I (I6989));
INVX1 gate3310(.O (g1549), .I (g878));
INVX1 gate3311(.O (g4107), .I (I5403));
INVX1 gate3312(.O (I7042), .I (g5310));
INVX1 gate3313(.O (g947), .I (g74));
INVX1 gate3314(.O (g6894), .I (I9149));
INVX1 gate3315(.O (g1834), .I (I2916));
INVX1 gate3316(.O (I4794), .I (g2814));
INVX1 gate3317(.O (g4307), .I (I5774));
INVX1 gate3318(.O (I5851), .I (g3739));
INVX1 gate3319(.O (g4536), .I (I6118));
INVX1 gate3320(.O (I3858), .I (g2197));
INVX1 gate3321(.O (I8702), .I (g6572));
INVX1 gate3322(.O (g2346), .I (I3496));
INVX1 gate3323(.O (g6735), .I (I8897));
INVX1 gate3324(.O (I3016), .I (g1754));
INVX1 gate3325(.O (I2970), .I (g1504));
INVX1 gate3326(.O (g5727), .I (I7490));
INVX1 gate3327(.O (I7164), .I (g5433));
INVX1 gate3328(.O (g2103), .I (I3225));
INVX1 gate3329(.O (g858), .I (g301));
INVX1 gate3330(.O (I2925), .I (g1762));
INVX1 gate3331(.O (g4858), .I (I6582));
INVX1 gate3332(.O (I3522), .I (g1664));
INVX1 gate3333(.O (g4016), .I (I5320));
INVX1 gate3334(.O (I3115), .I (g1519));
INVX1 gate3335(.O (I3251), .I (g1471));
INVX1 gate3336(.O (I3811), .I (g2145));
INVX1 gate3337(.O (I8276), .I (g6303));
INVX1 gate3338(.O (g1321), .I (I2318));
INVX1 gate3339(.O (I3047), .I (g1426));
INVX1 gate3340(.O (g1670), .I (I2648));
INVX1 gate3341(.O (g3228), .I (I4483));
INVX1 gate3342(.O (g3465), .I (g2986));
INVX1 gate3343(.O (g3322), .I (g3070));
INVX1 gate3344(.O (I5463), .I (g3783));
INVX1 gate3345(.O (g3230), .I (I4489));
INVX1 gate3346(.O (g4522), .I (I6078));
INVX1 gate3347(.O (g4115), .I (I5427));
INVX1 gate3348(.O (g2753), .I (I3927));
INVX1 gate3349(.O (g4251), .I (I5705));
INVX1 gate3350(.O (g1232), .I (I2228));
INVX1 gate3351(.O (I4300), .I (g2234));
INVX1 gate3352(.O (g6526), .I (I8494));
INVX1 gate3353(.O (g1813), .I (I2870));
INVX1 gate3354(.O (I8527), .I (g6440));
INVX1 gate3355(.O (I8647), .I (g6528));
INVX1 gate3356(.O (I2617), .I (key_out_127));
INVX1 gate3357(.O (I5720), .I (g4022));
INVX1 gate3358(.O (g2043), .I (I3158));
INVX1 gate3359(.O (g6039), .I (g5824));
INVX1 gate3360(.O (I8764), .I (g6564));
INVX1 gate3361(.O (g2443), .I (I3578));
INVX1 gate3362(.O (g6484), .I (g6361));
INVX1 gate3363(.O (g3096), .I (I4343));
INVX1 gate3364(.O (g5468), .I (I7150));
INVX1 gate3365(.O (g1519), .I (I2491));
INVX1 gate3366(.O (g1740), .I (g1116));
INVX1 gate3367(.O (I7012), .I (g5316));
INVX1 gate3368(.O (g6850), .I (I9077));
INVX1 gate3369(.O (I6895), .I (g5010));
INVX1 gate3370(.O (I1835), .I (g205));
INVX1 gate3371(.O (g3845), .I (I5050));
INVX1 gate3372(.O (I5843), .I (g3851));
INVX1 gate3373(.O (g2316), .I (I3468));
INVX1 gate3374(.O (I3537), .I (g1305));
INVX1 gate3375(.O (I8503), .I (g6434));
INVX1 gate3376(.O (g1552), .I (g1030));
INVX1 gate3377(.O (I5457), .I (g3766));
INVX1 gate3378(.O (g2565), .I (I3675));
INVX1 gate3379(.O (g6583), .I (I8617));
INVX1 gate3380(.O (g850), .I (g602));
INVX1 gate3381(.O (g5576), .I (g5415));
INVX1 gate3382(.O (g4537), .I (g4410));
INVX1 gate3383(.O (I7029), .I (g5149));
INVX1 gate3384(.O (g2347), .I (I3499));
INVX1 gate3385(.O (I5686), .I (g3942));
INVX1 gate3386(.O (I4123), .I (g2043));
INVX1 gate3387(.O (g3807), .I (I5006));
INVX1 gate3388(.O (g1586), .I (g1052));
INVX1 gate3389(.O (g3859), .I (I5078));
INVX1 gate3390(.O (g6276), .I (I7960));
INVX1 gate3391(.O (g4612), .I (g4320));
INVX1 gate3392(.O (g2914), .I (g1928));
INVX1 gate3393(.O (g6616), .I (I8710));
INVX1 gate3394(.O (I3629), .I (g1759));
INVX1 gate3395(.O (g6561), .I (I8567));
INVX1 gate3396(.O (I3328), .I (g1273));
INVX1 gate3397(.O (I2738), .I (key_out_120));
INVX1 gate3398(.O (I8617), .I (g6539));
INVX1 gate3399(.O (g1341), .I (I2376));
INVX1 gate3400(.O (g2413), .I (I3553));
INVX1 gate3401(.O (I4351), .I (g2233));
INVX1 gate3402(.O (g3342), .I (g3086));
INVX1 gate3403(.O (g4128), .I (I5466));
INVX1 gate3404(.O (g1710), .I (g1109));
INVX1 gate3405(.O (g4629), .I (g4276));
INVX1 gate3406(.O (I6485), .I (g4603));
INVX1 gate3407(.O (g6527), .I (I8497));
INVX1 gate3408(.O (g6404), .I (I8226));
INVX1 gate3409(.O (g4328), .I (g4092));
INVX1 gate3410(.O (I2140), .I (g28));
INVX1 gate3411(.O (g1645), .I (I2614));
INVX1 gate3412(.O (I2340), .I (g1142));
INVX1 gate3413(.O (g4130), .I (I5472));
INVX1 gate3414(.O (I5938), .I (g4351));
INVX1 gate3415(.O (I7963), .I (g6276));
INVX1 gate3416(.O (I3800), .I (g2145));
INVX1 gate3417(.O (g3481), .I (g2612));
INVX1 gate3418(.O (I2907), .I (g1498));
INVX1 gate3419(.O (g2820), .I (g2470));
INVX1 gate3420(.O (g2936), .I (g2026));
INVX1 gate3421(.O (g5524), .I (I7264));
INVX1 gate3422(.O (g6503), .I (I8429));
INVX1 gate3423(.O (g3354), .I (g3096));
INVX1 gate3424(.O (I4410), .I (g2088));
INVX1 gate3425(.O (I7808), .I (g5919));
INVX1 gate3426(.O (g2117), .I (I3244));
INVX1 gate3427(.O (g3960), .I (I5204));
INVX1 gate3428(.O (g2317), .I (I3471));
INVX1 gate3429(.O (g5119), .I (I6769));
INVX1 gate3430(.O (g6925), .I (I9208));
INVX1 gate3431(.O (I7707), .I (g5701));
INVX1 gate3432(.O (I5606), .I (g3821));
INVX1 gate3433(.O (g1659), .I (I2638));
INVX1 gate3434(.O (g1358), .I (g1119));
INVX1 gate3435(.O (g5352), .I (I7002));
INVX1 gate3436(.O (g5577), .I (g5420));
INVX1 gate3437(.O (g4213), .I (I5633));
INVX1 gate3438(.O (g5717), .I (I7478));
INVX1 gate3439(.O (I3902), .I (g2576));
INVX1 gate3440(.O (g6120), .I (I7832));
INVX1 gate3441(.O (g2922), .I (g1960));
INVX1 gate3442(.O (g1587), .I (key_out_122));
INVX1 gate3443(.O (I6812), .I (g5110));
INVX1 gate3444(.O (I8991), .I (g6788));
INVX1 gate3445(.O (g3783), .I (I4980));
INVX1 gate3446(.O (g1111), .I (I2143));
INVX1 gate3447(.O (I3090), .I (g1504));
INVX1 gate3448(.O (I9008), .I (g6818));
INVX1 gate3449(.O (g5893), .I (g5753));
INVX1 gate3450(.O (g1275), .I (g842));
INVX1 gate3451(.O (g6277), .I (I7963));
INVX1 gate3452(.O (g2581), .I (I3694));
INVX1 gate3453(.O (I3823), .I (g2125));
INVX1 gate3454(.O (g3267), .I (g3030));
INVX1 gate3455(.O (I4667), .I (g2908));
INVX1 gate3456(.O (g3312), .I (I4587));
INVX1 gate3457(.O (I7865), .I (g6095));
INVX1 gate3458(.O (I4343), .I (g2525));
INVX1 gate3459(.O (g2060), .I (g1369));
INVX1 gate3460(.O (g6617), .I (I8713));
INVX1 gate3461(.O (g6906), .I (I9185));
INVX1 gate3462(.O (g5975), .I (g5821));
INVX1 gate3463(.O (g4512), .I (I6048));
INVX1 gate3464(.O (I4282), .I (g2525));
INVX1 gate3465(.O (g2460), .I (I3590));
INVX1 gate3466(.O (I7604), .I (g5605));
INVX1 gate3467(.O (I8907), .I (g6702));
INVX1 gate3468(.O (I3056), .I (g1519));
INVX1 gate3469(.O (g3001), .I (I4198));
INVX1 gate3470(.O (g1174), .I (g37));
INVX1 gate3471(.O (g4823), .I (I6507));
INVX1 gate3472(.O (I2663), .I (g1006));
INVX1 gate3473(.O (g4166), .I (I5568));
INVX1 gate3474(.O (g6516), .I (g6409));
INVX1 gate3475(.O (g5274), .I (I6933));
INVX1 gate3476(.O (I8435), .I (g6413));
INVX1 gate3477(.O (I3148), .I (g1595));
INVX1 gate3478(.O (I8690), .I (g6571));
INVX1 gate3479(.O (g1985), .I (I3096));
INVX1 gate3480(.O (I4334), .I (g2256));
INVX1 gate3481(.O (I8482), .I (g6461));
INVX1 gate3482(.O (g2739), .I (I3906));
INVX1 gate3483(.O (g3761), .I (g3605));
INVX1 gate3484(.O (I3155), .I (g1612));
INVX1 gate3485(.O (I3355), .I (g1608));
INVX1 gate3486(.O (I2402), .I (g774));
INVX1 gate3487(.O (g4529), .I (I6099));
INVX1 gate3488(.O (g1284), .I (g851));
INVX1 gate3489(.O (g4148), .I (I5526));
INVX1 gate3490(.O (I6733), .I (g4773));
INVX1 gate3491(.O (I8656), .I (g6532));
INVX1 gate3492(.O (g3830), .I (I5019));
INVX1 gate3493(.O (I9122), .I (g6864));
INVX1 gate3494(.O (g2079), .I (g1348));
INVX1 gate3495(.O (g4155), .I (I5551));
INVX1 gate3496(.O (g4851), .I (I6561));
INVX1 gate3497(.O (g6892), .I (I9143));
INVX1 gate3498(.O (g1832), .I (I2910));
INVX1 gate3499(.O (I9230), .I (g6936));
INVX1 gate3500(.O (g1853), .I (I2955));
INVX1 gate3501(.O (g2840), .I (g2538));
INVX1 gate3502(.O (I2877), .I (key_out_122));
INVX1 gate3503(.O (I5879), .I (g3745));
INVX1 gate3504(.O (g5544), .I (g5331));
INVX1 gate3505(.O (g2390), .I (I3531));
INVX1 gate3506(.O (I6324), .I (g4450));
INVX1 gate3507(.O (g1559), .I (g965));
INVX1 gate3508(.O (I6069), .I (g4213));
INVX1 gate3509(.O (I8110), .I (g6143));
INVX1 gate3510(.O (g4463), .I (g4364));
INVX1 gate3511(.O (g943), .I (g496));
INVX1 gate3512(.O (g1931), .I (I3034));
INVX1 gate3513(.O (g6709), .I (I8837));
INVX1 gate3514(.O (g3932), .I (I5169));
INVX1 gate3515(.O (I6540), .I (g4714));
INVX1 gate3516(.O (I3720), .I (g2155));
INVX1 gate3517(.O (g6078), .I (g5801));
INVX1 gate3518(.O (I1871), .I (g281));
INVX1 gate3519(.O (I6377), .I (g4569));
INVX1 gate3520(.O (g5061), .I (I6701));
INVX1 gate3521(.O (g6478), .I (I8342));
INVX1 gate3522(.O (I2464), .I (g850));
INVX1 gate3523(.O (I3367), .I (g1283));
INVX1 gate3524(.O (g5387), .I (I7051));
INVX1 gate3525(.O (I9137), .I (g6864));
INVX1 gate3526(.O (g1905), .I (I3004));
INVX1 gate3527(.O (I8002), .I (g6110));
INVX1 gate3528(.O (g866), .I (g314));
INVX1 gate3529(.O (I2785), .I (key_out_124));
INVX1 gate3530(.O (I7086), .I (g5281));
INVX1 gate3531(.O (I5615), .I (g3914));
INVX1 gate3532(.O (g6035), .I (g5824));
INVX1 gate3533(.O (g4720), .I (I6340));
INVX1 gate3534(.O (I3843), .I (g2145));
INVX1 gate3535(.O (g4118), .I (I5436));
INVX1 gate3536(.O (g4619), .I (g4248));
INVX1 gate3537(.O (g6517), .I (I8467));
INVX1 gate3538(.O (g1204), .I (g39));
INVX1 gate3539(.O (g3677), .I (g3140));
INVX1 gate3540(.O (g6876), .I (I9095));
INVX1 gate3541(.O (g4843), .I (I6537));
INVX1 gate3542(.O (g3866), .I (I5091));
INVX1 gate3543(.O (g2954), .I (g2381));
INVX1 gate3544(.O (I4593), .I (g2966));
INVX1 gate3545(.O (g5046), .I (I6680));
INVX1 gate3546(.O (g2163), .I (I3288));
INVX1 gate3547(.O (g6656), .I (I8764));
INVX1 gate3548(.O (g4193), .I (I5609));
INVX1 gate3549(.O (I2237), .I (g465));
INVX1 gate3550(.O (g2032), .I (g1749));
INVX1 gate3551(.O (g4393), .I (I5882));
INVX1 gate3552(.O (I5545), .I (g3814));
INVX1 gate3553(.O (g5403), .I (I7069));
INVX1 gate3554(.O (I1838), .I (g206));
INVX1 gate3555(.O (g3848), .I (I5059));
INVX1 gate3556(.O (I5591), .I (g3821));
INVX1 gate3557(.O (I4264), .I (g2212));
INVX1 gate3558(.O (I2394), .I (g719));
INVX1 gate3559(.O (g5391), .I (I7055));
INVX1 gate3560(.O (g2568), .I (I3678));
INVX1 gate3561(.O (I2731), .I (g1117));
INVX1 gate3562(.O (I4050), .I (g2059));
INVX1 gate3563(.O (g3241), .I (I4522));
INVX1 gate3564(.O (g2912), .I (g2001));
INVX1 gate3565(.O (g4121), .I (I5445));
INVX1 gate3566(.O (g1969), .I (I3080));
INVX1 gate3567(.O (I3232), .I (g1782));
INVX1 gate3568(.O (g4321), .I (I5790));
INVX1 gate3569(.O (g5307), .I (I6959));
INVX1 gate3570(.O (g2157), .I (I3278));
INVX1 gate3571(.O (g5536), .I (g5467));
INVX1 gate3572(.O (g2357), .I (I3509));
INVX1 gate3573(.O (g1123), .I (I2165));
INVX1 gate3574(.O (g1323), .I (I2324));
INVX1 gate3575(.O (g4625), .I (g4267));
INVX1 gate3576(.O (I3909), .I (g2044));
INVX1 gate3577(.O (g4232), .I (I5674));
INVX1 gate3578(.O (g6402), .I (I8220));
INVX1 gate3579(.O (g6824), .I (I9005));
INVX1 gate3580(.O (g1666), .I (g1088));
INVX1 gate3581(.O (g4938), .I (I6630));
INVX1 gate3582(.O (I6819), .I (g5019));
INVX1 gate3583(.O (g6236), .I (g6070));
INVX1 gate3584(.O (I3519), .I (g1305));
INVX1 gate3585(.O (I8295), .I (g6295));
INVX1 gate3586(.O (I2955), .I (g1729));
INVX1 gate3587(.O (I7487), .I (g5684));
INVX1 gate3588(.O (g856), .I (g654));
INVX1 gate3589(.O (I6923), .I (g5124));
INVX1 gate3590(.O (g1528), .I (g878));
INVX1 gate3591(.O (I5204), .I (g3534));
INVX1 gate3592(.O (I5630), .I (g3914));
INVX1 gate3593(.O (I6488), .I (g4603));
INVX1 gate3594(.O (g1351), .I (I2388));
INVX1 gate3595(.O (g1648), .I (I2623));
INVX1 gate3596(.O (I2814), .I (key_out_124));
INVX1 gate3597(.O (g1875), .I (I2970));
INVX1 gate3598(.O (g4519), .I (I6069));
INVX1 gate3599(.O (g5115), .I (I6759));
INVX1 gate3600(.O (g6590), .I (I8638));
INVX1 gate3601(.O (g5251), .I (g5069));
INVX1 gate3602(.O (g6877), .I (I9098));
INVX1 gate3603(.O (g3258), .I (I4537));
INVX1 gate3604(.O (I4777), .I (g2962));
INVX1 gate3605(.O (I6701), .I (g4726));
INVX1 gate3606(.O (g5315), .I (g5116));
INVX1 gate3607(.O (g3867), .I (I5094));
INVX1 gate3608(.O (I2150), .I (g10));
INVX1 gate3609(.O (g1655), .I (g985));
INVX1 gate3610(.O (g6657), .I (I8767));
INVX1 gate3611(.O (g4606), .I (g4193));
INVX1 gate3612(.O (I3687), .I (g1814));
INVX1 gate3613(.O (I8089), .I (g6120));
INVX1 gate3614(.O (I2773), .I (g1191));
INVX1 gate3615(.O (g5874), .I (I7634));
INVX1 gate3616(.O (g1410), .I (g1233));
INVX1 gate3617(.O (I8966), .I (g6796));
INVX1 gate3618(.O (I5750), .I (g4022));
INVX1 gate3619(.O (I7045), .I (g5167));
INVX1 gate3620(.O (I6114), .I (g4405));
INVX1 gate3621(.O (g3975), .I (I5249));
INVX1 gate3622(.O (I7173), .I (g5436));
INVX1 gate3623(.O (g1884), .I (I2979));
INVX1 gate3624(.O (I7091), .I (g5281));
INVX1 gate3625(.O (g6899), .I (I9164));
INVX1 gate3626(.O (I4799), .I (g2967));
INVX1 gate3627(.O (I2212), .I (g123));
INVX1 gate3628(.O (g929), .I (g49));
INVX1 gate3629(.O (g6785), .I (I8943));
INVX1 gate3630(.O (g5880), .I (g5824));
INVX1 gate3631(.O (I5040), .I (key_out_5));
INVX1 gate3632(.O (I2967), .I (g1682));
INVX1 gate3633(.O (g5537), .I (g5385));
INVX1 gate3634(.O (g2778), .I (g2391));
INVX1 gate3635(.O (I1862), .I (g278));
INVX1 gate3636(.O (I3525), .I (g1461));
INVX1 gate3637(.O (g3370), .I (g3124));
INVX1 gate3638(.O (g2894), .I (g1891));
INVX1 gate3639(.O (I7007), .I (g5314));
INVX1 gate3640(.O (g1372), .I (I2408));
INVX1 gate3641(.O (g4141), .I (I5505));
INVX1 gate3642(.O (g6563), .I (I8573));
INVX1 gate3643(.O (I6008), .I (g4163));
INVX1 gate3644(.O (I3691), .I (g1732));
INVX1 gate3645(.O (g4525), .I (I6087));
INVX1 gate3646(.O (g1143), .I (I2172));
INVX1 gate3647(.O (g3984), .I (key_out_1));
INVX1 gate3648(.O (I8150), .I (g6185));
INVX1 gate3649(.O (g1282), .I (g849));
INVX1 gate3650(.O (I8438), .I (g6416));
INVX1 gate3651(.O (g3083), .I (I4318));
INVX1 gate3652(.O (g1988), .I (I3099));
INVX1 gate3653(.O (I4802), .I (g2877));
INVX1 gate3654(.O (I6972), .I (g5135));
INVX1 gate3655(.O (g3483), .I (g2716));
INVX1 gate3656(.O (I7261), .I (g5458));
INVX1 gate3657(.O (g6194), .I (I7906));
INVX1 gate3658(.O (g1334), .I (I2355));
INVX1 gate3659(.O (I3158), .I (g1829));
INVX1 gate3660(.O (I3659), .I (g1491));
INVX1 gate3661(.O (I3358), .I (g1323));
INVX1 gate3662(.O (g5328), .I (I6986));
INVX1 gate3663(.O (I1927), .I (g665));
INVX1 gate3664(.O (g6489), .I (g6369));
INVX1 gate3665(.O (g5542), .I (g5331));
INVX1 gate3666(.O (g5330), .I (I6992));
INVX1 gate3667(.O (g3306), .I (g3057));
INVX1 gate3668(.O (g2998), .I (I4195));
INVX1 gate3669(.O (g4158), .I (I5556));
INVX1 gate3670(.O (g4659), .I (I6250));
INVX1 gate3671(.O (g1555), .I (I2521));
INVX1 gate3672(.O (g3790), .I (g3388));
INVX1 gate3673(.O (I3587), .I (g1461));
INVX1 gate3674(.O (g1792), .I (I2848));
INVX1 gate3675(.O (g2603), .I (I3733));
INVX1 gate3676(.O (g2039), .I (I3148));
INVX1 gate3677(.O (g3187), .I (I4424));
INVX1 gate3678(.O (g2484), .I (I3611));
INVX1 gate3679(.O (g3387), .I (I4664));
INVX1 gate3680(.O (g3461), .I (g2986));
INVX1 gate3681(.O (g4587), .I (g4215));
INVX1 gate3682(.O (I6033), .I (g4179));
INVX1 gate3683(.O (g5554), .I (g5455));
INVX1 gate3684(.O (g3622), .I (I4821));
INVX1 gate3685(.O (g4111), .I (I5415));
INVX1 gate3686(.O (I8229), .I (g6330));
INVX1 gate3687(.O (I9149), .I (g6884));
INVX1 gate3688(.O (I2620), .I (key_out_125));
INVX1 gate3689(.O (g1113), .I (I2147));
INVX1 gate3690(.O (I4492), .I (g3001));
INVX1 gate3691(.O (g4615), .I (g4322));
INVX1 gate3692(.O (g2583), .I (g1830));
INVX1 gate3693(.O (g3904), .I (g3575));
INVX1 gate3694(.O (g3200), .I (I4437));
INVX1 gate3695(.O (I6096), .I (g4397));
INVX1 gate3696(.O (g3046), .I (I4267));
INVX1 gate3697(.O (g899), .I (I1924));
INVX1 gate3698(.O (g4374), .I (I5837));
INVX1 gate3699(.O (I3284), .I (g1702));
INVX1 gate3700(.O (g2919), .I (g1937));
INVX1 gate3701(.O (g1908), .I (I3007));
INVX1 gate3702(.O (I2788), .I (key_out_120));
INVX1 gate3703(.O (g1094), .I (I2122));
INVX1 gate3704(.O (I5618), .I (g3821));
INVX1 gate3705(.O (g2952), .I (g2381));
INVX1 gate3706(.O (I6337), .I (g4455));
INVX1 gate3707(.O (I5343), .I (g3599));
INVX1 gate3708(.O (g2276), .I (I3425));
INVX1 gate3709(.O (g1567), .I (I2537));
INVX1 gate3710(.O (g4284), .I (I5739));
INVX1 gate3711(.O (g5512), .I (I7254));
INVX1 gate3712(.O (g4545), .I (g4416));
INVX1 gate3713(.O (g5090), .I (g4741));
INVX1 gate3714(.O (g6409), .I (g6285));
INVX1 gate3715(.O (g5490), .I (I7190));
INVX1 gate3716(.O (I7689), .I (g5708));
INVX1 gate3717(.O (g4380), .I (I5851));
INVX1 gate3718(.O (I2842), .I (key_out_125));
INVX1 gate3719(.O (g1776), .I (I2821));
INVX1 gate3720(.O (g1593), .I (g1054));
INVX1 gate3721(.O (g2004), .I (I3115));
INVX1 gate3722(.O (g4853), .I (I6567));
INVX1 gate3723(.O (g6836), .I (I9031));
INVX1 gate3724(.O (I2485), .I (g766));
INVX1 gate3725(.O (I3794), .I (g2044));
INVX1 gate3726(.O (g2986), .I (g2010));
INVX1 gate3727(.O (g4020), .I (I5324));
INVX1 gate3728(.O (g6212), .I (I7910));
INVX1 gate3729(.O (I5548), .I (g4059));
INVX1 gate3730(.O (g5456), .I (g5300));
INVX1 gate3731(.O (g2647), .I (I3791));
INVX1 gate3732(.O (I8837), .I (g6665));
INVX1 gate3733(.O (g5148), .I (I6812));
INVX1 gate3734(.O (g5649), .I (I7404));
INVX1 gate3735(.O (g4507), .I (I6033));
INVX1 gate3736(.O (g3223), .I (I4468));
INVX1 gate3737(.O (I4623), .I (g2962));
INVX1 gate3738(.O (I1947), .I (g699));
INVX1 gate3739(.O (g2764), .I (g2357));
INVX1 gate3740(.O (I8620), .I (g6541));
INVX1 gate3741(.O (I8462), .I (g6430));
INVX1 gate3742(.O (I9119), .I (g6855));
INVX1 gate3743(.O (I2854), .I (key_out_120));
INVX1 gate3744(.O (g4559), .I (g4187));
INVX1 gate3745(.O (g5155), .I (g5099));
INVX1 gate3746(.O (g5355), .I (I7007));
INVX1 gate3747(.O (I9152), .I (g6889));
INVX1 gate3748(.O (g3016), .I (I4223));
INVX1 gate3749(.O (g6229), .I (g6036));
INVX1 gate3750(.O (g1160), .I (I2179));
INVX1 gate3751(.O (g5260), .I (g4938));
INVX1 gate3752(.O (I6081), .I (g4388));
INVX1 gate3753(.O (I4375), .I (g2254));
INVX1 gate3754(.O (g6822), .I (g6786));
INVX1 gate3755(.O (g1641), .I (I2604));
INVX1 gate3756(.O (g3251), .I (I4534));
INVX1 gate3757(.O (I6692), .I (g4720));
INVX1 gate3758(.O (g1450), .I (I2453));
INVX1 gate3759(.O (g5063), .I (g4799));
INVX1 gate3760(.O (I7910), .I (g5905));
INVX1 gate3761(.O (I8249), .I (g6289));
INVX1 gate3762(.O (g4628), .I (g4273));
INVX1 gate3763(.O (g4515), .I (I6057));
INVX1 gate3764(.O (g2120), .I (I3251));
INVX1 gate3765(.O (I4285), .I (g2555));
INVX1 gate3766(.O (g2320), .I (I3474));
INVX1 gate3767(.O (g4100), .I (I5382));
INVX1 gate3768(.O (g1724), .I (I2724));
INVX1 gate3769(.O (g3874), .I (I5103));
INVX1 gate3770(.O (I2958), .I (g1257));
INVX1 gate3771(.O (I5094), .I (g3705));
INVX1 gate3772(.O (I2376), .I (g729));
INVX1 gate3773(.O (I8485), .I (g6479));
INVX1 gate3774(.O (g5720), .I (I7481));
INVX1 gate3775(.O (I2405), .I (g1112));
INVX1 gate3776(.O (g2906), .I (g1911));
INVX1 gate3777(.O (g2789), .I (g2410));
INVX1 gate3778(.O (g1878), .I (I2973));
INVX1 gate3779(.O (g5118), .I (I6766));
INVX1 gate3780(.O (I9170), .I (g6883));
INVX1 gate3781(.O (I1917), .I (g48));
AN2X1 gate3782(.O (g2771), .I1 (g2497), .I2 (g1975));
AN2X1 gate3783(.O (g6620), .I1 (g6516), .I2 (g6117));
AN2X1 gate3784(.O (g5193), .I1 (g532), .I2 (g4967));
AN4X1 gate3785(.O (I5360), .I1 (g3532), .I2 (g3536), .I3 (g3539), .I4 (g3544));
AN2X1 gate3786(.O (g5598), .I1 (g5046), .I2 (g5509));
AN2X1 gate3787(.O (g6249), .I1 (g1332), .I2 (g5892));
AN2X1 gate3788(.O (g4666), .I1 (g4630), .I2 (g4627));
AN2X1 gate3789(.O (g3629), .I1 (g2809), .I2 (g2738));
AN2X1 gate3790(.O (g3328), .I1 (g2701), .I2 (g1894));
AN2X1 gate3791(.O (g6085), .I1 (key_out_126), .I2 (g5731));
AN2X1 gate3792(.O (g4351), .I1 (g166), .I2 (g3776));
AN2X1 gate3793(.O (g4648), .I1 (g4407), .I2 (g79));
AN2X1 gate3794(.O (g5232), .I1 (g548), .I2 (g4980));
AN2X1 gate3795(.O (g2340), .I1 (g1398), .I2 (g1387));
AN2X1 gate3796(.O (g5938), .I1 (g5114), .I2 (g5791));
AN2X1 gate3797(.O (g5909), .I1 (g5787), .I2 (g3384));
AN2X1 gate3798(.O (g1802), .I1 (g89), .I2 (g1064));
AN2X1 gate3799(.O (g3554), .I1 (g2941), .I2 (g179));
AN2X1 gate3800(.O (g4410), .I1 (g3903), .I2 (g1474));
AN2X1 gate3801(.O (g6640), .I1 (g1612), .I2 (g6549));
AN2X1 gate3802(.O (g4172), .I1 (g3930), .I2 (g1366));
AN2X1 gate3803(.O (g4372), .I1 (g406), .I2 (g3790));
AN2X1 gate3804(.O (g3512), .I1 (g2928), .I2 (g1764));
AN2X1 gate3805(.O (g3490), .I1 (g353), .I2 (g2959));
AN2X1 gate3806(.O (g4667), .I1 (g4653), .I2 (g4651));
AN2X1 gate3807(.O (g3166), .I1 (g2042), .I2 (g1233));
AN2X1 gate3808(.O (g3366), .I1 (g248), .I2 (g2893));
AN2X1 gate3809(.O (g6829), .I1 (g6806), .I2 (g5958));
AN2X1 gate3810(.O (g3649), .I1 (g3104), .I2 (g2764));
AN2X1 gate3811(.O (g6911), .I1 (g6904), .I2 (g6902));
AN2X1 gate3812(.O (g3155), .I1 (g248), .I2 (g2461));
AN2X1 gate3813(.O (g3698), .I1 (g2284), .I2 (g2835));
AN2X1 gate3814(.O (g6270), .I1 (key_out_45), .I2 (g6062));
AN2X1 gate3815(.O (g4792), .I1 (g1417), .I2 (g4471));
AN3X1 gate3816(.O (g6473), .I1 (g2036), .I2 (g6397), .I3 (g1628));
AN2X1 gate3817(.O (g4621), .I1 (g3953), .I2 (g4364));
AN2X1 gate3818(.O (g5158), .I1 (g504), .I2 (g4993));
AN2X1 gate3819(.O (g6124), .I1 (g5705), .I2 (g5958));
AN2X1 gate3820(.O (g6324), .I1 (g3880), .I2 (g6212));
AN3X1 gate3821(.O (g6469), .I1 (g2121), .I2 (g2032), .I3 (g6394));
AN2X1 gate3822(.O (g3279), .I1 (g2599), .I2 (g2612));
AN2X1 gate3823(.O (g3619), .I1 (g2449), .I2 (g3057));
AN2X1 gate3824(.O (g3167), .I1 (g1883), .I2 (g921));
AN2X1 gate3825(.O (g5311), .I1 (g5013), .I2 (g4468));
AN2X1 gate3826(.O (g3367), .I1 (g2809), .I2 (g1960));
AN2X1 gate3827(.O (g3652), .I1 (g2544), .I2 (g3096));
AN3X1 gate3828(.O (g3843), .I1 (g2856), .I2 (g945), .I3 (g3533));
AN2X1 gate3829(.O (g4593), .I1 (g4277), .I2 (g947));
AN2X1 gate3830(.O (g3686), .I1 (g2256), .I2 (g2819));
AN2X1 gate3831(.O (g5180), .I1 (g414), .I2 (g4950));
AN2X1 gate3832(.O (g5380), .I1 (g188), .I2 (g5264));
AN2X1 gate3833(.O (g4160), .I1 (g3923), .I2 (g1345));
AN2X1 gate3834(.O (g3321), .I1 (g2252), .I2 (g2713));
AN2X1 gate3835(.O (g2089), .I1 (key_out_122), .I2 (g1578));
AN2X1 gate3836(.O (g6245), .I1 (g1329), .I2 (g5889));
AN2X1 gate3837(.O (g4360), .I1 (g184), .I2 (g3785));
AN2X1 gate3838(.O (g3670), .I1 (g2234), .I2 (g2792));
AN2X1 gate3839(.O (g3625), .I1 (g2619), .I2 (g2320));
AN2X1 gate3840(.O (g6291), .I1 (g5210), .I2 (g6161));
AN2X1 gate3841(.O (g4050), .I1 (I5359), .I2 (I5360));
AN2X1 gate3842(.O (g5559), .I1 (g5024), .I2 (g5453));
AN2X1 gate3843(.O (g6144), .I1 (g3183), .I2 (g5997));
AN2X1 gate3844(.O (g6344), .I1 (g6272), .I2 (g6080));
AN2X1 gate3845(.O (g2948), .I1 (g2137), .I2 (g1595));
AN2X1 gate3846(.O (g6259), .I1 (key_out_42), .I2 (g6044));
AN2X1 gate3847(.O (g4179), .I1 (g390), .I2 (g3902));
AN2X1 gate3848(.O (g2955), .I1 (g2381), .I2 (g297));
AN2X1 gate3849(.O (g6088), .I1 (key_out_123), .I2 (g5753));
AN2X1 gate3850(.O (g6852), .I1 (g6847), .I2 (g2295));
AN2X1 gate3851(.O (g6923), .I1 (g6918), .I2 (g6917));
AN2X1 gate3852(.O (g5515), .I1 (g590), .I2 (g5364));
AN2X1 gate3853(.O (g1499), .I1 (g1101), .I2 (g1094));
AN2X1 gate3854(.O (g4835), .I1 (g4533), .I2 (g4530));
AN2X1 gate3855(.O (g3687), .I1 (g2245), .I2 (g2820));
AN3X1 gate3856(.O (g4271), .I1 (g2121), .I2 (g1749), .I3 (g4004));
AN3X1 gate3857(.O (g4611), .I1 (g3985), .I2 (g119), .I3 (g4300));
AN2X1 gate3858(.O (g3341), .I1 (g2998), .I2 (g2709));
AN2X1 gate3859(.O (g6650), .I1 (g6580), .I2 (g6235));
AN2X1 gate3860(.O (g4541), .I1 (g631), .I2 (g4199));
AN2X1 gate3861(.O (g3645), .I1 (g2497), .I2 (g3090));
AN2X1 gate3862(.O (g5123), .I1 (g4670), .I2 (g1936));
AN2X1 gate3863(.O (g3691), .I1 (g2268), .I2 (g2828));
AN2X1 gate3864(.O (g4209), .I1 (g3816), .I2 (g865));
AN2X1 gate3865(.O (g4353), .I1 (g3989), .I2 (g3332));
AN2X1 gate3866(.O (g6336), .I1 (g6246), .I2 (g6065));
AN2X1 gate3867(.O (g6768), .I1 (g6750), .I2 (g3477));
AN2X1 gate3868(.O (g4744), .I1 (g3434), .I2 (g4582));
AN2X1 gate3869(.O (g3659), .I1 (g2672), .I2 (g2361));
AN2X1 gate3870(.O (g5351), .I1 (g5326), .I2 (g3459));
AN2X1 gate3871(.O (g3358), .I1 (g2842), .I2 (g1369));
AN2X1 gate3872(.O (g5648), .I1 (g4507), .I2 (g5545));
AN2X1 gate3873(.O (g6934), .I1 (g6932), .I2 (g3605));
AN2X1 gate3874(.O (g3275), .I1 (g2172), .I2 (g2615));
AN2X1 gate3875(.O (g3311), .I1 (g218), .I2 (g2872));
AN2X1 gate3876(.O (g5410), .I1 (g378), .I2 (g5274));
AN2X1 gate3877(.O (g3615), .I1 (g2422), .I2 (g3046));
AN2X1 gate3878(.O (g2062), .I1 (g1499), .I2 (g1666));
AN2X1 gate3879(.O (g3374), .I1 (g2809), .I2 (g1969));
AN2X1 gate3880(.O (g4600), .I1 (g4054), .I2 (g4289));
AN2X1 gate3881(.O (g6096), .I1 (key_out_127), .I2 (g5753));
AN2X1 gate3882(.O (g1436), .I1 (g834), .I2 (g830));
AN2X1 gate3883(.O (g5172), .I1 (g441), .I2 (g4877));
AN2X1 gate3884(.O (g3180), .I1 (g260), .I2 (g2506));
AN2X1 gate3885(.O (g5618), .I1 (g5506), .I2 (g4933));
AN2X1 gate3886(.O (g5143), .I1 (g157), .I2 (g5099));
AN2X1 gate3887(.O (g6913), .I1 (g6900), .I2 (g6898));
AN2X1 gate3888(.O (g5235), .I1 (g554), .I2 (g4980));
AN2X1 gate3889(.O (g4580), .I1 (g706), .I2 (g4262));
AN2X1 gate3890(.O (g2085), .I1 (key_out_122), .I2 (g1567));
AN2X1 gate3891(.O (g6266), .I1 (key_out_46), .I2 (g6057));
AN2X1 gate3892(.O (g5555), .I1 (g5014), .I2 (g5442));
AN2X1 gate3893(.O (g2941), .I1 (g2166), .I2 (g170));
AN2X1 gate3894(.O (g6248), .I1 (g465), .I2 (g5894));
AN2X1 gate3895(.O (g6342), .I1 (g6264), .I2 (g6076));
AN2X1 gate3896(.O (g5621), .I1 (g5508), .I2 (g4943));
AN2X1 gate3897(.O (g3628), .I1 (g2449), .I2 (g3070));
AN2X1 gate3898(.O (g6255), .I1 (g1335), .I2 (g5895));
AN2X1 gate3899(.O (g6081), .I1 (key_out_125), .I2 (g5731));
AN2X1 gate3900(.O (g3630), .I1 (g3167), .I2 (g1756));
AN2X1 gate3901(.O (g6692), .I1 (g6616), .I2 (g6615));
AN2X1 gate3902(.O (g3300), .I1 (g2232), .I2 (g2682));
AN2X1 gate3903(.O (g6154), .I1 (g3219), .I2 (g6015));
AN2X1 gate3904(.O (g6354), .I1 (g5866), .I2 (g6193));
AN2X1 gate3905(.O (g4184), .I1 (g3934), .I2 (g2136));
AN2X1 gate3906(.O (g5494), .I1 (g5443), .I2 (g3455));
AN2X1 gate3907(.O (g4384), .I1 (g414), .I2 (g3797));
AN2X1 gate3908(.O (g4339), .I1 (g3971), .I2 (g3289));
AN2X1 gate3909(.O (g4838), .I1 (g4648), .I2 (g84));
AN2X1 gate3910(.O (g3123), .I1 (g230), .I2 (g2391));
AN2X1 gate3911(.O (g3323), .I1 (g2253), .I2 (g2716));
AN2X1 gate3912(.O (g4672), .I1 (g4635), .I2 (g4631));
AN2X1 gate3913(.O (g2733), .I1 (g2422), .I2 (g1943));
AN2X1 gate3914(.O (g3666), .I1 (g3128), .I2 (g2787));
AN2X1 gate3915(.O (g6129), .I1 (g5717), .I2 (g5975));
AN2X1 gate3916(.O (g6329), .I1 (g3888), .I2 (g6212));
AN2X1 gate3917(.O (g2073), .I1 (g1088), .I2 (g1499));
AN2X1 gate3918(.O (g5360), .I1 (g4431), .I2 (g5160));
AN2X1 gate3919(.O (g6828), .I1 (g6803), .I2 (g5958));
AN2X1 gate3920(.O (g5050), .I1 (g4285), .I2 (g4807));
AN2X1 gate3921(.O (g3351), .I1 (g2760), .I2 (g1931));
AN2X1 gate3922(.O (g6830), .I1 (g6809), .I2 (g5975));
AN2X1 gate3923(.O (g3648), .I1 (g2722), .I2 (g2343));
AN2X1 gate3924(.O (g3655), .I1 (g2197), .I2 (g2768));
AN3X1 gate3925(.O (g1706), .I1 (g766), .I2 (g719), .I3 (g729));
AN2X1 gate3926(.O (g6068), .I1 (g5824), .I2 (key_out_45));
AN2X1 gate3927(.O (g4044), .I1 (g410), .I2 (g3388));
AN3X1 gate3928(.O (g6468), .I1 (g2032), .I2 (g6394), .I3 (g1609));
AN2X1 gate3929(.O (g3172), .I1 (g2449), .I2 (g2491));
AN2X1 gate3930(.O (g3278), .I1 (g2175), .I2 (g2628));
AN2X1 gate3931(.O (g3372), .I1 (g254), .I2 (g2905));
AN2X1 gate3932(.O (g2781), .I1 (g2544), .I2 (g1982));
AN2X1 gate3933(.O (g3618), .I1 (g3016), .I2 (g2712));
AN2X1 gate3934(.O (g3667), .I1 (g2245), .I2 (g2789));
AN2X1 gate3935(.O (g3143), .I1 (g242), .I2 (g2437));
AN2X1 gate3936(.O (g3282), .I1 (g131), .I2 (g2863));
AN2X1 gate3937(.O (g6716), .I1 (g6682), .I2 (g932));
AN2X1 gate3938(.O (g6149), .I1 (g3200), .I2 (g5997));
AN2X1 gate3939(.O (g3693), .I1 (g2256), .I2 (g2830));
AN2X1 gate3940(.O (g3134), .I1 (g230), .I2 (g2413));
AN2X1 gate3941(.O (g3334), .I1 (g236), .I2 (g2883));
AN3X1 gate3942(.O (g6848), .I1 (g3741), .I2 (g328), .I3 (g6843));
AN2X1 gate3943(.O (g5153), .I1 (g492), .I2 (g4904));
AN2X1 gate3944(.O (g5209), .I1 (g560), .I2 (key_out_89));
AN2X1 gate3945(.O (g5353), .I1 (g5327), .I2 (g3463));
AN2X1 gate3946(.O (g6241), .I1 (g1325), .I2 (g5887));
AN2X1 gate3947(.O (g1808), .I1 (g706), .I2 (g49));
AN2X1 gate3948(.O (g3113), .I1 (g224), .I2 (g2364));
AN2X1 gate3949(.O (g5558), .I1 (g5018), .I2 (g5450));
AN2X1 gate3950(.O (g6644), .I1 (g6575), .I2 (g6230));
AN2X1 gate3951(.O (g6152), .I1 (g3212), .I2 (g6015));
AN2X1 gate3952(.O (g6258), .I1 (g512), .I2 (g5899));
AN2X1 gate3953(.O (g4178), .I1 (g3959), .I2 (g2110));
AN2X1 gate3954(.O (g1575), .I1 (g980), .I2 (g965));
AN2X1 gate3955(.O (g4378), .I1 (g410), .I2 (g3792));
AN2X1 gate3956(.O (g4831), .I1 (g4528), .I2 (g4524));
AN2X1 gate3957(.O (g4182), .I1 (g394), .I2 (g3904));
AN2X1 gate3958(.O (g5492), .I1 (g5441), .I2 (g3452));
AN2X1 gate3959(.O (g5600), .I1 (g5502), .I2 (g4900));
AN2X1 gate3960(.O (g6614), .I1 (g932), .I2 (g6556));
AN2X1 gate3961(.O (g4947), .I1 (g184), .I2 (g4741));
AN2X1 gate3962(.O (g3360), .I1 (g2783), .I2 (g1947));
AN2X1 gate3963(.O (g6125), .I1 (g5708), .I2 (g5975));
AN2X1 gate3964(.O (g1419), .I1 (g613), .I2 (g918));
AN2X1 gate3965(.O (g3641), .I1 (g2644), .I2 (g2333));
AN2X1 gate3966(.O (g4873), .I1 (g4838), .I2 (g4173));
AN2X1 gate3967(.O (g4037), .I1 (g2896), .I2 (g3388));
AN2X1 gate3968(.O (g3724), .I1 (g117), .I2 (g3251));
AN2X1 gate3969(.O (g4495), .I1 (g3913), .I2 (g4292));
AN2X1 gate3970(.O (g3379), .I1 (g3104), .I2 (g1988));
AN2X1 gate3971(.O (g5175), .I1 (g5094), .I2 (g1384));
AN2X1 gate3972(.O (g3658), .I1 (g3118), .I2 (g2776));
AN2X1 gate3973(.O (g6061), .I1 (g5824), .I2 (key_out_43));
AN2X1 gate3974(.O (g5500), .I1 (g5430), .I2 (g5074));
AN2X1 gate3975(.O (g3611), .I1 (g2370), .I2 (g3037));
AN2X1 gate3976(.O (g2137), .I1 (g760), .I2 (g1638));
AN2X1 gate3977(.O (g4042), .I1 (g406), .I2 (g3388));
AN2X1 gate3978(.O (g5184), .I1 (g453), .I2 (g4877));
AN2X1 gate3979(.O (g4442), .I1 (g4239), .I2 (g2882));
AN2X1 gate3980(.O (g4164), .I1 (g3958), .I2 (g2091));
AN2X1 gate3981(.O (g2807), .I1 (g2568), .I2 (g2001));
AN2X1 gate3982(.O (g5424), .I1 (g390), .I2 (g5296));
AN2X1 gate3983(.O (g6145), .I1 (g3187), .I2 (g6015));
AN2X1 gate3984(.O (g2859), .I1 (g2112), .I2 (g1649));
AN3X1 gate3985(.O (g3997), .I1 (g1250), .I2 (g3425), .I3 (g2849));
AN2X1 gate3986(.O (g4054), .I1 (g3694), .I2 (g69));
AN2X1 gate3987(.O (g6345), .I1 (g6273), .I2 (g6083));
AN2X1 gate3988(.O (g3132), .I1 (g2306), .I2 (g1206));
AN2X1 gate3989(.O (g3680), .I1 (g2245), .I2 (g2805));
AN2X1 gate3990(.O (g6637), .I1 (g1842), .I2 (g6549));
AN2X1 gate3991(.O (g3353), .I1 (g3162), .I2 (g2921));
AN2X1 gate3992(.O (g2142), .I1 (g1793), .I2 (g1777));
AN2X1 gate3993(.O (g2255), .I1 (g1706), .I2 (g736));
AN2X1 gate3994(.O (g6159), .I1 (g3177), .I2 (g6015));
AN2X1 gate3995(.O (g2081), .I1 (g1094), .I2 (g1546));
AN2X1 gate3996(.O (g3558), .I1 (g338), .I2 (g3199));
AN2X1 gate3997(.O (g5499), .I1 (g5451), .I2 (g3462));
AN2X1 gate3998(.O (g4389), .I1 (g449), .I2 (g3798));
AN2X1 gate3999(.O (g4171), .I1 (g3956), .I2 (g2104));
AN2X1 gate4000(.O (g6315), .I1 (g3849), .I2 (g6194));
AN2X1 gate4001(.O (g4371), .I1 (g461), .I2 (g3789));
AN3X1 gate4002(.O (g4429), .I1 (g923), .I2 (g4253), .I3 (g2936));
AN2X1 gate4003(.O (g4787), .I1 (g2937), .I2 (g4628));
AN2X1 gate4004(.O (g6047), .I1 (g5824), .I2 (key_out_48));
AN2X1 gate4005(.O (g6874), .I1 (g6873), .I2 (g2060));
AN2X1 gate4006(.O (g2267), .I1 (g1716), .I2 (g791));
AN3X1 gate4007(.O (g5444), .I1 (g4545), .I2 (g5256), .I3 (g1574));
AN2X1 gate4008(.O (g5269), .I1 (g557), .I2 (key_out_89));
AN2X1 gate4009(.O (g1407), .I1 (g301), .I2 (g866));
AN2X1 gate4010(.O (g4684), .I1 (g4584), .I2 (g1341));
AN2X1 gate4011(.O (g4791), .I1 (g3936), .I2 (g4636));
AN2X1 gate4012(.O (g6243), .I1 (g500), .I2 (g5890));
AN2X1 gate4013(.O (g6935), .I1 (g6933), .I2 (g3622));
AN2X1 gate4014(.O (g2746), .I1 (g2473), .I2 (g1954));
AN2X1 gate4015(.O (g4759), .I1 (g536), .I2 (g4500));
AN2X1 gate4016(.O (g6128), .I1 (g5590), .I2 (g5958));
AN2X1 gate4017(.O (g5414), .I1 (g382), .I2 (g5278));
AN2X1 gate4018(.O (g6130), .I1 (g5720), .I2 (g5958));
AN2X1 gate4019(.O (g5660), .I1 (g4509), .I2 (g5549));
AN2X1 gate4020(.O (g3375), .I1 (g260), .I2 (g2912));
AN2X1 gate4021(.O (g4449), .I1 (g4266), .I2 (g2887));
AN2X1 gate4022(.O (g3651), .I1 (g3064), .I2 (g2766));
AN2X1 gate4023(.O (g4865), .I1 (g4776), .I2 (g1849));
AN2X1 gate4024(.O (g2953), .I1 (g2381), .I2 (g293));
AN2X1 gate4025(.O (g2068), .I1 (g1541), .I2 (g1546));
AN2X1 gate4026(.O (g3285), .I1 (g2195), .I2 (g2653));
AN2X1 gate4027(.O (g4833), .I1 (g4521), .I2 (g4516));
AN2X1 gate4028(.O (g5178), .I1 (g516), .I2 (g4993));
AN2X1 gate4029(.O (g5679), .I1 (g74), .I2 (g5576));
AN2X1 gate4030(.O (g5378), .I1 (g179), .I2 (g5260));
AN2X1 gate4031(.O (g3339), .I1 (g2734), .I2 (g1914));
AN2X1 gate4032(.O (g1689), .I1 (g766), .I2 (g719));
AN2X1 gate4033(.O (g5182), .I1 (g520), .I2 (g4993));
AN2X1 gate4034(.O (g2699), .I1 (g2397), .I2 (g1905));
AN2X1 gate4035(.O (g2747), .I1 (g2449), .I2 (g1957));
AN2X1 gate4036(.O (g6090), .I1 (key_out_126), .I2 (g5742));
AN2X1 gate4037(.O (g4362), .I1 (g3996), .I2 (g3355));
AN2X1 gate4038(.O (g3672), .I1 (g3136), .I2 (g2800));
AN2X1 gate4039(.O (g4052), .I1 (g418), .I2 (g3388));
AN2X1 gate4040(.O (g3643), .I1 (g2518), .I2 (g3086));
AN2X1 gate4041(.O (g4452), .I1 (g3820), .I2 (g4227));
AN2X1 gate4042(.O (g6056), .I1 (g5824), .I2 (key_out_42));
AN2X1 gate4043(.O (g1826), .I1 (g714), .I2 (g710));
AN2X1 gate4044(.O (g6148), .I1 (g3196), .I2 (g6015));
AN2X1 gate4045(.O (g6348), .I1 (g5869), .I2 (g6211));
AN2X1 gate4046(.O (g5560), .I1 (g5044), .I2 (g5456));
AN2X1 gate4047(.O (g3634), .I1 (g2179), .I2 (g2744));
AN2X1 gate4048(.O (g6155), .I1 (g2588), .I2 (g5997));
AN2X1 gate4049(.O (g6851), .I1 (g6846), .I2 (g2293));
AN2X1 gate4050(.O (g3551), .I1 (g2937), .I2 (g938));
AN2X1 gate4051(.O (g3099), .I1 (g218), .I2 (g2350));
AN2X1 gate4052(.O (g3304), .I1 (g2857), .I2 (g1513));
AN2X1 gate4053(.O (g4486), .I1 (g716), .I2 (g4195));
AN2X1 gate4054(.O (g3499), .I1 (g357), .I2 (g2961));
AN2X1 gate4055(.O (g4730), .I1 (g1423), .I2 (g4565));
AN2X1 gate4056(.O (g5632), .I1 (g4494), .I2 (g5538));
AN2X1 gate4057(.O (g5095), .I1 (g4794), .I2 (g951));
AN2X1 gate4058(.O (g6260), .I1 (key_out_41), .I2 (g6048));
AN2X1 gate4059(.O (g4185), .I1 (g398), .I2 (g3906));
AN2X1 gate4060(.O (g1609), .I1 (g760), .I2 (g754));
AN2X1 gate4061(.O (g5495), .I1 (g5444), .I2 (g3456));
AN4X1 gate4062(.O (g2577), .I1 (g1743), .I2 (g1797), .I3 (g1793), .I4 (g1138));
AN2X1 gate4063(.O (g3613), .I1 (g2604), .I2 (g2312));
AN2X1 gate4064(.O (g6619), .I1 (g6515), .I2 (g6115));
AN2X1 gate4065(.O (g6318), .I1 (g3865), .I2 (g6212));
AN4X1 gate4066(.O (g2026), .I1 (g1359), .I2 (g1402), .I3 (g1398), .I4 (g901));
AN2X1 gate4067(.O (g5164), .I1 (g437), .I2 (g4877));
AN2X1 gate4068(.O (g5364), .I1 (g574), .I2 (g5194));
AN2X1 gate4069(.O (g5233), .I1 (g551), .I2 (g4980));
AN2X1 gate4070(.O (g2821), .I1 (g1890), .I2 (g910));
AN2X1 gate4071(.O (g3729), .I1 (g327), .I2 (g3441));
AN2X1 gate4072(.O (g5454), .I1 (g5256), .I2 (g4549));
AN2X1 gate4073(.O (g5553), .I1 (g5012), .I2 (g5440));
AN2X1 gate4074(.O (g6321), .I1 (g3873), .I2 (g6212));
AN2X1 gate4075(.O (g3660), .I1 (g2568), .I2 (g3110));
AN3X1 gate4076(.O (g6625), .I1 (g2121), .I2 (g1595), .I3 (g6538));
AN2X1 gate4077(.O (g4045), .I1 (g3425), .I2 (g123));
AN2X1 gate4078(.O (g4445), .I1 (g4235), .I2 (g1854));
AN2X1 gate4079(.O (g6253), .I1 (g508), .I2 (g5896));
AN2X1 gate4080(.O (g4373), .I1 (g4001), .I2 (g3370));
AN2X1 gate4081(.O (g5189), .I1 (g528), .I2 (g4993));
AN2X1 gate4082(.O (g4491), .I1 (g3554), .I2 (g4215));
AN2X1 gate4083(.O (g6909), .I1 (g6896), .I2 (g6894));
AN2X1 gate4084(.O (g4169), .I1 (g3966), .I2 (g2099));
AN2X1 gate4085(.O (g5171), .I1 (g406), .I2 (g4950));
AN2X1 gate4086(.O (g4369), .I1 (g3999), .I2 (g3364));
AN2X1 gate4087(.O (g3679), .I1 (g2245), .I2 (g2803));
AN2X1 gate4088(.O (g4602), .I1 (g4407), .I2 (g4293));
AN2X1 gate4089(.O (g5371), .I1 (g152), .I2 (g5248));
AN2X1 gate4090(.O (g3378), .I1 (g3136), .I2 (g2932));
AN2X1 gate4091(.O (g5429), .I1 (g398), .I2 (g5304));
AN2X1 gate4092(.O (g4407), .I1 (g4054), .I2 (g74));
AN2X1 gate4093(.O (g5956), .I1 (g5783), .I2 (g5425));
AN2X1 gate4094(.O (g4868), .I1 (g4774), .I2 (g2891));
AN2X1 gate4095(.O (g5675), .I1 (g64), .I2 (g5574));
AN2X1 gate4096(.O (g3135), .I1 (g2370), .I2 (g2416));
AN2X1 gate4097(.O (g4459), .I1 (g4245), .I2 (g1899));
AN2X1 gate4098(.O (g3335), .I1 (g230), .I2 (g2884));
AN2X1 gate4099(.O (g3831), .I1 (g2330), .I2 (g3425));
AN2X1 gate4100(.O (g3182), .I1 (g2473), .I2 (g2512));
AN2X1 gate4101(.O (g3288), .I1 (g2631), .I2 (g2634));
AN2X1 gate4102(.O (g3382), .I1 (g3136), .I2 (g2934));
AN2X1 gate4103(.O (g4793), .I1 (g4277), .I2 (g4639));
AN2X1 gate4104(.O (g4015), .I1 (g445), .I2 (g3388));
AN2X1 gate4105(.O (g2107), .I1 (g1583), .I2 (g1543));
AN2X1 gate4106(.O (g6141), .I1 (g3173), .I2 (g5997));
AN2X1 gate4107(.O (g6341), .I1 (g6261), .I2 (g6074));
AN2X1 gate4108(.O (g6645), .I1 (g6576), .I2 (g6231));
AN2X1 gate4109(.O (g3632), .I1 (g3043), .I2 (g2743));
AN2X1 gate4110(.O (g3437), .I1 (g837), .I2 (g2853));
AN2X1 gate4111(.O (g3653), .I1 (g2215), .I2 (g2767));
AN2X1 gate4112(.O (g5201), .I1 (g4859), .I2 (g5084));
AN2X1 gate4113(.O (g3208), .I1 (g895), .I2 (g2551));
AN2X1 gate4114(.O (g3302), .I1 (g212), .I2 (g2867));
AN2X1 gate4115(.O (g6158), .I1 (g2594), .I2 (g6015));
AN2X1 gate4116(.O (g5449), .I1 (g4545), .I2 (g5246));
AN2X1 gate4117(.O (g5604), .I1 (g5059), .I2 (g5521));
AN2X1 gate4118(.O (g5098), .I1 (g4021), .I2 (g4837));
AN2X1 gate4119(.O (g5498), .I1 (g5449), .I2 (g3460));
AN2X1 gate4120(.O (g1585), .I1 (g1017), .I2 (g1011));
AN2X1 gate4121(.O (g6275), .I1 (key_out_47), .I2 (g6070));
AN2X1 gate4122(.O (g6311), .I1 (g3837), .I2 (g6194));
AN2X1 gate4123(.O (g4671), .I1 (g4645), .I2 (g4641));
AN3X1 gate4124(.O (g4247), .I1 (g1764), .I2 (g4007), .I3 (g1628));
AN2X1 gate4125(.O (g3454), .I1 (g2933), .I2 (g1660));
AN2X1 gate4126(.O (g4826), .I1 (g4209), .I2 (g4463));
AN2X1 gate4127(.O (g5162), .I1 (g5088), .I2 (g2105));
AN2X1 gate4128(.O (g5362), .I1 (g4437), .I2 (g5174));
AN2X1 gate4129(.O (g3296), .I1 (g3054), .I2 (g2650));
AN2X1 gate4130(.O (g5419), .I1 (g386), .I2 (g5292));
AN2X1 gate4131(.O (g3725), .I1 (g118), .I2 (g3251));
AN2X1 gate4132(.O (g2935), .I1 (g2291), .I2 (g1788));
AN2X1 gate4133(.O (g5452), .I1 (g5315), .I2 (g4612));
AN2X1 gate4134(.O (g6559), .I1 (g1612), .I2 (g6474));
AN2X1 gate4135(.O (g5728), .I1 (g5623), .I2 (g3889));
AN2X1 gate4136(.O (g5486), .I1 (g386), .I2 (g5331));
AN2X1 gate4137(.O (g5185), .I1 (g524), .I2 (g4993));
AN2X1 gate4138(.O (g3171), .I1 (g248), .I2 (g2488));
AN2X1 gate4139(.O (g3371), .I1 (g260), .I2 (g2904));
AN3X1 gate4140(.O (g6628), .I1 (g2138), .I2 (g1612), .I3 (g6540));
AN2X1 gate4141(.O (g4165), .I1 (g3927), .I2 (g1352));
AN2X1 gate4142(.O (g4048), .I1 (g414), .I2 (g3388));
AN2X1 gate4143(.O (g4448), .I1 (g3815), .I2 (g4225));
AN2X1 gate4144(.O (g3281), .I1 (g2178), .I2 (g2640));
AN2X1 gate4145(.O (g4827), .I1 (g4520), .I2 (g4515));
AN2X1 gate4146(.O (g4333), .I1 (g3964), .I2 (g3284));
AN3X1 gate4147(.O (I2566), .I1 (g749), .I2 (g743), .I3 (g736));
AN2X1 gate4148(.O (g2166), .I1 (g1633), .I2 (g161));
AN2X1 gate4149(.O (g3684), .I1 (g2268), .I2 (g2817));
AN2X1 gate4150(.O (g4396), .I1 (g422), .I2 (g3801));
AN2X1 gate4151(.O (g3338), .I1 (g3162), .I2 (g2914));
AN2X1 gate4152(.O (g2056), .I1 (g1672), .I2 (g1675));
AN2X1 gate4153(.O (g5406), .I1 (g374), .I2 (g5270));
AN2X1 gate4154(.O (g3309), .I1 (g2243), .I2 (g2695));
AN2X1 gate4155(.O (g5635), .I1 (g4498), .I2 (g5542));
AN2X1 gate4156(.O (g5682), .I1 (g84), .I2 (g5578));
AN2X1 gate4157(.O (g5487), .I1 (g390), .I2 (g5331));
AN2X1 gate4158(.O (g6123), .I1 (g5702), .I2 (g5958));
AN2X1 gate4159(.O (g6323), .I1 (g3877), .I2 (g6194));
AN2X1 gate4160(.O (g3759), .I1 (g2644), .I2 (g3498));
AN2X1 gate4161(.O (g5226), .I1 (g672), .I2 (g5054));
AN2X1 gate4162(.O (g6151), .I1 (g3209), .I2 (g5997));
AN2X1 gate4163(.O (g3449), .I1 (g128), .I2 (g2946));
AN2X1 gate4164(.O (g6648), .I1 (g6579), .I2 (g6234));
AN2X1 gate4165(.O (g5173), .I1 (g512), .I2 (g4993));
AN2X1 gate4166(.O (g5373), .I1 (g161), .I2 (g5250));
AN2X1 gate4167(.O (g4181), .I1 (g3939), .I2 (g1381));
AN2X1 gate4168(.O (g2720), .I1 (g2422), .I2 (g1919));
AN2X1 gate4169(.O (g4685), .I1 (g4591), .I2 (g2079));
AN2X1 gate4170(.O (g5169), .I1 (g5093), .I2 (g1375));
AN2X1 gate4171(.O (g5369), .I1 (g143), .I2 (g5247));
AN2X1 gate4172(.O (g5602), .I1 (g594), .I2 (g5515));
AN4X1 gate4173(.O (g2834), .I1 (g1263), .I2 (g1257), .I3 (g1270), .I4 (I4040));
AN2X1 gate4174(.O (g3362), .I1 (g3031), .I2 (g2740));
AN2X1 gate4175(.O (g6343), .I1 (g6268), .I2 (g6078));
AN2X1 gate4176(.O (g2121), .I1 (g1632), .I2 (g754));
AN2X1 gate4177(.O (g2670), .I1 (g2029), .I2 (g1503));
AN2X1 gate4178(.O (g6693), .I1 (g6618), .I2 (g6617));
AN2X1 gate4179(.O (g1633), .I1 (g716), .I2 (g152));
AN2X1 gate4180(.O (g6334), .I1 (g3858), .I2 (g6212));
AN2X1 gate4181(.O (g3728), .I1 (g326), .I2 (g3441));
AN2X1 gate4182(.O (g6555), .I1 (g1838), .I2 (g6469));
AN2X1 gate4183(.O (g3730), .I1 (g328), .I2 (g3441));
AN2X1 gate4184(.O (g2909), .I1 (g606), .I2 (g2092));
AN2X1 gate4185(.O (g4041), .I1 (g461), .I2 (g3388));
AN2X1 gate4186(.O (g3425), .I1 (g2296), .I2 (g3208));
AN2X1 gate4187(.O (g6313), .I1 (g3841), .I2 (g6194));
AN2X1 gate4188(.O (g5940), .I1 (g5115), .I2 (g5794));
AN2X1 gate4189(.O (g4673), .I1 (g4656), .I2 (g4654));
AN2X1 gate4190(.O (g5188), .I1 (g1043), .I2 (g4894));
AN2X1 gate4191(.O (g6908), .I1 (g6907), .I2 (g3886));
AN2X1 gate4192(.O (g5216), .I1 (g563), .I2 (key_out_89));
AN2X1 gate4193(.O (g6094), .I1 (key_out_125), .I2 (g5753));
AN2X1 gate4194(.O (g4168), .I1 (g3925), .I2 (g1355));
AN2X1 gate4195(.O (g4368), .I1 (g3998), .I2 (g3363));
AN2X1 gate4196(.O (g5671), .I1 (g54), .I2 (g5572));
AN2X1 gate4197(.O (g3678), .I1 (g2256), .I2 (g2802));
AN2X1 gate4198(.O (g5428), .I1 (g394), .I2 (g5300));
AN2X1 gate4199(.O (g4058), .I1 (g3424), .I2 (g1246));
AN2X1 gate4200(.O (g3635), .I1 (g2473), .I2 (g3079));
AN2X1 gate4201(.O (g2860), .I1 (g710), .I2 (g2296));
AN2X1 gate4202(.O (g3682), .I1 (g2772), .I2 (g2430));
AN2X1 gate4203(.O (g3305), .I1 (g2960), .I2 (g2296));
AN2X1 gate4204(.O (g5910), .I1 (g5816), .I2 (g5667));
AN2X1 gate4205(.O (g3755), .I1 (g2604), .I2 (g3481));
AN2X1 gate4206(.O (g2659), .I1 (g1686), .I2 (g2296));
AN2X1 gate4207(.O (g5883), .I1 (g5824), .I2 (g3752));
AN2X1 gate4208(.O (g3373), .I1 (g3118), .I2 (g2927));
AN2X1 gate4209(.O (g5217), .I1 (g4866), .I2 (g5092));
AN2X1 gate4210(.O (g4863), .I1 (g4777), .I2 (g2874));
AN2X1 gate4211(.O (g3283), .I1 (g2609), .I2 (g2622));
AN2X1 gate4212(.O (g3602), .I1 (g2688), .I2 (g2663));
AN3X1 gate4213(.O (I2574), .I1 (g804), .I2 (g798), .I3 (g791));
AN2X1 gate4214(.O (g5165), .I1 (g508), .I2 (g4993));
AN2X1 gate4215(.O (g6777), .I1 (g6762), .I2 (g3488));
AN3X1 gate4216(.O (g3718), .I1 (g1743), .I2 (g3140), .I3 (g1157));
AN2X1 gate4217(.O (g3767), .I1 (g2706), .I2 (g3504));
AN2X1 gate4218(.O (g4688), .I1 (g1474), .I2 (g4568));
AN2X1 gate4219(.O (g1784), .I1 (g858), .I2 (g889));
AN2X1 gate4220(.O (g2853), .I1 (g836), .I2 (g2021));
AN2X1 gate4221(.O (g6799), .I1 (g4948), .I2 (g6782));
AN2X1 gate4222(.O (g2794), .I1 (g2544), .I2 (g1994));
AN2X1 gate4223(.O (g3203), .I1 (g2497), .I2 (g2565));
AN2X1 gate4224(.O (g6132), .I1 (g3752), .I2 (g5880));
AN2X1 gate4225(.O (g6238), .I1 (g528), .I2 (g5886));
AN2X1 gate4226(.O (g6153), .I1 (g3216), .I2 (g5997));
AN2X1 gate4227(.O (g4183), .I1 (g3965), .I2 (g1391));
AN2X1 gate4228(.O (g4383), .I1 (g453), .I2 (g3796));
AN2X1 gate4229(.O (g6558), .I1 (g1842), .I2 (g6474));
AN2X1 gate4230(.O (g5181), .I1 (g449), .I2 (g4877));
AN2X1 gate4231(.O (g3689), .I1 (g3162), .I2 (g2826));
AN2X1 gate4232(.O (g4588), .I1 (g2419), .I2 (g4273));
AN2X1 gate4233(.O (g5197), .I1 (g465), .I2 (g4967));
AN2X1 gate4234(.O (g4161), .I1 (g3931), .I2 (g2087));
AN2X1 gate4235(.O (g4361), .I1 (g3995), .I2 (g3354));
AN2X1 gate4236(.O (g3671), .I1 (g2760), .I2 (g2405));
AN2X1 gate4237(.O (g4051), .I1 (g449), .I2 (g3388));
AN2X1 gate4238(.O (g6092), .I1 (key_out_122), .I2 (g5731));
AN2X1 gate4239(.O (g4346), .I1 (g157), .I2 (g3773));
AN2X1 gate4240(.O (g2323), .I1 (g471), .I2 (g1358));
AN2X1 gate4241(.O (g5562), .I1 (g5228), .I2 (g5457));
AN2X1 gate4242(.O (g3910), .I1 (key_out_3), .I2 (g1049));
AN2X1 gate4243(.O (g3609), .I1 (g2706), .I2 (g2678));
AN2X1 gate4244(.O (g6262), .I1 (g516), .I2 (g5901));
AN3X1 gate4245(.O (g6736), .I1 (g6712), .I2 (g754), .I3 (g5237));
AN2X1 gate4246(.O (g3758), .I1 (g545), .I2 (g3461));
AN2X1 gate4247(.O (g4043), .I1 (g457), .I2 (g3388));
AN2X1 gate4248(.O (g3365), .I1 (g254), .I2 (g2892));
AN3X1 gate4249(.O (g5441), .I1 (g4537), .I2 (g5251), .I3 (g1558));
AN2X1 gate4250(.O (g5673), .I1 (g59), .I2 (g5573));
AN2X1 gate4251(.O (g4347), .I1 (g3986), .I2 (g3320));
AN2X1 gate4252(.O (g3133), .I1 (g236), .I2 (g2410));
AN2X1 gate4253(.O (g3333), .I1 (g2264), .I2 (g2728));
AN2X1 gate4254(.O (g3774), .I1 (g3016), .I2 (g3510));
AN2X1 gate4255(.O (g4697), .I1 (g4589), .I2 (g1363));
AN2X1 gate4256(.O (g3780), .I1 (g3043), .I2 (g3519));
AN3X1 gate4257(.O (g6737), .I1 (g6714), .I2 (g760), .I3 (g5237));
AN2X1 gate4258(.O (g6077), .I1 (g5824), .I2 (key_out_47));
AN2X1 gate4259(.O (g3662), .I1 (g2544), .I2 (g3114));
AN2X1 gate4260(.O (g6643), .I1 (g6574), .I2 (g6229));
AN2X1 gate4261(.O (g3290), .I1 (g2213), .I2 (g2664));
AN2X1 gate4262(.O (g6634), .I1 (g1595), .I2 (g6545));
AN2X1 gate4263(.O (g3816), .I1 (g3434), .I2 (g861));
AN2X1 gate4264(.O (g2113), .I1 (g1576), .I2 (g1535));
AN2X1 gate4265(.O (g6099), .I1 (key_out_124), .I2 (g5753));
AN2X1 gate4266(.O (g6304), .I1 (g5915), .I2 (g6165));
AN2X1 gate4267(.O (g3181), .I1 (g254), .I2 (g2509));
AN2X1 gate4268(.O (g3381), .I1 (g3128), .I2 (g1998));
AN2X1 gate4269(.O (g3685), .I1 (g2256), .I2 (g2818));
AN2X1 gate4270(.O (g3700), .I1 (g2276), .I2 (g2837));
AN2X1 gate4271(.O (g3421), .I1 (g622), .I2 (g2846));
AN2X1 gate4272(.O (g5569), .I1 (g5348), .I2 (g3772));
AN2X1 gate4273(.O (g4460), .I1 (g4218), .I2 (g1539));
AN2X1 gate4274(.O (g4597), .I1 (g3694), .I2 (g4286));
AN2X1 gate4275(.O (g6613), .I1 (g932), .I2 (g6554));
AN2X1 gate4276(.O (g4739), .I1 (g2850), .I2 (g4579));
AN2X1 gate4277(.O (g6269), .I1 (g524), .I2 (g5908));
AN2X1 gate4278(.O (g4937), .I1 (g166), .I2 (g4732));
AN2X1 gate4279(.O (g4668), .I1 (g4642), .I2 (g4638));
AN2X1 gate4280(.O (g3631), .I1 (g2631), .I2 (g2324));
AN2X1 gate4281(.O (g2160), .I1 (g1624), .I2 (g929));
AN2X1 gate4282(.O (g4390), .I1 (g418), .I2 (g3799));
AN2X1 gate4283(.O (g3301), .I1 (g218), .I2 (g2866));
AN2X1 gate4284(.O (g4501), .I1 (g4250), .I2 (g1671));
AN2X1 gate4285(.O (g4156), .I1 (g3926), .I2 (g2078));
AN2X1 gate4286(.O (g4356), .I1 (g175), .I2 (g3779));
AN2X1 gate4287(.O (g4942), .I1 (g175), .I2 (g4736));
AN2X1 gate4288(.O (g5183), .I1 (g418), .I2 (g4950));
AN2X1 gate4289(.O (g4163), .I1 (g374), .I2 (g3892));
AN2X1 gate4290(.O (g5023), .I1 (g3935), .I2 (g4804));
AN2X1 gate4291(.O (g4363), .I1 (g402), .I2 (g3786));
AN2X1 gate4292(.O (g4032), .I1 (g441), .I2 (g3388));
AN2X1 gate4293(.O (g4053), .I1 (g3387), .I2 (g1415));
AN2X1 gate4294(.O (g4453), .I1 (g4238), .I2 (g1858));
AN2X1 gate4295(.O (g5161), .I1 (g5095), .I2 (g4535));
AN2X1 gate4296(.O (g3669), .I1 (g2234), .I2 (g2790));
AN2X1 gate4297(.O (g5361), .I1 (g4435), .I2 (g5168));
AN2X1 gate4298(.O (g3368), .I1 (g2822), .I2 (g2923));
AN2X1 gate4299(.O (g6135), .I1 (g5584), .I2 (g5958));
AN2X1 gate4300(.O (g5665), .I1 (g361), .I2 (g5570));
AN2X1 gate4301(.O (g6831), .I1 (g6812), .I2 (g5975));
AN2X1 gate4302(.O (g5451), .I1 (g5251), .I2 (g4544));
AN2X1 gate4303(.O (g6288), .I1 (g5615), .I2 (g6160));
AN2X1 gate4304(.O (g4157), .I1 (g3830), .I2 (g1533));
AN2X1 gate4305(.O (g4357), .I1 (g3990), .I2 (g3342));
AN2X1 gate4306(.O (g5146), .I1 (g184), .I2 (g5099));
AN2X1 gate4307(.O (g6916), .I1 (g6903), .I2 (g6901));
AN2X1 gate4308(.O (g5633), .I1 (g4496), .I2 (g5539));
AN2X1 gate4309(.O (g3505), .I1 (g2924), .I2 (g1749));
AN2X1 gate4310(.O (g6749), .I1 (g6735), .I2 (g6734));
AN2X1 gate4311(.O (g6798), .I1 (g4946), .I2 (g6781));
AN2X1 gate4312(.O (g5944), .I1 (g5778), .I2 (g5403));
AN2X1 gate4313(.O (g5240), .I1 (g293), .I2 (g4915));
AN2X1 gate4314(.O (g5043), .I1 (g3941), .I2 (g4805));
AN3X1 gate4315(.O (g5443), .I1 (g4537), .I2 (g5251), .I3 (g2307));
AN2X1 gate4316(.O (g6302), .I1 (g5740), .I2 (g6164));
AN2X1 gate4317(.O (g6719), .I1 (g4518), .I2 (g6665));
AN2X1 gate4318(.O (g2092), .I1 (g642), .I2 (g1570));
AN2X1 gate4319(.O (g4683), .I1 (g4585), .I2 (g2066));
AN2X1 gate4320(.O (g5681), .I1 (g79), .I2 (g5577));
AN2X1 gate4321(.O (g3688), .I1 (g2783), .I2 (g2457));
AN2X1 gate4322(.O (g4735), .I1 (g2018), .I2 (g4577));
AN2X1 gate4323(.O (g6265), .I1 (g520), .I2 (g5903));
AN2X1 gate4324(.O (g4782), .I1 (g1624), .I2 (g4623));
AN2X1 gate4325(.O (g4661), .I1 (g4637), .I2 (g4634));
AN2X1 gate4326(.O (g4949), .I1 (g193), .I2 (g4753));
AN2X1 gate4327(.O (g3326), .I1 (g2734), .I2 (g1891));
AN2X1 gate4328(.O (g6770), .I1 (g6754), .I2 (g3482));
AN2X1 gate4329(.O (g3760), .I1 (g548), .I2 (g3465));
AN2X1 gate4330(.O (g5936), .I1 (g5113), .I2 (g5788));
AN2X1 gate4331(.O (g4039), .I1 (g402), .I2 (g3388));
AN2X1 gate4332(.O (g5317), .I1 (g148), .I2 (g4869));
AN2X1 gate4333(.O (g3383), .I1 (g3128), .I2 (g2004));
AN2X1 gate4334(.O (g5601), .I1 (g5052), .I2 (g5518));
AN2X1 gate4335(.O (g3608), .I1 (g2599), .I2 (g2308));
AN2X1 gate4336(.O (g3924), .I1 (g3505), .I2 (g471));
AN2X1 gate4337(.O (g4583), .I1 (g1808), .I2 (g4267));
AN2X1 gate4338(.O (g3161), .I1 (g2397), .I2 (g2470));
AN2X1 gate4339(.O (g2339), .I1 (g1603), .I2 (g197));
AN2X1 gate4340(.O (g3361), .I1 (g3150), .I2 (g1950));
AN2X1 gate4341(.O (g4616), .I1 (g4231), .I2 (g3761));
AN2X1 gate4342(.O (g3665), .I1 (g2748), .I2 (g2378));
AN2X1 gate4343(.O (g3127), .I1 (g224), .I2 (g2394));
AN2X1 gate4344(.O (g3327), .I1 (g2772), .I2 (g2906));
AN2X1 gate4345(.O (g3146), .I1 (g2370), .I2 (g2446));
AN2X1 gate4346(.O (g3633), .I1 (g2497), .I2 (g3076));
AN2X1 gate4347(.O (g5937), .I1 (g5775), .I2 (g5392));
AN2X1 gate4348(.O (g3103), .I1 (g212), .I2 (g2353));
AN2X1 gate4349(.O (g3303), .I1 (g2722), .I2 (g2890));
AN2X1 gate4350(.O (g5668), .I1 (g49), .I2 (g5571));
AN2X1 gate4351(.O (g6338), .I1 (g6251), .I2 (g6067));
AN2X1 gate4352(.O (g5190), .I1 (g426), .I2 (g4950));
AN2X1 gate4353(.O (g5501), .I1 (g5454), .I2 (g3478));
AN2X1 gate4354(.O (g2551), .I1 (g715), .I2 (g1826));
AN2X1 gate4355(.O (g5156), .I1 (g434), .I2 (g4877));
AN2X1 gate4356(.O (g5356), .I1 (g5265), .I2 (g1902));
AN2X1 gate4357(.O (g4277), .I1 (g3936), .I2 (g942));
AN2X1 gate4358(.O (g5942), .I1 (g5117), .I2 (g5797));
AN2X1 gate4359(.O (g4789), .I1 (g3551), .I2 (g4632));
AN2X1 gate4360(.O (g3316), .I1 (g2748), .I2 (g2894));
AN2X1 gate4361(.O (g3434), .I1 (g2850), .I2 (g857));
AN2X1 gate4362(.O (g5954), .I1 (g5121), .I2 (g5813));
AN2X1 gate4363(.O (g5163), .I1 (g402), .I2 (g4950));
AN2X1 gate4364(.O (g6098), .I1 (key_out_128), .I2 (g5753));
AN2X1 gate4365(.O (g3147), .I1 (g2419), .I2 (g59));
AN2X1 gate4366(.O (g5363), .I1 (g4439), .I2 (g5179));
AN2X1 gate4367(.O (g3681), .I1 (g2234), .I2 (g2806));
AN2X1 gate4368(.O (g5053), .I1 (g4599), .I2 (g4808));
AN2X1 gate4369(.O (g3697), .I1 (g2796), .I2 (g2481));
AN2X1 gate4370(.O (g5157), .I1 (g496), .I2 (g4904));
AN2X1 gate4371(.O (g5357), .I1 (g398), .I2 (g5220));
AN3X1 gate4372(.O (g4244), .I1 (g1749), .I2 (g4004), .I3 (g1609));
AN2X1 gate4373(.O (g4340), .I1 (g3972), .I2 (g3291));
AN2X1 gate4374(.O (g3936), .I1 (g3551), .I2 (g940));
AN2X1 gate4375(.O (g3117), .I1 (g218), .I2 (g2367));
AN2X1 gate4376(.O (g3317), .I1 (g2722), .I2 (g2895));
AN2X1 gate4377(.O (g4035), .I1 (g437), .I2 (g3388));
AN2X1 gate4378(.O (g918), .I1 (g610), .I2 (g602));
AN2X1 gate4379(.O (g6086), .I1 (key_out_123), .I2 (g5742));
AN2X1 gate4380(.O (g4214), .I1 (g1822), .I2 (g4045));
AN2X1 gate4381(.O (g1620), .I1 (g1056), .I2 (g1084));
AN2X1 gate4382(.O (g3784), .I1 (g114), .I2 (g3251));
AN2X1 gate4383(.O (g2916), .I1 (g1030), .I2 (g2113));
AN2X1 gate4384(.O (g3479), .I1 (g345), .I2 (g2957));
AN2X1 gate4385(.O (g6131), .I1 (g5593), .I2 (g5975));
AN2X1 gate4386(.O (g3668), .I1 (g2568), .I2 (g3124));
AN2X1 gate4387(.O (g6331), .I1 (g3891), .I2 (g6212));
AN2X1 gate4388(.O (g4236), .I1 (g654), .I2 (g3907));
AN2X1 gate4389(.O (g3294), .I1 (g139), .I2 (g2870));
AN2X1 gate4390(.O (g5949), .I1 (g5119), .I2 (g5805));
AN2X1 gate4391(.O (g3190), .I1 (g260), .I2 (g2535));
AN2X1 gate4392(.O (g6766), .I1 (g6750), .I2 (g2986));
AN2X1 gate4393(.O (g3156), .I1 (g242), .I2 (g2464));
AN2X1 gate4394(.O (g3356), .I1 (g248), .I2 (g2888));
AN2X1 gate4395(.O (g5646), .I1 (g4502), .I2 (g5544));
AN2X1 gate4396(.O (g2873), .I1 (g1845), .I2 (g1861));
AN2X1 gate4397(.O (g6748), .I1 (g6733), .I2 (g6732));
AN2X1 gate4398(.O (g5603), .I1 (g5504), .I2 (g4911));
AN2X1 gate4399(.O (g5484), .I1 (g378), .I2 (g5331));
AN2X1 gate4400(.O (g4928), .I1 (g148), .I2 (g4723));
AN2X1 gate4401(.O (g3704), .I1 (g2276), .I2 (g2841));
AN2X1 gate4402(.O (g4464), .I1 (g4272), .I2 (g1937));
AN2X1 gate4403(.O (g4785), .I1 (g2160), .I2 (g4625));
AN2X1 gate4404(.O (g6091), .I1 (key_out_126), .I2 (g5753));
AN2X1 gate4405(.O (g3810), .I1 (g625), .I2 (g3421));
AN2X1 gate4406(.O (g5952), .I1 (g5120), .I2 (g5809));
AN2X1 gate4407(.O (g5616), .I1 (g5505), .I2 (g4929));
AN2X1 gate4408(.O (g6718), .I1 (g4511), .I2 (g6661));
AN2X1 gate4409(.O (g6767), .I1 (g6754), .I2 (g2986));
AN2X1 gate4410(.O (g3157), .I1 (g2422), .I2 (g2467));
AN2X1 gate4411(.O (g3357), .I1 (g242), .I2 (g2889));
AN2X1 gate4412(.O (g4489), .I1 (g2166), .I2 (g4206));
AN2X1 gate4413(.O (g2770), .I1 (g2518), .I2 (g1972));
AN2X1 gate4414(.O (g4471), .I1 (g4253), .I2 (g332));
AN2X1 gate4415(.O (g5503), .I1 (g366), .I2 (g5384));
AN2X1 gate4416(.O (g3626), .I1 (g3031), .I2 (g2727));
AN2X1 gate4417(.O (g4038), .I1 (g430), .I2 (g3388));
AN2X1 gate4418(.O (g5617), .I1 (g5061), .I2 (g5524));
AN2X1 gate4419(.O (g3683), .I1 (g3150), .I2 (g2813));
AN2X1 gate4420(.O (g4836), .I1 (g4527), .I2 (g4523));
AN2X1 gate4421(.O (g2138), .I1 (g1639), .I2 (g809));
AN2X1 gate4422(.O (g3661), .I1 (g2234), .I2 (g2778));
AN2X1 gate4423(.O (g6247), .I1 (g504), .I2 (g5893));
AN2X1 gate4424(.O (g3627), .I1 (g2473), .I2 (g3067));
AN2X1 gate4425(.O (g5945), .I1 (g5118), .I2 (g5801));
AN2X1 gate4426(.O (g2808), .I1 (g2009), .I2 (g1581));
AN2X1 gate4427(.O (g3292), .I1 (g2214), .I2 (g2667));
AN2X1 gate4428(.O (g3646), .I1 (g2179), .I2 (g2756));
AN2X1 gate4429(.O (g2759), .I1 (g2473), .I2 (g1966));
AN2X1 gate4430(.O (g6910), .I1 (g6892), .I2 (g6891));
AN2X1 gate4431(.O (g3603), .I1 (g2370), .I2 (g3019));
AN2X1 gate4432(.O (g3484), .I1 (g349), .I2 (g2958));
AN2X1 gate4433(.O (g5482), .I1 (g370), .I2 (g5331));
AN2X1 gate4434(.O (g3702), .I1 (g2284), .I2 (g2839));
AN2X1 gate4435(.O (g6066), .I1 (g5824), .I2 (key_out_46));
AN2X1 gate4436(.O (g5214), .I1 (g562), .I2 (key_out_89));
AN2X1 gate4437(.O (g3616), .I1 (g2397), .I2 (g3049));
AN2X1 gate4438(.O (g6055), .I1 (g5824), .I2 (key_out_44));
AN2X1 gate4439(.O (g6133), .I1 (g5723), .I2 (g5975));
AN2X1 gate4440(.O (g5663), .I1 (g4513), .I2 (g5550));
AN2X1 gate4441(.O (g6333), .I1 (g3896), .I2 (g6212));
AN2X1 gate4442(.O (g2419), .I1 (g1808), .I2 (g54));
AN2X1 gate4443(.O (g3764), .I1 (g551), .I2 (g3480));
AN2X1 gate4444(.O (g5402), .I1 (g370), .I2 (g5266));
AN2X1 gate4445(.O (g5236), .I1 (g269), .I2 (g4915));
AN2X1 gate4446(.O (g4708), .I1 (g578), .I2 (g4541));
AN2X1 gate4447(.O (g5556), .I1 (g5015), .I2 (g5445));
AN2X1 gate4448(.O (g4219), .I1 (g3911), .I2 (g1655));
AN2X1 gate4449(.O (g3277), .I1 (g2174), .I2 (g2625));
AN2X1 gate4450(.O (g3617), .I1 (g2609), .I2 (g2317));
AN2X1 gate4451(.O (g6093), .I1 (key_out_125), .I2 (g5742));
AN2X1 gate4452(.O (g2897), .I1 (g1030), .I2 (g2062));
AN2X1 gate4453(.O (g6256), .I1 (key_out_44), .I2 (g6040));
AN2X1 gate4454(.O (g4176), .I1 (g386), .I2 (g3901));
AN2X1 gate4455(.O (g6816), .I1 (g6784), .I2 (g3346));
AN2X1 gate4456(.O (g4829), .I1 (g4526), .I2 (g4522));
AN2X1 gate4457(.O (g6263), .I1 (key_out_43), .I2 (g6052));
AN2X1 gate4458(.O (g5194), .I1 (g586), .I2 (g4874));
AN2X1 gate4459(.O (g3709), .I1 (g2284), .I2 (g2845));
AN2X1 gate4460(.O (g5557), .I1 (g5016), .I2 (g5448));
AN2X1 gate4461(.O (g3340), .I1 (g2772), .I2 (g2915));
AN2X1 gate4462(.O (g6631), .I1 (g1838), .I2 (g6545));
AN2X1 gate4463(.O (g3907), .I1 (g650), .I2 (g3522));
AN2X1 gate4464(.O (g4177), .I1 (g3933), .I2 (g1372));
AN2X1 gate4465(.O (g5948), .I1 (g5779), .I2 (g5407));
AN2X1 gate4466(.O (g4377), .I1 (g457), .I2 (g3791));
AN2X1 gate4467(.O (g3690), .I1 (g2276), .I2 (g2827));
AN2X1 gate4468(.O (g5955), .I1 (g5782), .I2 (g5420));
AN2X1 gate4469(.O (g5350), .I1 (g5325), .I2 (g3453));
AN2X1 gate4470(.O (g4199), .I1 (g628), .I2 (g3810));
AN2X1 gate4471(.O (g5438), .I1 (g5224), .I2 (g3769));
AN2X1 gate4472(.O (g2868), .I1 (g1316), .I2 (g1861));
AN2X1 gate4473(.O (g3310), .I1 (g224), .I2 (g2871));
AN2X1 gate4474(.O (g4797), .I1 (g4593), .I2 (g4643));
AN2X1 gate4475(.O (g5212), .I1 (g561), .I2 (key_out_89));
AN2X1 gate4476(.O (g3663), .I1 (g2215), .I2 (g2779));
AN2X1 gate4477(.O (g2793), .I1 (g2568), .I2 (g1991));
AN2X1 gate4478(.O (g2015), .I1 (g616), .I2 (g1419));
AN2X1 gate4479(.O (g4344), .I1 (g3981), .I2 (g3306));
AN2X1 gate4480(.O (g5229), .I1 (g545), .I2 (g4980));
AN2X1 gate4481(.O (g6772), .I1 (g6746), .I2 (g3312));
AN2X1 gate4482(.O (g3762), .I1 (g2672), .I2 (g3500));
AN2X1 gate4483(.O (g4694), .I1 (g1481), .I2 (g4578));
AN2X1 gate4484(.O (g3657), .I1 (g2734), .I2 (g2357));
AN2X1 gate4485(.O (g2721), .I1 (g2397), .I2 (g1922));
AN2X1 gate4486(.O (g4488), .I1 (g1633), .I2 (g4202));
AN2X1 gate4487(.O (g4701), .I1 (g4596), .I2 (g1378));
AN2X1 gate4488(.O (g3928), .I1 (g3512), .I2 (g478));
AN3X1 gate4489(.O (g6474), .I1 (g2138), .I2 (g2036), .I3 (g6397));
AN2X1 gate4490(.O (g3899), .I1 (g323), .I2 (g3441));
AN2X1 gate4491(.O (g3464), .I1 (g341), .I2 (g2956));
AN2X1 gate4492(.O (g5620), .I1 (g5507), .I2 (g4938));
AN2X1 gate4493(.O (g4870), .I1 (g4779), .I2 (g1884));
AN2X1 gate4494(.O (g3295), .I1 (g2660), .I2 (g2647));
AN2X1 gate4495(.O (g2671), .I1 (g2263), .I2 (g2296));
AN2X1 gate4496(.O (g1576), .I1 (g1101), .I2 (g1094));
AN2X1 gate4497(.O (g3844), .I1 (g3540), .I2 (g1665));
AN3X1 gate4498(.O (g1716), .I1 (g821), .I2 (g774), .I3 (g784));
AN2X1 gate4499(.O (g3089), .I1 (g212), .I2 (g2336));
AN2X1 gate4500(.O (g3731), .I1 (g331), .I2 (g3441));
AN2X1 gate4501(.O (g3489), .I1 (g2607), .I2 (g1861));
AN2X1 gate4502(.O (g5192), .I1 (g1046), .I2 (g4894));
AN2X1 gate4503(.O (g5485), .I1 (g382), .I2 (g5331));
AN2X1 gate4504(.O (g5941), .I1 (g5777), .I2 (g5399));
AN2X1 gate4505(.O (g4230), .I1 (g3756), .I2 (g1861));
AN2X1 gate4506(.O (g6126), .I1 (g5711), .I2 (g5958));
AN2X1 gate4507(.O (g6326), .I1 (g3833), .I2 (g6194));
AN2X1 gate4508(.O (g4033), .I1 (g426), .I2 (g3388));
AN2X1 gate4509(.O (g3814), .I1 (g913), .I2 (key_out_3));
AN2X1 gate4510(.O (g2758), .I1 (g2497), .I2 (g1963));
AN2X1 gate4511(.O (g3350), .I1 (g3150), .I2 (g1928));
AN2X1 gate4512(.O (g2861), .I1 (g2120), .I2 (g1654));
AN2X1 gate4513(.O (g6924), .I1 (g6920), .I2 (g6919));
AN2X1 gate4514(.O (g5176), .I1 (g410), .I2 (g4950));
AN2X1 gate4515(.O (g4395), .I1 (g445), .I2 (g3800));
AN2X1 gate4516(.O (g5376), .I1 (g170), .I2 (g5255));
AN2X1 gate4517(.O (g5911), .I1 (g5817), .I2 (g5670));
AN2X1 gate4518(.O (g2846), .I1 (g619), .I2 (g2015));
AN2X1 gate4519(.O (g6127), .I1 (g5714), .I2 (g5975));
AN2X1 gate4520(.O (g6327), .I1 (g3884), .I2 (g6212));
AN2X1 gate4521(.O (g5225), .I1 (g669), .I2 (g5054));
AN2X1 gate4522(.O (g4342), .I1 (g3978), .I2 (g3299));
AN2X1 gate4523(.O (g6146), .I1 (g3192), .I2 (g5997));
AN2X1 gate4524(.O (g6346), .I1 (g6274), .I2 (g6087));
AN2X1 gate4525(.O (g2018), .I1 (g1423), .I2 (g1254));
AN2X1 gate4526(.O (g4354), .I1 (g437), .I2 (g3777));
AN4X1 gate4527(.O (I5352), .I1 (g3529), .I2 (g3531), .I3 (g3535), .I4 (g3538));
AN2X1 gate4528(.O (g5177), .I1 (g445), .I2 (g4877));
AN2X1 gate4529(.O (g6240), .I1 (g4205), .I2 (g5888));
AN2X1 gate4530(.O (g3620), .I1 (g2422), .I2 (g3060));
AN2X1 gate4531(.O (g1027), .I1 (g598), .I2 (key_out_32));
AN2X1 gate4532(.O (g2685), .I1 (g2370), .I2 (g1887));
AN2X1 gate4533(.O (g2700), .I1 (g2370), .I2 (g1908));
AN2X1 gate4534(.O (g2021), .I1 (g835), .I2 (g1436));
AN2X1 gate4535(.O (g6316), .I1 (g3855), .I2 (g6194));
AN2X1 gate4536(.O (g5898), .I1 (g5800), .I2 (g5647));
AN2X1 gate4537(.O (g4401), .I1 (g426), .I2 (g3802));
AN2X1 gate4538(.O (g1514), .I1 (g1017), .I2 (g1011));
AN2X1 gate4539(.O (g5900), .I1 (g5804), .I2 (g5658));
AN2X1 gate4540(.O (g2950), .I1 (g2156), .I2 (g1612));
AN2X1 gate4541(.O (g4761), .I1 (g4567), .I2 (g1674));
AN2X1 gate4542(.O (g5245), .I1 (g297), .I2 (g4915));
AN2X1 gate4543(.O (g1763), .I1 (g478), .I2 (g1119));
AN2X1 gate4544(.O (g4828), .I1 (g4510), .I2 (g4508));
AN2X1 gate4545(.O (g3298), .I1 (g2231), .I2 (g2679));
AN2X1 gate4546(.O (g4830), .I1 (g4529), .I2 (g4525));
AN2X1 gate4547(.O (g5144), .I1 (g166), .I2 (g5099));
AN2X1 gate4548(.O (g4592), .I1 (g3147), .I2 (g4281));
AN2X1 gate4549(.O (g6914), .I1 (g6895), .I2 (g6893));
AN2X1 gate4550(.O (g2101), .I1 (g1001), .I2 (g1543));
AN2X1 gate4551(.O (g5488), .I1 (g394), .I2 (g5331));
AN2X1 gate4552(.O (g4932), .I1 (g157), .I2 (g4727));
AN2X1 gate4553(.O (g1416), .I1 (g913), .I2 (g266));
AN2X1 gate4554(.O (g5701), .I1 (g5683), .I2 (g3813));
AN2X1 gate4555(.O (g6317), .I1 (g3862), .I2 (g6194));
AN2X1 gate4556(.O (g5215), .I1 (g4864), .I2 (g5090));
AN2X1 gate4557(.O (g5951), .I1 (g5780), .I2 (g5411));
AN2X1 gate4558(.O (g4677), .I1 (g4652), .I2 (g4646));
AN2X1 gate4559(.O (g3176), .I1 (g2422), .I2 (g2494));
AN2X1 gate4560(.O (g3376), .I1 (g3104), .I2 (g1979));
AN2X1 gate4561(.O (g3286), .I1 (g2196), .I2 (g2656));
AN2X1 gate4562(.O (g3765), .I1 (g554), .I2 (g3485));
AN2X1 gate4563(.O (g4349), .I1 (g441), .I2 (g3775));
AN2X1 gate4564(.O (g6060), .I1 (g5824), .I2 (key_out_41));
AN4X1 gate4565(.O (g1595), .I1 (g729), .I2 (g719), .I3 (g766), .I4 (I2566));
AN4X1 gate4566(.O (I5359), .I1 (g3518), .I2 (g3521), .I3 (g3526), .I4 (g3530));
AN2X1 gate4567(.O (g3610), .I1 (g2397), .I2 (g3034));
AN3X1 gate4568(.O (g6739), .I1 (g6715), .I2 (g815), .I3 (g5242));
AN4X1 gate4569(.O (g1612), .I1 (g784), .I2 (g774), .I3 (g821), .I4 (I2574));
AN2X1 gate4570(.O (g3324), .I1 (g230), .I2 (g2875));
AN2X1 gate4571(.O (g6079), .I1 (key_out_120), .I2 (g5753));
AN2X1 gate4572(.O (g5122), .I1 (g193), .I2 (g4662));
AN2X1 gate4573(.O (g3377), .I1 (g3118), .I2 (g2931));
AN2X1 gate4574(.O (g4352), .I1 (g3988), .I2 (g3331));
AN2X1 gate4575(.O (g4867), .I1 (g4811), .I2 (g3872));
AN2X1 gate4576(.O (g6156), .I1 (g2591), .I2 (g6015));
AN2X1 gate4577(.O (g3287), .I1 (g135), .I2 (g2865));
AN2X1 gate4578(.O (g5096), .I1 (g4794), .I2 (g4647));
AN2X1 gate4579(.O (g4186), .I1 (g3973), .I2 (g1395));
AN2X1 gate4580(.O (g5496), .I1 (g5446), .I2 (g3457));
AN2X1 gate4581(.O (g6250), .I1 (key_out_48), .I2 (g6036));
AN2X1 gate4582(.O (g4170), .I1 (g382), .I2 (g3900));
AN3X1 gate4583(.O (g4280), .I1 (g2138), .I2 (g1764), .I3 (g4007));
AN2X1 gate4584(.O (g3144), .I1 (g236), .I2 (g2440));
AN2X1 gate4585(.O (g3344), .I1 (g242), .I2 (g2885));
AN2X1 gate4586(.O (g5142), .I1 (g148), .I2 (g5099));
AN2X1 gate4587(.O (g3819), .I1 (g964), .I2 (g3437));
AN2X1 gate4588(.O (g6912), .I1 (g6899), .I2 (g6897));
AN2X1 gate4589(.O (g3694), .I1 (g3147), .I2 (g64));
AN2X1 gate4590(.O (g6157), .I1 (g3158), .I2 (g5997));
AN2X1 gate4591(.O (g5481), .I1 (g366), .I2 (g5331));
AN2X1 gate4592(.O (g3701), .I1 (g2268), .I2 (g2838));
AN2X1 gate4593(.O (g5497), .I1 (g5447), .I2 (g3458));
AN2X1 gate4594(.O (g5154), .I1 (g500), .I2 (g4993));
AN2X1 gate4595(.O (g5354), .I1 (g5249), .I2 (g2903));
AN2X1 gate4596(.O (g4461), .I1 (g4241), .I2 (g2919));
AN2X1 gate4597(.O (g4756), .I1 (g3816), .I2 (g4587));
AN2X1 gate4598(.O (g4046), .I1 (I5351), .I2 (I5352));
AN2X1 gate4599(.O (g5218), .I1 (key_out_12), .I2 (key_out_89));
AN2X1 gate4600(.O (g3650), .I1 (g2660), .I2 (g2347));
AN2X1 gate4601(.O (g4345), .I1 (g3982), .I2 (g3308));
AN2X1 gate4602(.O (g3336), .I1 (g2760), .I2 (g1911));
AN2X1 gate4603(.O (g3768), .I1 (g3448), .I2 (g1528));
AN2X1 gate4604(.O (g4159), .I1 (g370), .I2 (g3890));
AN2X1 gate4605(.O (g4359), .I1 (g434), .I2 (g3782));
AN2X1 gate4606(.O (g3806), .I1 (g3384), .I2 (g2024));
AN2X1 gate4607(.O (g4416), .I1 (g3905), .I2 (g1481));
AN2X1 gate4608(.O (g3887), .I1 (g3276), .I2 (g1861));
AN2X1 gate4609(.O (g3122), .I1 (g2435), .I2 (g1394));
AN2X1 gate4610(.O (g2732), .I1 (g2449), .I2 (g1940));
AN2X1 gate4611(.O (g4047), .I1 (g453), .I2 (g3388));
AN2X1 gate4612(.O (g6646), .I1 (g6577), .I2 (g6232));
AN3X1 gate4613(.O (g3433), .I1 (g1359), .I2 (g2831), .I3 (g905));
AN2X1 gate4614(.O (g5953), .I1 (g5781), .I2 (g5415));
AN2X1 gate4615(.O (g6084), .I1 (key_out_122), .I2 (g5753));
AN2X1 gate4616(.O (g6603), .I1 (g6581), .I2 (g6236));
AN2X1 gate4617(.O (g4874), .I1 (g582), .I2 (g4708));
AN2X1 gate4618(.O (g5677), .I1 (g69), .I2 (g5575));
AN2X1 gate4619(.O (g3195), .I1 (g2473), .I2 (g2541));
AN2X1 gate4620(.O (g3337), .I1 (g2796), .I2 (g2913));
AN3X1 gate4621(.O (I4040), .I1 (g1279), .I2 (g2025), .I3 (g1267));
AN2X1 gate4622(.O (g5149), .I1 (g4910), .I2 (g1480));
AN2X1 gate4623(.O (g5349), .I1 (g5324), .I2 (g3451));
AN2X1 gate4624(.O (g5198), .I1 (g558), .I2 (key_out_89));
AN2X1 gate4625(.O (g5398), .I1 (g366), .I2 (g5261));
AN2X1 gate4626(.O (g1570), .I1 (g634), .I2 (g1027));
AN2X1 gate4627(.O (g6647), .I1 (g6578), .I2 (g6233));
AN2X1 gate4628(.O (g1691), .I1 (g821), .I2 (g774));
AN2X1 gate4629(.O (g3692), .I1 (g2268), .I2 (g2829));
AN2X1 gate4630(.O (g3726), .I1 (g119), .I2 (g3251));
AN2X1 gate4631(.O (g3154), .I1 (g2039), .I2 (g1410));
AN2X1 gate4632(.O (g4800), .I1 (g4648), .I2 (g4296));
AN2X1 gate4633(.O (g5152), .I1 (g430), .I2 (g4950));
AN2X1 gate4634(.O (g6320), .I1 (g3869), .I2 (g6194));
AN2X1 gate4635(.O (g5211), .I1 (g4860), .I2 (g5086));
AN2X1 gate4636(.O (g5186), .I1 (g422), .I2 (g4950));
AN2X1 gate4637(.O (g5599), .I1 (g5049), .I2 (g5512));
AN2X1 gate4638(.O (g4490), .I1 (g2941), .I2 (g4210));
AN2X1 gate4639(.O (g3293), .I1 (g212), .I2 (g2864));
AN2X1 gate4640(.O (g6771), .I1 (g6758), .I2 (g3483));
AN2X1 gate4641(.O (g3329), .I1 (g2748), .I2 (g2907));
AN2X1 gate4642(.O (g5170), .I1 (g5091), .I2 (g2111));
AN2X1 gate4643(.O (g4456), .I1 (g3829), .I2 (g4229));
AN2X1 gate4644(.O (g6299), .I1 (g5530), .I2 (g6163));
AN2X1 gate4645(.O (g4348), .I1 (g3987), .I2 (g3322));
AN2X1 gate4646(.O (g3727), .I1 (g122), .I2 (g3251));
AN2X1 gate4647(.O (g2937), .I1 (g2160), .I2 (g931));
AN2X1 gate4648(.O (g4355), .I1 (g430), .I2 (g3778));
AN2X1 gate4649(.O (g5939), .I1 (g5776), .I2 (g5395));
AN3X1 gate4650(.O (g2294), .I1 (g1716), .I2 (g791), .I3 (g798));
AN2X1 gate4651(.O (g4698), .I1 (g4586), .I2 (g2106));
AN2X1 gate4652(.O (g5483), .I1 (g374), .I2 (g5331));
AN2X1 gate4653(.O (g3703), .I1 (g2284), .I2 (g2840));
AN3X1 gate4654(.O (g6738), .I1 (g6713), .I2 (g809), .I3 (g5242));
AN2X1 gate4655(.O (g2156), .I1 (g815), .I2 (g1642));
AN2X1 gate4656(.O (g6244), .I1 (g4759), .I2 (g5891));
AN2X1 gate4657(.O (g2356), .I1 (g1603), .I2 (g269));
AN2X1 gate4658(.O (g6140), .I1 (g5587), .I2 (g5975));
AN2X1 gate4659(.O (g3953), .I1 (g3554), .I2 (g188));
AN2X1 gate4660(.O (g6340), .I1 (g6257), .I2 (g6069));
AN2X1 gate4661(.O (g5187), .I1 (g457), .I2 (g4877));
AN2X1 gate4662(.O (g1628), .I1 (g815), .I2 (g809));
AN2X1 gate4663(.O (g4167), .I1 (g378), .I2 (g3898));
AN2X1 gate4664(.O (g6082), .I1 (key_out_122), .I2 (g5742));
AN2X1 gate4665(.O (g4367), .I1 (g193), .I2 (g3788));
AN2X1 gate4666(.O (g4872), .I1 (g4760), .I2 (g1549));
AN2X1 gate4667(.O (g4057), .I1 (g422), .I2 (g3388));
AN2X1 gate4668(.O (g5904), .I1 (g5812), .I2 (g5664));
AN2X1 gate4669(.O (g5200), .I1 (g559), .I2 (key_out_89));
AN2X1 gate4670(.O (g4457), .I1 (g4261), .I2 (g2902));
AN2X1 gate4671(.O (g5446), .I1 (g4537), .I2 (g5241));
AN2X1 gate4672(.O (g3349), .I1 (g2783), .I2 (g1925));
AN2X1 gate4673(.O (g2053), .I1 (g1094), .I2 (g1675));
AN2X1 gate4674(.O (g5145), .I1 (g175), .I2 (g5099));
AN2X1 gate4675(.O (g6915), .I1 (g6906), .I2 (g6905));
AN2X1 gate4676(.O (g4834), .I1 (g4534), .I2 (g4531));
AN2X1 gate4677(.O (g4686), .I1 (g4590), .I2 (g1348));
AN2X1 gate4678(.O (g5191), .I1 (g461), .I2 (g4877));
AN2X1 gate4679(.O (g3699), .I1 (g2276), .I2 (g2836));
AN2X1 gate4680(.O (g4598), .I1 (g1978), .I2 (g4253));
AN2X1 gate4681(.O (g5637), .I1 (g4499), .I2 (g5543));
AN2X1 gate4682(.O (g5159), .I1 (g536), .I2 (g4967));
AN2X1 gate4683(.O (g5359), .I1 (g4428), .I2 (g5155));
AN2X1 gate4684(.O (g4253), .I1 (g1861), .I2 (g3819));
AN2X1 gate4685(.O (g3644), .I1 (g2197), .I2 (g2755));
AN2X1 gate4686(.O (g3319), .I1 (g2688), .I2 (g2675));
AN2X1 gate4687(.O (g3352), .I1 (g2796), .I2 (g2920));
AN2X1 gate4688(.O (g5047), .I1 (g3954), .I2 (g4806));
AN3X1 gate4689(.O (g5447), .I1 (g4545), .I2 (g5256), .I3 (g2311));
AN2X1 gate4690(.O (g4687), .I1 (g4493), .I2 (g1542));
AN2X1 gate4691(.O (g3186), .I1 (g2449), .I2 (g2515));
AN2X1 gate4692(.O (g3170), .I1 (g254), .I2 (g2485));
AN2X1 gate4693(.O (g3614), .I1 (g2998), .I2 (g2691));
AN2X1 gate4694(.O (g3325), .I1 (g224), .I2 (g2876));
AN2X1 gate4695(.O (g4341), .I1 (g3977), .I2 (g3297));
AN2X1 gate4696(.O (g2782), .I1 (g2518), .I2 (g1985));
AN2X1 gate4697(.O (g6295), .I1 (g5379), .I2 (g6162));
AN2X1 gate4698(.O (g3280), .I1 (g2177), .I2 (g2637));
AN2X1 gate4699(.O (g5017), .I1 (g4784), .I2 (g1679));
AN2X1 gate4700(.O (g4691), .I1 (g4581), .I2 (g2098));
AN2X1 gate4701(.O (g5935), .I1 (g5112), .I2 (g5784));
AN2X1 gate4702(.O (g2949), .I1 (g830), .I2 (g1861));
AN4X1 gate4703(.O (I5351), .I1 (g3511), .I2 (g3517), .I3 (g3520), .I4 (g3525));
AN2X1 gate4704(.O (g5234), .I1 (g197), .I2 (g4915));
AN2X1 gate4705(.O (g3636), .I1 (g2701), .I2 (g2327));
AN3X1 gate4706(.O (g2292), .I1 (g1706), .I2 (g736), .I3 (g743));
AN2X1 gate4707(.O (g6089), .I1 (key_out_123), .I2 (g5731));
AN2X1 gate4708(.O (g6731), .I1 (g6717), .I2 (g4427));
AN2X1 gate4709(.O (g6557), .I1 (g1595), .I2 (g6469));
AN2X1 gate4710(.O (g4358), .I1 (g3991), .I2 (g3343));
AN2X1 gate4711(.O (g2084), .I1 (g1577), .I2 (g1563));
AN2X1 gate4712(.O (g2850), .I1 (g2018), .I2 (g1255));
AN2X1 gate4713(.O (g5213), .I1 (g4862), .I2 (g5087));
AN2X1 gate4714(.O (g6254), .I1 (g532), .I2 (g5897));
AN2X1 gate4715(.O (g6150), .I1 (g3204), .I2 (g6015));
AN2X1 gate4716(.O (g5902), .I1 (g5808), .I2 (g5661));
AN2X1 gate4717(.O (g3145), .I1 (g2397), .I2 (g2443));
AN2X1 gate4718(.O (g3345), .I1 (g236), .I2 (g2886));
AN2X1 gate4719(.O (g6773), .I1 (g6762), .I2 (g2986));
AN2X1 gate4720(.O (g3763), .I1 (g3064), .I2 (g3501));
AN2X1 gate4721(.O (g3191), .I1 (g2497), .I2 (g2538));
AN2X1 gate4722(.O (g4180), .I1 (g3929), .I2 (g2119));
AN2X1 gate4723(.O (g5166), .I1 (g541), .I2 (g4967));
AN2X1 gate4724(.O (g3637), .I1 (g2822), .I2 (g2752));
AN2X1 gate4725(.O (g4832), .I1 (g4517), .I2 (g4512));
AN2X1 gate4726(.O (g6769), .I1 (g6758), .I2 (g2986));
AN2X1 gate4727(.O (g3307), .I1 (g2242), .I2 (g2692));
AN2X1 gate4728(.O (g3359), .I1 (g2822), .I2 (g2922));
AN2X1 gate4729(.O (g4794), .I1 (g4593), .I2 (g949));
AN2X1 gate4730(.O (g3757), .I1 (g2619), .I2 (g3487));
AN2X1 gate4731(.O (g3522), .I1 (g646), .I2 (g2909));
AN2X1 gate4732(.O (g3315), .I1 (g2701), .I2 (g1875));
AN2X1 gate4733(.O (g3642), .I1 (g3054), .I2 (g2754));
AN2X1 gate4734(.O (g3654), .I1 (g2518), .I2 (g3100));
AN2X1 gate4735(.O (g5619), .I1 (g5064), .I2 (g5527));
AN2X1 gate4736(.O (g5167), .I1 (g5011), .I2 (g1556));
OR2X1 gate4737(.O (g3880), .I1 (g3658), .I2 (g3665));
OR2X1 gate4738(.O (g4440), .I1 (g4371), .I2 (g4038));
OR2X1 gate4739(.O (g3978), .I1 (g3655), .I2 (g3117));
OR2X1 gate4740(.O (g6788), .I1 (g3760), .I2 (g6767));
OR2X1 gate4741(.O (g3935), .I1 (g3464), .I2 (g2868));
OR2X1 gate4742(.O (g3982), .I1 (g3663), .I2 (g3127));
OR4X1 gate4743(.O (I8376), .I1 (g6315), .I2 (g6126), .I3 (g6129), .I4 (g6146));
OR2X1 gate4744(.O (g5625), .I1 (g5495), .I2 (g3281));
OR2X1 gate4745(.O (g6298), .I1 (g6255), .I2 (g6093));
OR3X1 gate4746(.O (g6485), .I1 (I8393), .I2 (I8394), .I3 (key_out_119));
OR2X1 gate4747(.O (g4655), .I1 (g4368), .I2 (g3660));
OR2X1 gate4748(.O (g6252), .I1 (g5905), .I2 (g2381));
OR2X1 gate4749(.O (g6176), .I1 (key_out_66), .I2 (key_out_16));
OR4X1 gate4750(.O (I8377), .I1 (g6150), .I2 (g6324), .I3 (g5180), .I4 (g5181));
OR2X1 gate4751(.O (g6286), .I1 (g6238), .I2 (g6079));
OR2X1 gate4752(.O (g3851), .I1 (g3681), .I2 (g3146));
OR2X1 gate4753(.O (g3964), .I1 (g3634), .I2 (g3089));
OR2X1 gate4754(.O (g5659), .I1 (g5551), .I2 (g5398));
OR2X1 gate4755(.O (g2928), .I1 (g2100), .I2 (g1582));
OR2X1 gate4756(.O (g6287), .I1 (g6241), .I2 (g6082));
OR2X1 gate4757(.O (g3989), .I1 (g3679), .I2 (g3144));
OR2X1 gate4758(.O (g5374), .I1 (g5215), .I2 (g4947));
OR2X1 gate4759(.O (g3971), .I1 (g3644), .I2 (g3099));
OR2X1 gate4760(.O (g6781), .I1 (g6718), .I2 (g6748));
OR2X1 gate4761(.O (g3598), .I1 (g2808), .I2 (g2821));
OR2X1 gate4762(.O (g4641), .I1 (g4347), .I2 (g3627));
OR2X1 gate4763(.O (g4450), .I1 (g4389), .I2 (g4047));
OR2X1 gate4764(.O (g3740), .I1 (g3335), .I2 (g2747));
OR4X1 gate4765(.O (I8136), .I1 (g6015), .I2 (g6212), .I3 (g4950), .I4 (g4877));
OR2X1 gate4766(.O (g5628), .I1 (g5498), .I2 (g3292));
OR2X1 gate4767(.O (g5630), .I1 (g5501), .I2 (g3309));
OR2X1 gate4768(.O (g6114), .I1 (g5904), .I2 (g5604));
OR2X1 gate4769(.O (g5323), .I1 (g5098), .I2 (g4802));
OR2X1 gate4770(.O (g5666), .I1 (g5555), .I2 (g5406));
OR4X1 gate4771(.O (I8137), .I1 (g4894), .I2 (g4904), .I3 (g4993), .I4 (g4967));
OR3X1 gate4772(.O (I8395), .I1 (g5182), .I2 (g5200), .I3 (key_out_86));
OR2X1 gate4773(.O (g3879), .I1 (g3704), .I2 (g3195));
OR4X1 gate4774(.O (I9057), .I1 (g6320), .I2 (g6828), .I3 (g6830), .I4 (g6153));
OR2X1 gate4775(.O (g4092), .I1 (g3311), .I2 (g2721));
OR4X1 gate4776(.O (I8081), .I1 (g4894), .I2 (g4904), .I3 (g4993), .I4 (g4967));
OR2X1 gate4777(.O (g4864), .I1 (g4744), .I2 (g4490));
OR3X1 gate4778(.O (g6845), .I1 (I9064), .I2 (I9065), .I3 (key_out_114));
OR2X1 gate4779(.O (g5372), .I1 (g5213), .I2 (g4942));
OR2X1 gate4780(.O (g5693), .I1 (g5632), .I2 (g5481));
OR2X1 gate4781(.O (g5804), .I1 (g5371), .I2 (g5603));
OR2X1 gate4782(.O (g6142), .I1 (g5909), .I2 (g3806));
OR2X1 gate4783(.O (I8129), .I1 (g4915), .I2 (key_out_89));
OR4X1 gate4784(.O (g6481), .I1 (I8367), .I2 (I8368), .I3 (I8369), .I4 (key_out_117));
OR2X1 gate4785(.O (g4651), .I1 (g4357), .I2 (g3643));
OR2X1 gate4786(.O (g4285), .I1 (g3490), .I2 (g3887));
OR2X1 gate4787(.O (g4500), .I1 (g4243), .I2 (g2010));
OR3X1 gate4788(.O (g5202), .I1 (g4904), .I2 (g4914), .I3 (g4894));
OR2X1 gate4789(.O (g3750), .I1 (g3372), .I2 (g2794));
OR2X1 gate4790(.O (g6267), .I1 (g2953), .I2 (g5884));
OR2X1 gate4791(.O (g4231), .I1 (g3997), .I2 (g4000));
OR2X1 gate4792(.O (g6676), .I1 (g6631), .I2 (g6555));
OR2X1 gate4793(.O (g6293), .I1 (g6244), .I2 (g6085));
OR2X1 gate4794(.O (g4205), .I1 (g3843), .I2 (g541));
OR2X1 gate4795(.O (g4634), .I1 (g4341), .I2 (g3615));
OR4X1 gate4796(.O (I8349), .I1 (I8345), .I2 (I8346), .I3 (I8347), .I4 (I8348));
OR2X1 gate4797(.O (g6703), .I1 (g6692), .I2 (g4831));
OR2X1 gate4798(.O (g3884), .I1 (g3666), .I2 (g3671));
OR2X1 gate4799(.O (g4444), .I1 (g4378), .I2 (g4042));
OR2X1 gate4800(.O (g4862), .I1 (g4739), .I2 (g4489));
OR4X1 gate4801(.O (I8119), .I1 (key_out_87), .I2 (g4993), .I3 (g4967), .I4 (g4980));
OR2X1 gate4802(.O (g3988), .I1 (g3678), .I2 (g3143));
OR2X1 gate4803(.O (g5674), .I1 (g5558), .I2 (g5419));
OR2X1 gate4804(.O (g6747), .I1 (g6614), .I2 (g6731));
OR2X1 gate4805(.O (g6855), .I1 (g6851), .I2 (g2085));
OR2X1 gate4806(.O (I8211), .I1 (g4915), .I2 (key_out_89));
OR4X1 gate4807(.O (I8386), .I1 (g6152), .I2 (g6327), .I3 (g5183), .I4 (g5177));
OR2X1 gate4808(.O (g5680), .I1 (g5562), .I2 (g5429));
OR2X1 gate4809(.O (g4946), .I1 (g4830), .I2 (g4833));
OR2X1 gate4810(.O (I8370), .I1 (g5214), .I2 (key_out_84));
OR2X1 gate4811(.O (g4436), .I1 (g4359), .I2 (g4035));
OR3X1 gate4812(.O (I8387), .I1 (g5178), .I2 (g5209), .I3 (key_out_85));
OR2X1 gate4813(.O (g6274), .I1 (g5682), .I2 (g5956));
OR2X1 gate4814(.O (g6426), .I1 (g6288), .I2 (g6119));
OR2X1 gate4815(.O (g6170), .I1 (key_out_69), .I2 (key_out_19));
OR2X1 gate4816(.O (g3996), .I1 (g3691), .I2 (g3171));
OR4X1 gate4817(.O (I8345), .I1 (g6326), .I2 (g6135), .I3 (g6140), .I4 (g6157));
OR2X1 gate4818(.O (g5623), .I1 (g5503), .I2 (g5357));
OR3X1 gate4819(.O (g6483), .I1 (I8385), .I2 (I8386), .I3 (key_out_118));
OR2X1 gate4820(.O (g4653), .I1 (g4361), .I2 (g3652));
OR2X1 gate4821(.O (g3878), .I1 (g3703), .I2 (g3191));
OR2X1 gate4822(.O (g6790), .I1 (g3765), .I2 (g6773));
OR4X1 gate4823(.O (I8359), .I1 (g5232), .I2 (g5236), .I3 (g5216), .I4 (g5226));
OR2X1 gate4824(.O (g4752), .I1 (g4452), .I2 (g4155));
OR2X1 gate4825(.O (g6461), .I1 (g6353), .I2 (g6351));
OR2X1 gate4826(.O (g3981), .I1 (g3661), .I2 (g3123));
OR2X1 gate4827(.O (g5024), .I1 (g4793), .I2 (g4600));
OR2X1 gate4828(.O (g4233), .I1 (g3912), .I2 (g471));
OR2X1 gate4829(.O (g4454), .I1 (g4395), .I2 (g4051));
OR2X1 gate4830(.O (g5672), .I1 (g5557), .I2 (g5414));
OR2X1 gate4831(.O (g5077), .I1 (g1612), .I2 (g4694));
OR2X1 gate4832(.O (g5231), .I1 (g5048), .I2 (g672));
OR2X1 gate4833(.O (g6307), .I1 (g6262), .I2 (g6096));
OR2X1 gate4834(.O (g3744), .I1 (g3345), .I2 (g2759));
OR2X1 gate4835(.O (g6251), .I1 (g5668), .I2 (g5939));
OR2X1 gate4836(.O (g6447), .I1 (g6340), .I2 (g5938));
OR4X1 gate4837(.O (I8128), .I1 (key_out_87), .I2 (g4993), .I3 (g4967), .I4 (g4980));
OR2X1 gate4838(.O (g3864), .I1 (g3693), .I2 (g3176));
OR2X1 gate4839(.O (g5044), .I1 (g4797), .I2 (g4602));
OR2X1 gate4840(.O (g4745), .I1 (g4468), .I2 (g4569));
OR2X1 gate4841(.O (g6272), .I1 (g5679), .I2 (g5953));
OR2X1 gate4842(.O (g5014), .I1 (g4785), .I2 (g4583));
OR2X1 gate4843(.O (g3871), .I1 (g3701), .I2 (g3186));
OR4X1 gate4844(.O (I7970), .I1 (g6015), .I2 (g6212), .I3 (g4950), .I4 (g4877));
OR4X1 gate4845(.O (I8348), .I1 (g5229), .I2 (g5234), .I3 (g5218), .I4 (g5225));
OR2X1 gate4846(.O (g6554), .I1 (g6337), .I2 (g6466));
OR4X1 gate4847(.O (I7987), .I1 (g6194), .I2 (g5958), .I3 (g5975), .I4 (g5997));
OR2X1 gate4848(.O (g5916), .I1 (g5728), .I2 (g3781));
OR4X1 gate4849(.O (I8118), .I1 (g6015), .I2 (g6212), .I3 (g4950), .I4 (g4877));
OR4X1 gate4850(.O (I8367), .I1 (g6313), .I2 (g6124), .I3 (g6127), .I4 (g6144));
OR2X1 gate4851(.O (g6456), .I1 (g6346), .I2 (g5954));
OR4X1 gate4852(.O (I8393), .I1 (g6317), .I2 (g6130), .I3 (g6133), .I4 (g6151));
OR2X1 gate4853(.O (g4086), .I1 (g3310), .I2 (g2720));
OR2X1 gate4854(.O (g1589), .I1 (g1059), .I2 (g1045));
OR2X1 gate4855(.O (g6118), .I1 (g5911), .I2 (g5619));
OR2X1 gate4856(.O (g6167), .I1 (key_out_70), .I2 (key_out_20));
OR2X1 gate4857(.O (g3862), .I1 (g3632), .I2 (g3641));
OR2X1 gate4858(.O (g6457), .I1 (g6352), .I2 (g6347));
OR2X1 gate4859(.O (g4635), .I1 (g4342), .I2 (g3616));
OR2X1 gate4860(.O (g6549), .I1 (g6473), .I2 (g4247));
OR2X1 gate4861(.O (g6686), .I1 (key_out_51), .I2 (g6645));
OR2X1 gate4862(.O (g5532), .I1 (g5350), .I2 (g3278));
OR4X1 gate4863(.O (g6670), .I1 (g6557), .I2 (g6634), .I3 (g4410), .I4 (g2948));
OR2X1 gate4864(.O (g5012), .I1 (g4782), .I2 (g4580));
OR2X1 gate4865(.O (g4059), .I1 (g3466), .I2 (g3425));
OR2X1 gate4866(.O (g5281), .I1 (g5074), .I2 (g5124));
OR4X1 gate4867(.O (I8358), .I1 (g5192), .I2 (g5153), .I3 (g5158), .I4 (g5197));
OR2X1 gate4868(.O (g6687), .I1 (key_out_50), .I2 (g6646));
OR2X1 gate4869(.O (g3749), .I1 (g3371), .I2 (g2793));
OR2X1 gate4870(.O (g5808), .I1 (g5373), .I2 (g5616));
OR2X1 gate4871(.O (g6691), .I1 (key_out_56), .I2 (g6603));
OR2X1 gate4872(.O (g3873), .I1 (g3649), .I2 (g3657));
OR2X1 gate4873(.O (g3869), .I1 (g3642), .I2 (g3650));
OR2X1 gate4874(.O (g6659), .I1 (g6634), .I2 (g6631));
OR2X1 gate4875(.O (g4430), .I1 (g4349), .I2 (g4015));
OR2X1 gate4876(.O (g6239), .I1 (g2339), .I2 (g6073));
OR2X1 gate4877(.O (g6545), .I1 (g6468), .I2 (g4244));
OR2X1 gate4878(.O (g4638), .I1 (g4345), .I2 (g3620));
OR2X1 gate4879(.O (g6794), .I1 (g6777), .I2 (g3333));
OR2X1 gate4880(.O (g6931), .I1 (g6741), .I2 (g6929));
OR2X1 gate4881(.O (g3990), .I1 (g3684), .I2 (g3155));
OR2X1 gate4882(.O (g5385), .I1 (g3992), .I2 (g5318));
OR2X1 gate4883(.O (g3888), .I1 (g3672), .I2 (g3682));
OR2X1 gate4884(.O (g5470), .I1 (g5359), .I2 (g5142));
OR2X1 gate4885(.O (g6300), .I1 (g6253), .I2 (g6091));
OR2X1 gate4886(.O (g4455), .I1 (g4396), .I2 (g4052));
OR3X1 gate4887(.O (g6750), .I1 (g6670), .I2 (g6625), .I3 (g6736));
OR2X1 gate4888(.O (g5678), .I1 (g5560), .I2 (g5428));
OR2X1 gate4889(.O (g3745), .I1 (g3356), .I2 (g2770));
OR2X1 gate4890(.O (g6440), .I1 (g6336), .I2 (g5935));
OR2X1 gate4891(.O (g3865), .I1 (g3637), .I2 (g3648));
OR2X1 gate4892(.O (g3833), .I1 (g3602), .I2 (g3608));
OR2X1 gate4893(.O (g4021), .I1 (g3558), .I2 (g2949));
OR2X1 gate4894(.O (g3896), .I1 (g3689), .I2 (key_out_101));
OR2X1 gate4895(.O (g5535), .I1 (g5353), .I2 (g3300));
OR2X1 gate4896(.O (g5015), .I1 (g4787), .I2 (g4588));
OR2X1 gate4897(.O (g4631), .I1 (g4340), .I2 (g3611));
OR2X1 gate4898(.O (g5246), .I1 (g5077), .I2 (g2080));
OR2X1 gate4899(.O (g6792), .I1 (g6770), .I2 (g3321));
OR4X1 gate4900(.O (I7980), .I1 (key_out_87), .I2 (g4993), .I3 (g4967), .I4 (g4980));
OR4X1 gate4901(.O (I8360), .I1 (I8356), .I2 (I8357), .I3 (I8358), .I4 (I8359));
OR2X1 gate4902(.O (g4441), .I1 (g4372), .I2 (g4039));
OR2X1 gate4903(.O (g6113), .I1 (g5902), .I2 (g5601));
OR3X1 gate4904(.O (g5388), .I1 (g5318), .I2 (g1589), .I3 (key_out_10));
OR2X1 gate4905(.O (I8379), .I1 (g5212), .I2 (key_out_83));
OR2X1 gate4906(.O (g5430), .I1 (g5161), .I2 (g4873));
OR2X1 gate4907(.O (g4458), .I1 (g4401), .I2 (g4057));
OR2X1 gate4908(.O (g3748), .I1 (g3366), .I2 (g2782));
OR2X1 gate4909(.O (g6264), .I1 (g5675), .I2 (g5948));
OR2X1 gate4910(.O (g4074), .I1 (g3301), .I2 (g2699));
OR2X1 gate4911(.O (g6450), .I1 (g6341), .I2 (g5940));
OR2X1 gate4912(.O (g4080), .I1 (g3302), .I2 (g2700));
OR2X1 gate4913(.O (g5066), .I1 (g4668), .I2 (g4672));
OR2X1 gate4914(.O (g6179), .I1 (key_out_64), .I2 (key_out_14));
OR4X1 gate4915(.O (I8209), .I1 (g6015), .I2 (g6212), .I3 (g4950), .I4 (g4877));
OR2X1 gate4916(.O (g6289), .I1 (g6240), .I2 (g6081));
OR2X1 gate4917(.O (g6658), .I1 (key_out_49), .I2 (g6620));
OR2X1 gate4918(.O (g6271), .I1 (g2955), .I2 (g5885));
OR2X1 gate4919(.O (g5662), .I1 (g5553), .I2 (g5402));
OR2X1 gate4920(.O (g5018), .I1 (g4791), .I2 (g4597));
OR2X1 gate4921(.O (I7972), .I1 (g4915), .I2 (key_out_89));
OR3X1 gate4922(.O (g5467), .I1 (g3868), .I2 (g5318), .I3 (g3992));
OR2X1 gate4923(.O (g5816), .I1 (g5378), .I2 (g5620));
OR2X1 gate4924(.O (g5700), .I1 (g5663), .I2 (g5488));
OR2X1 gate4925(.O (g4451), .I1 (g4390), .I2 (g4048));
OR2X1 gate4926(.O (g6864), .I1 (g6852), .I2 (g2089));
OR2X1 gate4927(.O (g5817), .I1 (g5380), .I2 (g5621));
OR2X1 gate4928(.O (g3883), .I1 (g3709), .I2 (g3203));
OR2X1 gate4929(.O (g5605), .I1 (g3575), .I2 (g5500));
OR3X1 gate4930(.O (I9059), .I1 (g5185), .I2 (g5198), .I3 (key_out_82));
OR2X1 gate4931(.O (g4443), .I1 (g4377), .I2 (g4041));
OR2X1 gate4932(.O (g4434), .I1 (g4355), .I2 (g4033));
OR2X1 gate4933(.O (g5669), .I1 (g5556), .I2 (g5410));
OR2X1 gate4934(.O (g5368), .I1 (g5201), .I2 (g4932));
OR4X1 gate4935(.O (I7979), .I1 (g6015), .I2 (g6212), .I3 (g4950), .I4 (g4877));
OR2X1 gate4936(.O (g5531), .I1 (g5349), .I2 (g3275));
OR2X1 gate4937(.O (g5458), .I1 (g3466), .I2 (g5311));
OR2X1 gate4938(.O (g6795), .I1 (g4867), .I2 (g6772));
OR2X1 gate4939(.O (g4936), .I1 (g4827), .I2 (g4828));
OR2X1 gate4940(.O (g5074), .I1 (g4792), .I2 (g4598));
OR2X1 gate4941(.O (g5474), .I1 (g5363), .I2 (g5146));
OR2X1 gate4942(.O (g6926), .I1 (g6798), .I2 (g6923));
OR3X1 gate4943(.O (g6754), .I1 (g6676), .I2 (g6625), .I3 (g6737));
OR2X1 gate4944(.O (g6273), .I1 (g5681), .I2 (g5955));
OR2X1 gate4945(.O (g6444), .I1 (g6338), .I2 (g5936));
OR4X1 gate4946(.O (I8378), .I1 (g5173), .I2 (g5166), .I3 (g5235), .I4 (g5245));
OR4X1 gate4947(.O (I8135), .I1 (g6194), .I2 (g5958), .I3 (g5975), .I4 (g5997));
OR3X1 gate4948(.O (g5326), .I1 (g5069), .I2 (g4410), .I3 (g3012));
OR3X1 gate4949(.O (I9066), .I1 (g5189), .I2 (g5269), .I3 (key_out_79));
OR2X1 gate4950(.O (g6927), .I1 (g6799), .I2 (g6924));
OR2X1 gate4951(.O (g3751), .I1 (g3375), .I2 (g2807));
OR2X1 gate4952(.O (g6660), .I1 (g6640), .I2 (g6637));
OR2X1 gate4953(.O (g6679), .I1 (g6637), .I2 (g6558));
OR4X1 gate4954(.O (I8208), .I1 (g6194), .I2 (g5958), .I3 (g5975), .I4 (g5997));
OR2X1 gate4955(.O (g6182), .I1 (key_out_63), .I2 (key_out_13));
OR3X1 gate4956(.O (g5327), .I1 (g5077), .I2 (g4416), .I3 (g3028));
OR2X1 gate4957(.O (g3743), .I1 (g3344), .I2 (g2758));
OR2X1 gate4958(.O (g3856), .I1 (g3686), .I2 (g3157));
OR2X1 gate4959(.O (g5303), .I1 (g5053), .I2 (g4768));
OR2X1 gate4960(.O (g5696), .I1 (g5637), .I2 (g5484));
OR2X1 gate4961(.O (g3992), .I1 (key_out_113), .I2 (key_out_9));
OR2X1 gate4962(.O (g5472), .I1 (g5361), .I2 (g5144));
OR2X1 gate4963(.O (g3863), .I1 (g3692), .I2 (g3172));
OR2X1 gate4964(.O (g6437), .I1 (g6302), .I2 (g6121));
OR2X1 gate4965(.O (g6917), .I1 (g6909), .I2 (g6910));
OR2X1 gate4966(.O (g3857), .I1 (g3687), .I2 (g3161));
OR2X1 gate4967(.O (g5533), .I1 (g5351), .I2 (g3290));
OR2X1 gate4968(.O (g5697), .I1 (g5646), .I2 (g5485));
OR2X1 gate4969(.O (g5013), .I1 (g4826), .I2 (g4621));
OR2X1 gate4970(.O (g4627), .I1 (g4333), .I2 (g3603));
OR2X1 gate4971(.O (g6454), .I1 (g6344), .I2 (g5949));
OR2X1 gate4972(.O (g6296), .I1 (g6247), .I2 (g6088));
OR2X1 gate4973(.O (g4646), .I1 (g4353), .I2 (g3635));
OR4X1 gate4974(.O (I8138), .I1 (g4980), .I2 (g4915), .I3 (key_out_89), .I4 (g5054));
OR2X1 gate4975(.O (g6189), .I1 (key_out_71), .I2 (key_out_21));
OR2X1 gate4976(.O (g3977), .I1 (g3653), .I2 (g3113));
OR4X1 gate4977(.O (I9058), .I1 (g6156), .I2 (g6331), .I3 (g5190), .I4 (g5164));
OR2X1 gate4978(.O (g6787), .I1 (g3758), .I2 (g6766));
OR2X1 gate4979(.O (g5060), .I1 (key_out_10), .I2 (g4819));
OR2X1 gate4980(.O (g6297), .I1 (g6248), .I2 (g6089));
OR2X1 gate4981(.O (g3999), .I1 (g3699), .I2 (g3181));
OR2X1 gate4982(.O (g6684), .I1 (key_out_57), .I2 (g6643));
OR4X1 gate4983(.O (I7978), .I1 (g6194), .I2 (g5958), .I3 (g5975), .I4 (g5997));
OR2X1 gate4984(.O (g6109), .I1 (g5900), .I2 (g5599));
OR2X1 gate4985(.O (g6791), .I1 (g6768), .I2 (g3307));
OR2X1 gate4986(.O (g6309), .I1 (g6265), .I2 (g6098));
OR2X1 gate4987(.O (g3732), .I1 (g3324), .I2 (g2732));
OR2X1 gate4988(.O (g3533), .I1 (g3154), .I2 (g3166));
OR4X1 gate4989(.O (I8385), .I1 (g6316), .I2 (g6128), .I3 (g6131), .I4 (g6149));
OR2X1 gate4990(.O (g6268), .I1 (g5677), .I2 (g5951));
OR2X1 gate4991(.O (g3820), .I1 (g3287), .I2 (g2671));
OR2X1 gate4992(.O (g6452), .I1 (g6342), .I2 (g5942));
OR2X1 gate4993(.O (g5626), .I1 (g5496), .I2 (g3285));
OR2X1 gate4994(.O (g4656), .I1 (g4369), .I2 (g3662));
OR2X1 gate4995(.O (g6185), .I1 (key_out_67), .I2 (key_out_17));
OR2X1 gate4996(.O (g3739), .I1 (g3334), .I2 (g2746));
OR4X1 gate4997(.O (I7989), .I1 (key_out_87), .I2 (g4993), .I3 (g4967), .I4 (g4980));
OR2X1 gate4998(.O (g3995), .I1 (g3690), .I2 (g3170));
OR4X1 gate4999(.O (I8369), .I1 (g5165), .I2 (g5159), .I3 (g5233), .I4 (g5240));
OR4X1 gate5000(.O (I7971), .I1 (key_out_87), .I2 (g4993), .I3 (g4967), .I4 (g4980));
OR2X1 gate5001(.O (g5627), .I1 (g5497), .I2 (g3286));
OR3X1 gate5002(.O (g6682), .I1 (g6478), .I2 (g6624), .I3 (g6623));
OR2X1 gate5003(.O (g3942), .I1 (g3215), .I2 (g3575));
OR2X1 gate5004(.O (g5583), .I1 (g5569), .I2 (g4020));
OR2X1 gate5005(.O (g6173), .I1 (key_out_65), .I2 (key_out_15));
OR2X1 gate5006(.O (g3954), .I1 (g3484), .I2 (g3489));
OR2X1 gate5007(.O (g6920), .I1 (g6915), .I2 (g6916));
OR2X1 gate5008(.O (g6261), .I1 (g5673), .I2 (g5944));
OR2X1 gate5009(.O (g6793), .I1 (g6771), .I2 (g3323));
OR2X1 gate5010(.O (g4948), .I1 (g4834), .I2 (g4836));
OR2X1 gate5011(.O (g6246), .I1 (g5665), .I2 (g5937));
OR2X1 gate5012(.O (g5224), .I1 (g5123), .I2 (g3630));
OR2X1 gate5013(.O (g5277), .I1 (g5023), .I2 (g4763));
OR2X1 gate5014(.O (g4438), .I1 (g4363), .I2 (g4037));
OR2X1 gate5015(.O (g4773), .I1 (g4495), .I2 (g4220));
OR2X1 gate5016(.O (g6689), .I1 (key_out_55), .I2 (g6648));
OR2X1 gate5017(.O (g3998), .I1 (g3698), .I2 (g3180));
OR4X1 gate5018(.O (I8774), .I1 (g6655), .I2 (g6653), .I3 (g6651), .I4 (g6649));
OR2X1 gate5019(.O (g3850), .I1 (g3680), .I2 (g3145));
OR2X1 gate5020(.O (g6108), .I1 (g5898), .I2 (g5598));
OR3X1 gate5021(.O (g6758), .I1 (g6673), .I2 (g6628), .I3 (g6738));
OR2X1 gate5022(.O (g2896), .I1 (g2323), .I2 (g1763));
OR2X1 gate5023(.O (g6455), .I1 (g6345), .I2 (g5952));
OR2X1 gate5024(.O (g3986), .I1 (g3667), .I2 (g3133));
OR2X1 gate5025(.O (g6846), .I1 (g5860), .I2 (g6834));
OR2X1 gate5026(.O (g3503), .I1 (g3122), .I2 (g3132));
OR4X1 gate5027(.O (I7969), .I1 (g6194), .I2 (g5958), .I3 (g5975), .I4 (g5997));
OR2X1 gate5028(.O (g4941), .I1 (g4829), .I2 (g4832));
OR2X1 gate5029(.O (g6290), .I1 (g6245), .I2 (g6086));
OR2X1 gate5030(.O (g3987), .I1 (g3669), .I2 (g3134));
OR2X1 gate5031(.O (g6847), .I1 (g5861), .I2 (g6837));
OR2X1 gate5032(.O (g6685), .I1 (key_out_53), .I2 (g6644));
OR2X1 gate5033(.O (g5295), .I1 (g5047), .I2 (g4766));
OR2X1 gate5034(.O (g4473), .I1 (g3575), .I2 (g4253));
OR2X1 gate5035(.O (g3991), .I1 (g3685), .I2 (g3156));
OR4X1 gate5036(.O (I7988), .I1 (g6015), .I2 (g6212), .I3 (g4950), .I4 (g4877));
OR2X1 gate5037(.O (g5471), .I1 (g5360), .I2 (g5143));
OR4X1 gate5038(.O (I8368), .I1 (g6148), .I2 (g6321), .I3 (g5176), .I4 (g5184));
OR2X1 gate5039(.O (g6257), .I1 (g5671), .I2 (g5941));
OR2X1 gate5040(.O (g6301), .I1 (g6254), .I2 (g6092));
OR4X1 gate5041(.O (g6673), .I1 (g6559), .I2 (g6640), .I3 (g4416), .I4 (g2950));
OR4X1 gate5042(.O (I8080), .I1 (g6015), .I2 (g6212), .I3 (g4950), .I4 (g4877));
OR2X1 gate5043(.O (g6669), .I1 (g6613), .I2 (g4679));
OR2X1 gate5044(.O (g3877), .I1 (g3651), .I2 (g3659));
OR4X1 gate5045(.O (I8126), .I1 (g6194), .I2 (g5958), .I3 (g5975), .I4 (g5997));
OR2X1 gate5046(.O (g5062), .I1 (g4661), .I2 (g4666));
OR2X1 gate5047(.O (g6480), .I1 (key_out_94), .I2 (key_out_81));
OR4X1 gate5048(.O (I8779), .I1 (g6605), .I2 (g6656), .I3 (g6654), .I4 (g6652));
OR2X1 gate5049(.O (g6688), .I1 (key_out_52), .I2 (g6647));
OR2X1 gate5050(.O (g5085), .I1 (g4694), .I2 (g4280));
OR2X1 gate5051(.O (I7981), .I1 (g4915), .I2 (key_out_89));
OR4X1 gate5052(.O (I8127), .I1 (g6015), .I2 (g6212), .I3 (g4950), .I4 (g4877));
OR2X1 gate5053(.O (g4433), .I1 (g4354), .I2 (g4032));
OR4X1 gate5054(.O (I8346), .I1 (g6159), .I2 (g6334), .I3 (g5163), .I4 (g5191));
OR2X1 gate5055(.O (g5812), .I1 (g5376), .I2 (g5618));
OR2X1 gate5056(.O (g4859), .I1 (g4730), .I2 (g4486));
OR2X1 gate5057(.O (g6665), .I1 (I8778), .I2 (I8779));
OR2X1 gate5058(.O (g5473), .I1 (g5362), .I2 (g5145));
OR4X1 gate5059(.O (I8347), .I1 (g5188), .I2 (g5157), .I3 (g5154), .I4 (g5193));
OR2X1 gate5060(.O (g6303), .I1 (g6258), .I2 (g6094));
OR2X1 gate5061(.O (g5069), .I1 (g1595), .I2 (g4688));
OR4X1 gate5062(.O (I9064), .I1 (g6323), .I2 (g6829), .I3 (g6831), .I4 (g6155));
OR2X1 gate5063(.O (g4497), .I1 (g4166), .I2 (g3784));
OR4X1 gate5064(.O (I8210), .I1 (key_out_87), .I2 (g4993), .I3 (g4967), .I4 (g4980));
OR2X1 gate5065(.O (g5377), .I1 (g5217), .I2 (g4949));
OR2X1 gate5066(.O (g3837), .I1 (g3609), .I2 (g3613));
OR2X1 gate5067(.O (g6116), .I1 (g5910), .I2 (g5617));
OR4X1 gate5068(.O (I8117), .I1 (g6194), .I2 (g5958), .I3 (g5975), .I4 (g5997));
OR2X1 gate5069(.O (g4001), .I1 (g3702), .I2 (g3190));
OR2X1 gate5070(.O (g3842), .I1 (g3670), .I2 (g3135));
OR2X1 gate5071(.O (g5291), .I1 (g5043), .I2 (g4764));
OR2X1 gate5072(.O (g3941), .I1 (g3479), .I2 (g2873));
OR2X1 gate5073(.O (g5694), .I1 (g5633), .I2 (g5482));
OR2X1 gate5074(.O (g6936), .I1 (g5438), .I2 (g6935));
OR2X1 gate5075(.O (g4068), .I1 (g3293), .I2 (g2685));
OR4X1 gate5076(.O (I8079), .I1 (g6194), .I2 (g5958), .I3 (g5975), .I4 (g5997));
OR2X1 gate5077(.O (g4468), .I1 (g4214), .I2 (g3831));
OR2X1 gate5078(.O (g4866), .I1 (g4756), .I2 (g4491));
OR2X1 gate5079(.O (g3829), .I1 (g3294), .I2 (g3305));
OR4X1 gate5080(.O (I8356), .I1 (g6311), .I2 (g6123), .I3 (g6125), .I4 (g6141));
OR2X1 gate5081(.O (g3733), .I1 (g3325), .I2 (g2733));
OR2X1 gate5082(.O (g6937), .I1 (g4616), .I2 (g6934));
OR2X1 gate5083(.O (g6479), .I1 (key_out_121), .I2 (key_out_80));
OR2X1 gate5084(.O (g6294), .I1 (g6249), .I2 (g6090));
OR2X1 gate5085(.O (g5065), .I1 (g4667), .I2 (g4671));
OR2X1 gate5086(.O (g5228), .I1 (g5096), .I2 (g4800));
OR4X1 gate5087(.O (I8357), .I1 (g6145), .I2 (g6318), .I3 (g5171), .I4 (g5187));
OR2X1 gate5088(.O (g3849), .I1 (g3618), .I2 (g3625));
OR2X1 gate5089(.O (g6704), .I1 (g6660), .I2 (g492));
OR2X1 gate5090(.O (g4599), .I1 (g3499), .I2 (g4230));
OR2X1 gate5091(.O (g6453), .I1 (g6343), .I2 (g5945));
OR2X1 gate5092(.O (g4544), .I1 (g4410), .I2 (g2995));
OR4X1 gate5093(.O (I8778), .I1 (g6612), .I2 (g6611), .I3 (g6609), .I4 (g6607));
OR2X1 gate5094(.O (g2924), .I1 (g2095), .I2 (g1573));
OR2X1 gate5095(.O (g4427), .I1 (g4373), .I2 (g3668));
OR2X1 gate5096(.O (g4446), .I1 (g4383), .I2 (g4043));
OR2X1 gate5097(.O (g3870), .I1 (g3700), .I2 (g3182));
OR3X1 gate5098(.O (g6683), .I1 (g6465), .I2 (g6622), .I3 (g6621));
OR2X1 gate5099(.O (g5676), .I1 (g5559), .I2 (g5424));
OR2X1 gate5100(.O (g4637), .I1 (g4344), .I2 (g3619));
OR2X1 gate5101(.O (g3972), .I1 (g3646), .I2 (g3103));
OR2X1 gate5102(.O (g6782), .I1 (g6719), .I2 (g6749));
OR2X1 gate5103(.O (g6661), .I1 (I8773), .I2 (I8774));
OR2X1 gate5104(.O (g4757), .I1 (g4456), .I2 (g4158));
OR2X1 gate5105(.O (g6292), .I1 (g6243), .I2 (g6084));
OR2X1 gate5106(.O (g4811), .I1 (g4429), .I2 (g4432));
OR2X1 gate5107(.O (g4642), .I1 (g4348), .I2 (g3628));
OR2X1 gate5108(.O (g4447), .I1 (g4384), .I2 (g4044));
OR2X1 gate5109(.O (g5624), .I1 (g5494), .I2 (g3280));
OR2X1 gate5110(.O (g5068), .I1 (g4673), .I2 (g4677));
OR2X1 gate5111(.O (g4654), .I1 (g4362), .I2 (g3654));
OR2X1 gate5112(.O (g3891), .I1 (g3683), .I2 (g3688));
OR2X1 gate5113(.O (g3913), .I1 (g3449), .I2 (g2860));
OR2X1 gate5114(.O (I7990), .I1 (g4915), .I2 (key_out_89));
OR2X1 gate5115(.O (g6702), .I1 (g6659), .I2 (g496));
OR2X1 gate5116(.O (g6919), .I1 (g6912), .I2 (g6914));
OR2X1 gate5117(.O (I8120), .I1 (g4915), .I2 (key_out_89));
OR2X1 gate5118(.O (g4243), .I1 (g4053), .I2 (g4058));
OR2X1 gate5119(.O (g5699), .I1 (g5660), .I2 (g5487));
OR2X1 gate5120(.O (g5241), .I1 (g5069), .I2 (g2067));
OR2X1 gate5121(.O (g4234), .I1 (g3921), .I2 (g478));
OR2X1 gate5122(.O (g3815), .I1 (g3282), .I2 (g2659));
OR2X1 gate5123(.O (g5386), .I1 (g5227), .I2 (g669));
OR2X1 gate5124(.O (g6789), .I1 (g3764), .I2 (g6769));
OR4X1 gate5125(.O (I8082), .I1 (g4980), .I2 (g4915), .I3 (key_out_89), .I4 (g5054));
OR2X1 gate5126(.O (g5370), .I1 (g5211), .I2 (g4937));
OR2X1 gate5127(.O (g3828), .I1 (g3304), .I2 (g1351));
OR4X1 gate5128(.O (I9065), .I1 (g6158), .I2 (g6333), .I3 (g5152), .I4 (g5156));
OR2X1 gate5129(.O (g3746), .I1 (g3357), .I2 (g2771));
OR2X1 gate5130(.O (g5083), .I1 (g4688), .I2 (g4271));
OR2X1 gate5131(.O (g6907), .I1 (g6874), .I2 (g3358));
OR2X1 gate5132(.O (g5622), .I1 (g5492), .I2 (g3277));
OR2X1 gate5133(.O (g6690), .I1 (key_out_54), .I2 (g6650));
OR4X1 gate5134(.O (g6482), .I1 (I8376), .I2 (I8377), .I3 (I8378), .I4 (key_out_116));
OR2X1 gate5135(.O (g4652), .I1 (g4358), .I2 (g3645));
OR2X1 gate5136(.O (g4549), .I1 (g4416), .I2 (g3013));
OR2X1 gate5137(.O (g3747), .I1 (g3365), .I2 (g2781));
OR2X1 gate5138(.O (g3855), .I1 (g3626), .I2 (g3631));
OR2X1 gate5139(.O (g5695), .I1 (g5635), .I2 (g5483));
OR2X1 gate5140(.O (g6110), .I1 (key_out_68), .I2 (key_out_18));
OR2X1 gate5141(.O (g6310), .I1 (g6269), .I2 (g6099));
OR2X1 gate5142(.O (g5016), .I1 (g4789), .I2 (g4592));
OR3X1 gate5143(.O (g6762), .I1 (g6679), .I2 (g6628), .I3 (g6739));
OR2X1 gate5144(.O (g4740), .I1 (g4448), .I2 (g4154));
OR4X1 gate5145(.O (I8394), .I1 (g6154), .I2 (g6329), .I3 (g5186), .I4 (g5172));
OR2X1 gate5146(.O (g6556), .I1 (g6339), .I2 (g6467));
OR2X1 gate5147(.O (g6930), .I1 (g6740), .I2 (g6928));
OR2X1 gate5148(.O (g3599), .I1 (g2935), .I2 (g1637));
OR2X1 gate5149(.O (g3821), .I1 (g2951), .I2 (g3466));
OR2X1 gate5150(.O (g4860), .I1 (g4735), .I2 (g4488));
OR2X1 gate5151(.O (g6237), .I1 (g5912), .I2 (g2381));
OR2X1 gate5152(.O (g4645), .I1 (g4352), .I2 (g3633));
OR3X1 gate5153(.O (g6844), .I1 (I9057), .I2 (I9058), .I3 (key_out_115));
OR4X1 gate5154(.O (I8773), .I1 (g6610), .I2 (g6608), .I3 (g6606), .I4 (g6604));
OR2X1 gate5155(.O (g5629), .I1 (g5499), .I2 (g3298));
OR2X1 gate5156(.O (g4607), .I1 (g4232), .I2 (g3899));
OR2X1 gate5157(.O (g6705), .I1 (g6693), .I2 (g4835));
OR2X1 gate5158(.O (g5800), .I1 (g5369), .I2 (g5600));
OR2X1 gate5159(.O (g6242), .I1 (g2356), .I2 (g6075));
OR2X1 gate5160(.O (g3841), .I1 (g3614), .I2 (g3617));
OR2X1 gate5161(.O (g6918), .I1 (g6911), .I2 (g6913));
OR2X1 gate5162(.O (g5348), .I1 (g5317), .I2 (g5122));
OR2X1 gate5163(.O (g3858), .I1 (g3629), .I2 (g3636));
OR2X1 gate5164(.O (g5698), .I1 (g5648), .I2 (g5486));
OR2X1 gate5165(.O (g4630), .I1 (g4339), .I2 (g3610));
OR2X1 gate5166(.O (g6921), .I1 (g6908), .I2 (g6816));
OR2X1 gate5167(.O (g5367), .I1 (g5199), .I2 (g4928));
ND3X1 gate5168(.O (g1777), .I1 (g1060), .I2 (g102), .I3 (g89));
ND2X1 gate5169(.O (I7217), .I1 (g152), .I2 (I7216));
ND2X1 gate5170(.O (I7571), .I1 (g5678), .I2 (I7569));
ND4X1 gate5171(.O (g5686), .I1 (g5546), .I2 (g1017), .I3 (g1551), .I4 (g2916));
ND2X1 gate5172(.O (I2073), .I1 (g15), .I2 (key_out_25));
ND2X1 gate5173(.O (I2796), .I1 (g804), .I2 (I2795));
ND2X1 gate5174(.O (g948), .I1 (I2014), .I2 (I2015));
ND2X1 gate5175(.O (I4205), .I1 (g743), .I2 (I4203));
ND2X1 gate5176(.O (I3875), .I1 (g285), .I2 (I3874));
ND3X1 gate5177(.O (g3330), .I1 (g1815), .I2 (g1797), .I3 (g3109));
ND2X1 gate5178(.O (g4151), .I1 (I5536), .I2 (I5537));
ND3X1 gate5179(.O (g2435), .I1 (g1138), .I2 (g1777), .I3 (g1157));
ND2X1 gate5180(.O (I5658), .I1 (key_out_105), .I2 (I5657));
ND2X1 gate5181(.O (g1558), .I1 (I2527), .I2 (I2528));
ND2X1 gate5182(.O (I4444), .I1 (g2092), .I2 (g606));
ND2X1 gate5183(.O (I5271), .I1 (g3710), .I2 (key_out_22));
ND2X1 gate5184(.O (I2898), .I1 (g1027), .I2 (I2897));
ND2X1 gate5185(.O (I2797), .I1 (g798), .I2 (I2795));
ND2X1 gate5186(.O (I2245), .I1 (key_out_32), .I2 (I2244));
ND2X1 gate5187(.O (I3988), .I1 (g291), .I2 (g2544));
ND2X1 gate5188(.O (g1574), .I1 (I2543), .I2 (I2544));
ND4X1 gate5189(.O (g3529), .I1 (g3200), .I2 (g2215), .I3 (g2976), .I4 (g2968));
ND2X1 gate5190(.O (I1963), .I1 (g242), .I2 (I1961));
ND2X1 gate5191(.O (I5209), .I1 (key_out_5), .I2 (key_out_37));
ND2X1 gate5192(.O (I7562), .I1 (g74), .I2 (g5676));
ND2X1 gate5193(.O (g5506), .I1 (I7231), .I2 (I7232));
ND2X1 gate5194(.O (g5111), .I1 (I6744), .I2 (I6745));
ND2X1 gate5195(.O (I4182), .I1 (g2292), .I2 (g749));
ND2X1 gate5196(.O (I6186), .I1 (g4301), .I2 (key_out_36));
ND2X1 gate5197(.O (I7441), .I1 (g594), .I2 (I7439));
ND2X1 gate5198(.O (I6026), .I1 (g4223), .I2 (g4221));
ND2X1 gate5199(.O (I2768), .I1 (g743), .I2 (I2766));
ND2X1 gate5200(.O (I3933), .I1 (g288), .I2 (g2473));
ND3X1 gate5201(.O (g5853), .I1 (g5638), .I2 (g2053), .I3 (g1076));
ND2X1 gate5202(.O (g2731), .I1 (I3894), .I2 (I3895));
ND2X1 gate5203(.O (g5507), .I1 (I7238), .I2 (I7239));
ND2X1 gate5204(.O (g2966), .I1 (I4160), .I2 (I4161));
ND2X1 gate5205(.O (I2934), .I1 (g1436), .I2 (I2933));
ND2X1 gate5206(.O (I3179), .I1 (g736), .I2 (I3177));
ND2X1 gate5207(.O (I6187), .I1 (g3955), .I2 (key_out_36));
ND2X1 gate5208(.O (I6027), .I1 (g4223), .I2 (I6026));
ND3X1 gate5209(.O (g2009), .I1 (g901), .I2 (g1387), .I3 (g905));
ND2X1 gate5210(.O (I4233), .I1 (g2267), .I2 (g798));
ND2X1 gate5211(.O (g2769), .I1 (I3953), .I2 (I3954));
ND2X1 gate5212(.O (g1044), .I1 (I2081), .I2 (I2082));
ND4X1 gate5213(.O (g4674), .I1 (g4550), .I2 (g1514), .I3 (g2107), .I4 (g2897));
ND2X1 gate5214(.O (I7569), .I1 (g79), .I2 (g5678));
ND2X1 gate5215(.O (I6391), .I1 (g4504), .I2 (key_out_59));
ND4X1 gate5216(.O (g3525), .I1 (g3192), .I2 (g3002), .I3 (g2197), .I4 (g2179));
ND4X1 gate5217(.O (g4680), .I1 (g4550), .I2 (g1514), .I3 (g1006), .I4 (g2897));
ND2X1 gate5218(.O (I2081), .I1 (g25), .I2 (key_out_24));
ND2X1 gate5219(.O (I8195), .I1 (g471), .I2 (I8194));
ND2X1 gate5220(.O (g1534), .I1 (I2498), .I2 (I2499));
ND2X1 gate5221(.O (I2497), .I1 (key_out_109), .I2 (key_out_108));
ND2X1 gate5222(.O (g939), .I1 (I1987), .I2 (I1988));
ND2X1 gate5223(.O (I5269), .I1 (g3705), .I2 (g3710));
ND3X1 gate5224(.O (g3985), .I1 (g1138), .I2 (g3718), .I3 (g2142));
ND2X1 gate5225(.O (g1036), .I1 (I2061), .I2 (I2062));
ND2X1 gate5226(.O (I2676), .I1 (g131), .I2 (I2674));
ND2X1 gate5227(.O (g1749), .I1 (I2767), .I2 (I2768));
ND2X1 gate5228(.O (g6097), .I1 (g2954), .I2 (g5857));
ND3X1 gate5229(.O (g6783), .I1 (g6747), .I2 (g5068), .I3 (g5066));
ND2X1 gate5230(.O (g5776), .I1 (I7528), .I2 (I7529));
ND2X1 gate5231(.O (I7434), .I1 (g5554), .I2 (I7432));
ND2X1 gate5232(.O (g1042), .I1 (I2073), .I2 (I2074));
ND2X1 gate5233(.O (I7210), .I1 (g5367), .I2 (I7208));
ND4X1 gate5234(.O (g3530), .I1 (g3204), .I2 (g3023), .I3 (g2197), .I4 (g2179));
ND2X1 gate5235(.O (I6964), .I1 (g586), .I2 (I6962));
ND2X1 gate5236(.O (I5208), .I1 (key_out_2), .I2 (key_out_37));
ND2X1 gate5237(.O (I5302), .I1 (g3505), .I2 (I5300));
ND2X1 gate5238(.O (g5777), .I1 (I7535), .I2 (I7536));
ND2X1 gate5239(.O (g4613), .I1 (I6195), .I2 (I6196));
ND2X1 gate5240(.O (I2544), .I1 (g774), .I2 (I2542));
ND2X1 gate5241(.O (g1138), .I1 (g102), .I2 (g98));
ND2X1 gate5242(.O (I1994), .I1 (g504), .I2 (g218));
ND2X1 gate5243(.O (I4445), .I1 (g2092), .I2 (I4444));
ND2X1 gate5244(.O (I2061), .I1 (g7), .I2 (key_out_26));
ND2X1 gate5245(.O (I5189), .I1 (key_out_6), .I2 (key_out_61));
ND2X1 gate5246(.O (g4903), .I1 (g4717), .I2 (g858));
ND2X1 gate5247(.O (I3178), .I1 (g1706), .I2 (I3177));
ND2X1 gate5248(.O (I4920), .I1 (g3522), .I2 (I4919));
ND2X1 gate5249(.O (g2951), .I1 (g2142), .I2 (g1797));
ND4X1 gate5250(.O (g3518), .I1 (g3177), .I2 (g3023), .I3 (g3007), .I4 (g2981));
ND2X1 gate5251(.O (I2003), .I1 (g500), .I2 (g212));
ND3X1 gate5252(.O (g6717), .I1 (g6669), .I2 (g5065), .I3 (g5062));
ND2X1 gate5253(.O (I3916), .I1 (g2449), .I2 (I3914));
ND4X1 gate5254(.O (g5864), .I1 (g5649), .I2 (g1529), .I3 (g1088), .I4 (g2068));
ND3X1 gate5255(.O (g2008), .I1 (g866), .I2 (g873), .I3 (g1784));
ND2X1 gate5256(.O (I5309), .I1 (g3512), .I2 (I5307));
ND2X1 gate5257(.O (I7432), .I1 (g111), .I2 (g5554));
ND2X1 gate5258(.O (I4203), .I1 (g2255), .I2 (g743));
ND4X1 gate5259(.O (g3521), .I1 (g3187), .I2 (g3023), .I3 (g3007), .I4 (g2179));
ND2X1 gate5260(.O (I5759), .I1 (g3836), .I2 (g3503));
ND2X1 gate5261(.O (I6962), .I1 (g4874), .I2 (g586));
ND2X1 gate5262(.O (I6659), .I1 (g4762), .I2 (g3541));
ND2X1 gate5263(.O (I4940), .I1 (g3437), .I2 (I4939));
ND2X1 gate5264(.O (I2935), .I1 (g345), .I2 (I2933));
ND2X1 gate5265(.O (g2266), .I1 (I3412), .I2 (I3413));
ND2X1 gate5266(.O (I2542), .I1 (g821), .I2 (g774));
ND2X1 gate5267(.O (I3412), .I1 (g1419), .I2 (I3411));
ND2X1 gate5268(.O (I3189), .I1 (g1716), .I2 (I3188));
ND2X1 gate5269(.O (g5634), .I1 (g5563), .I2 (g4767));
ND2X1 gate5270(.O (I3990), .I1 (g2544), .I2 (I3988));
ND2X1 gate5271(.O (g2960), .I1 (I4151), .I2 (I4152));
ND2X1 gate5272(.O (g5926), .I1 (g5741), .I2 (g639));
ND4X1 gate5273(.O (g3511), .I1 (g3158), .I2 (g3002), .I3 (g2976), .I4 (g2968));
ND2X1 gate5274(.O (I7439), .I1 (g5515), .I2 (g594));
ND2X1 gate5275(.O (I2090), .I1 (g33), .I2 (key_out_23));
ND4X1 gate5276(.O (g5862), .I1 (g5649), .I2 (g1529), .I3 (g1535), .I4 (g2068));
ND2X1 gate5277(.O (I9050), .I1 (g6832), .I2 (g3598));
ND2X1 gate5278(.O (I5766), .I1 (g3961), .I2 (g3957));
ND3X1 gate5279(.O (g1582), .I1 (g784), .I2 (g774), .I3 (g821));
ND2X1 gate5280(.O (g1793), .I1 (g94), .I2 (g1084));
ND2X1 gate5281(.O (g3968), .I1 (I5227), .I2 (I5228));
ND2X1 gate5282(.O (I7527), .I1 (g49), .I2 (g5662));
ND2X1 gate5283(.O (I5226), .I1 (g3259), .I2 (g3263));
ND2X1 gate5284(.O (g4049), .I1 (g3677), .I2 (g3425));
ND2X1 gate5285(.O (I7224), .I1 (g161), .I2 (I7223));
ND2X1 gate5286(.O (I5767), .I1 (g3961), .I2 (key_out_34));
ND2X1 gate5287(.O (I5535), .I1 (g3907), .I2 (g654));
ND2X1 gate5288(.O (I5227), .I1 (g3259), .I2 (key_out_29));
ND2X1 gate5289(.O (g5947), .I1 (g5821), .I2 (g2944));
ND2X1 gate5290(.O (g3742), .I1 (I4920), .I2 (I4921));
ND4X1 gate5291(.O (g5873), .I1 (g5649), .I2 (g1017), .I3 (g1564), .I4 (g2113));
ND2X1 gate5292(.O (g4504), .I1 (I6027), .I2 (I6028));
ND2X1 gate5293(.O (I7244), .I1 (g188), .I2 (g5377));
ND3X1 gate5294(.O (g5869), .I1 (g5649), .I2 (g1076), .I3 (g2081));
ND2X1 gate5295(.O (I5188), .I1 (key_out_8), .I2 (key_out_61));
ND2X1 gate5296(.O (g3983), .I1 (I5270), .I2 (I5271));
ND4X1 gate5297(.O (g4678), .I1 (g2897), .I2 (g2101), .I3 (g1514), .I4 (g4550));
ND2X1 gate5298(.O (g6843), .I1 (I9051), .I2 (I9052));
ND2X1 gate5299(.O (g3961), .I1 (key_out_78), .I2 (key_out_72));
ND2X1 gate5300(.O (I5308), .I1 (g478), .I2 (I5307));
ND2X1 gate5301(.O (I2506), .I1 (key_out_107), .I2 (key_out_106));
ND2X1 gate5302(.O (I3445), .I1 (g1689), .I2 (g729));
ND2X1 gate5303(.O (g2061), .I1 (I3169), .I2 (I3170));
ND2X1 gate5304(.O (I3169), .I1 (g1540), .I2 (I3168));
ND3X1 gate5305(.O (g6740), .I1 (g6703), .I2 (g6457), .I3 (g4936));
ND2X1 gate5306(.O (I7556), .I1 (g69), .I2 (I7555));
ND2X1 gate5307(.O (g4007), .I1 (I5308), .I2 (I5309));
ND2X1 gate5308(.O (I5196), .I1 (key_out_7), .I2 (key_out_35));
ND2X1 gate5309(.O (I7563), .I1 (g74), .I2 (I7562));
ND2X1 gate5310(.O (g5684), .I1 (I7440), .I2 (I7441));
ND2X1 gate5311(.O (I2507), .I1 (key_out_107), .I2 (I2506));
ND2X1 gate5312(.O (I1995), .I1 (g504), .I2 (I1994));
ND2X1 gate5313(.O (g2307), .I1 (I3446), .I2 (I3447));
ND2X1 gate5314(.O (I7237), .I1 (g179), .I2 (g5374));
ND2X1 gate5315(.O (g2858), .I1 (g1815), .I2 (g2577));
ND2X1 gate5316(.O (g2757), .I1 (I3934), .I2 (I3935));
ND2X1 gate5317(.O (I6744), .I1 (g4708), .I2 (I6743));
ND2X1 gate5318(.O (I4183), .I1 (g2292), .I2 (I4182));
ND2X1 gate5319(.O (I7557), .I1 (g5674), .I2 (I7555));
ND2X1 gate5320(.O (I2300), .I1 (g830), .I2 (I2299));
ND2X1 gate5321(.O (I3188), .I1 (g1716), .I2 (g791));
ND4X1 gate5322(.O (g5865), .I1 (g5649), .I2 (g1088), .I3 (g1076), .I4 (g2068));
ND2X1 gate5323(.O (I5197), .I1 (key_out_4), .I2 (key_out_35));
ND2X1 gate5324(.O (I4161), .I1 (g619), .I2 (I4159));
ND2X1 gate5325(.O (I3741), .I1 (g349), .I2 (I3739));
ND2X1 gate5326(.O (g5019), .I1 (I6660), .I2 (key_out_62));
ND2X1 gate5327(.O (I5257), .I1 (g3714), .I2 (g3719));
ND4X1 gate5328(.O (g3532), .I1 (g3212), .I2 (g2215), .I3 (g3007), .I4 (g2981));
ND2X1 gate5329(.O (I2528), .I1 (g719), .I2 (I2526));
ND2X1 gate5330(.O (I5301), .I1 (g471), .I2 (I5300));
ND2X1 gate5331(.O (g1743), .I1 (g1064), .I2 (g94));
ND2X1 gate5332(.O (g1411), .I1 (g314), .I2 (g873));
ND2X1 gate5333(.O (g3012), .I1 (I4204), .I2 (I4205));
ND2X1 gate5334(.O (g5504), .I1 (I7217), .I2 (I7218));
ND2X1 gate5335(.O (I6175), .I1 (g4236), .I2 (g571));
ND2X1 gate5336(.O (I3455), .I1 (g1691), .I2 (g784));
ND2X1 gate5337(.O (I6500), .I1 (g4504), .I2 (key_out_91));
ND3X1 gate5338(.O (g1573), .I1 (g729), .I2 (g719), .I3 (g766));
ND2X1 gate5339(.O (I3846), .I1 (g284), .I2 (g2370));
ND2X1 gate5340(.O (I4210), .I1 (g2294), .I2 (g804));
ND2X1 gate5341(.O (g4803), .I1 (I6474), .I2 (I6475));
ND2X1 gate5342(.O (g3109), .I1 (g2360), .I2 (g1064));
ND2X1 gate5343(.O (g2698), .I1 (I3847), .I2 (I3848));
ND2X1 gate5344(.O (g3957), .I1 (key_out_76), .I2 (key_out_74));
ND2X1 gate5345(.O (I6499), .I1 (g4504), .I2 (g3541));
ND4X1 gate5346(.O (g4816), .I1 (g996), .I2 (g4550), .I3 (g1518), .I4 (g2073));
ND2X1 gate5347(.O (I3847), .I1 (g284), .I2 (I3846));
ND2X1 gate5348(.O (I7520), .I1 (g361), .I2 (g5659));
ND2X1 gate5349(.O (I4784), .I1 (g622), .I2 (I4782));
ND2X1 gate5350(.O (I1952), .I1 (g524), .I2 (I1951));
ND4X1 gate5351(.O (g3539), .I1 (g2591), .I2 (g2215), .I3 (g2197), .I4 (g2981));
ND2X1 gate5352(.O (I8202), .I1 (g478), .I2 (I8201));
ND2X1 gate5353(.O (I1986), .I1 (g508), .I2 (g224));
ND2X1 gate5354(.O (I2933), .I1 (g1436), .I2 (g345));
ND2X1 gate5355(.O (I5760), .I1 (g3836), .I2 (I5759));
ND2X1 gate5356(.O (g4301), .I1 (key_out_77), .I2 (key_out_88));
ND2X1 gate5357(.O (I1970), .I1 (g516), .I2 (I1969));
ND2X1 gate5358(.O (I7225), .I1 (g5370), .I2 (I7223));
ND2X1 gate5359(.O (I6660), .I1 (g4762), .I2 (key_out_33));
ND2X1 gate5360(.O (g5502), .I1 (I7209), .I2 (I7210));
ND2X1 gate5361(.O (I3168), .I1 (g1540), .I2 (g1534));
ND2X1 gate5362(.O (I1987), .I1 (g508), .I2 (I1986));
ND2X1 gate5363(.O (g1316), .I1 (I2300), .I2 (I2301));
ND2X1 gate5364(.O (I2674), .I1 (g710), .I2 (g131));
ND4X1 gate5365(.O (g4669), .I1 (g4550), .I2 (g1017), .I3 (g1680), .I4 (g2897));
ND2X1 gate5366(.O (I3411), .I1 (g1419), .I2 (g616));
ND2X1 gate5367(.O (I7245), .I1 (g188), .I2 (I7244));
ND2X1 gate5368(.O (g2607), .I1 (I3740), .I2 (I3741));
ND2X1 gate5369(.O (g5308), .I1 (I6963), .I2 (I6964));
ND2X1 gate5370(.O (g2311), .I1 (I3456), .I2 (I3457));
ND4X1 gate5371(.O (g3535), .I1 (g3216), .I2 (g2215), .I3 (g2197), .I4 (g2968));
ND2X1 gate5372(.O (g5455), .I1 (g2330), .I2 (g5311));
ND2X1 gate5373(.O (I4782), .I1 (g2846), .I2 (g622));
ND2X1 gate5374(.O (I9052), .I1 (g3598), .I2 (I9050));
ND2X1 gate5375(.O (I3126), .I1 (g1279), .I2 (I3125));
ND2X1 gate5376(.O (I3400), .I1 (g135), .I2 (I3398));
ND2X1 gate5377(.O (I4526), .I1 (g2909), .I2 (g646));
ND2X1 gate5378(.O (g5780), .I1 (I7556), .I2 (I7557));
ND2X1 gate5379(.O (g3246), .I1 (I4527), .I2 (I4528));
ND3X1 gate5380(.O (g3502), .I1 (g1411), .I2 (g1402), .I3 (g2795));
ND2X1 gate5381(.O (g4608), .I1 (I6176), .I2 (I6177));
ND2X1 gate5382(.O (I4919), .I1 (g3522), .I2 (g650));
ND3X1 gate5383(.O (g2100), .I1 (g1588), .I2 (g804), .I3 (g791));
ND2X1 gate5384(.O (I7230), .I1 (g170), .I2 (g5372));
ND2X1 gate5385(.O (I7433), .I1 (g111), .I2 (I7432));
ND2X1 gate5386(.O (I3127), .I1 (g1276), .I2 (I3125));
ND2X1 gate5387(.O (g3028), .I1 (I4234), .I2 (I4235));
ND2X1 gate5388(.O (I2795), .I1 (g804), .I2 (g798));
ND2X1 gate5389(.O (I5784), .I1 (g628), .I2 (I5782));
ND2X1 gate5390(.O (I4527), .I1 (g2909), .I2 (I4526));
ND2X1 gate5391(.O (I7550), .I1 (g5672), .I2 (I7548));
ND2X1 gate5392(.O (I4546), .I1 (g2853), .I2 (I4545));
ND2X1 gate5393(.O (I6745), .I1 (g582), .I2 (I6743));
ND2X1 gate5394(.O (I5294), .I1 (g625), .I2 (I5292));
ND2X1 gate5395(.O (I6963), .I1 (g4874), .I2 (I6962));
ND3X1 gate5396(.O (g3741), .I1 (g901), .I2 (g3433), .I3 (g2340));
ND2X1 gate5397(.O (g1157), .I1 (g89), .I2 (g107));
ND2X1 gate5398(.O (I2499), .I1 (key_out_108), .I2 (I2497));
ND2X1 gate5399(.O (g937), .I1 (I1979), .I2 (I1980));
ND2X1 gate5400(.O (g4472), .I1 (g3380), .I2 (g4253));
ND3X1 gate5401(.O (g2010), .I1 (g1473), .I2 (g1470), .I3 (g1459));
ND2X1 gate5402(.O (g928), .I1 (I1962), .I2 (I1963));
ND2X1 gate5403(.O (I7097), .I1 (g5194), .I2 (g574));
ND2X1 gate5404(.O (I4547), .I1 (g353), .I2 (I4545));
ND2X1 gate5405(.O (I3697), .I1 (g1570), .I2 (g642));
ND2X1 gate5406(.O (I3914), .I1 (g287), .I2 (g2449));
ND2X1 gate5407(.O (I2543), .I1 (g821), .I2 (I2542));
ND2X1 gate5408(.O (I3413), .I1 (g616), .I2 (I3411));
ND2X1 gate5409(.O (I7218), .I1 (g5368), .I2 (I7216));
ND2X1 gate5410(.O (I7312), .I1 (g5364), .I2 (I7311));
ND4X1 gate5411(.O (g3538), .I1 (g2588), .I2 (g2215), .I3 (g2197), .I4 (g2179));
ND2X1 gate5412(.O (g5505), .I1 (I7224), .I2 (I7225));
ND2X1 gate5413(.O (g1075), .I1 (I2109), .I2 (I2110));
ND2X1 gate5414(.O (I2014), .I1 (g532), .I2 (I2013));
ND2X1 gate5415(.O (g2804), .I1 (I4009), .I2 (I4010));
ND3X1 gate5416(.O (g6742), .I1 (g6683), .I2 (g932), .I3 (g6716));
ND2X1 gate5417(.O (I6185), .I1 (g4301), .I2 (g3955));
ND4X1 gate5418(.O (g5863), .I1 (g5649), .I2 (g1076), .I3 (g1535), .I4 (g2068));
ND2X1 gate5419(.O (I3739), .I1 (g2021), .I2 (g349));
ND2X1 gate5420(.O (I2022), .I1 (g528), .I2 (I2021));
ND2X1 gate5421(.O (I5782), .I1 (g3810), .I2 (g628));
ND2X1 gate5422(.O (I7576), .I1 (g84), .I2 (g5680));
ND4X1 gate5423(.O (g5688), .I1 (g5546), .I2 (g1585), .I3 (g2084), .I4 (g2916));
ND4X1 gate5424(.O (g5857), .I1 (g5638), .I2 (g1552), .I3 (g1017), .I4 (g2062));
ND2X1 gate5425(.O (I3190), .I1 (g791), .I2 (I3188));
ND2X1 gate5426(.O (I5292), .I1 (g3421), .I2 (g625));
ND2X1 gate5427(.O (g1764), .I1 (I2796), .I2 (I2797));
ND2X1 gate5428(.O (I3954), .I1 (g2497), .I2 (I3952));
ND2X1 gate5429(.O (g5779), .I1 (I7549), .I2 (I7550));
ND2X1 gate5430(.O (I7577), .I1 (g84), .I2 (I7576));
ND2X1 gate5431(.O (I5647), .I1 (key_out_111), .I2 (key_out_110));
ND4X1 gate5432(.O (g3531), .I1 (g3209), .I2 (g2215), .I3 (g2976), .I4 (g2179));
ND2X1 gate5433(.O (I1980), .I1 (g230), .I2 (I1978));
ND2X1 gate5434(.O (g5508), .I1 (I7245), .I2 (I7246));
ND2X1 gate5435(.O (I4150), .I1 (g2551), .I2 (g139));
ND2X1 gate5436(.O (g6873), .I1 (g6848), .I2 (g3621));
ND2X1 gate5437(.O (g6095), .I1 (g2952), .I2 (g5854));
ND2X1 gate5438(.O (I4009), .I1 (g292), .I2 (I4008));
ND2X1 gate5439(.O (I2675), .I1 (g710), .I2 (I2674));
ND2X1 gate5440(.O (g926), .I1 (I1952), .I2 (I1953));
ND2X1 gate5441(.O (I3894), .I1 (g286), .I2 (I3893));
ND2X1 gate5442(.O (I4212), .I1 (g804), .I2 (I4210));
ND2X1 gate5443(.O (g5565), .I1 (I7312), .I2 (I7313));
ND2X1 gate5444(.O (I6028), .I1 (g4221), .I2 (I6026));
ND2X1 gate5445(.O (I2109), .I1 (g602), .I2 (I2108));
ND2X1 gate5446(.O (I5244), .I1 (g3247), .I2 (key_out_28));
ND3X1 gate5447(.O (g1402), .I1 (g310), .I2 (g866), .I3 (g873));
ND2X1 gate5448(.O (I4921), .I1 (g650), .I2 (I4919));
ND2X1 gate5449(.O (I7536), .I1 (g5666), .I2 (I7534));
ND2X1 gate5450(.O (I7223), .I1 (g161), .I2 (g5370));
ND2X1 gate5451(.O (I2498), .I1 (key_out_109), .I2 (I2497));
ND2X1 gate5452(.O (I1951), .I1 (g524), .I2 (g248));
ND2X1 gate5453(.O (I7522), .I1 (g5659), .I2 (I7520));
ND2X1 gate5454(.O (I3952), .I1 (g289), .I2 (g2497));
ND2X1 gate5455(.O (g5775), .I1 (I7521), .I2 (I7522));
ND2X1 gate5456(.O (I8201), .I1 (g478), .I2 (g6192));
ND2X1 gate5457(.O (g2024), .I1 (I3126), .I2 (I3127));
ND2X1 gate5458(.O (g2795), .I1 (g1997), .I2 (g866));
ND2X1 gate5459(.O (g4004), .I1 (I5301), .I2 (I5302));
ND2X1 gate5460(.O (I6196), .I1 (g631), .I2 (I6194));
ND2X1 gate5461(.O (I3970), .I1 (g290), .I2 (g2518));
ND2X1 gate5462(.O (I4941), .I1 (g357), .I2 (I4939));
ND2X1 gate5463(.O (I5657), .I1 (key_out_105), .I2 (key_out_104));
ND2X1 gate5464(.O (I7542), .I1 (g59), .I2 (I7541));
ND2X1 gate5465(.O (I2897), .I1 (g1027), .I2 (g634));
ND2X1 gate5466(.O (I2682), .I1 (g918), .I2 (I2681));
ND2X1 gate5467(.O (I2766), .I1 (g749), .I2 (g743));
ND2X1 gate5468(.O (g3013), .I1 (I4211), .I2 (I4212));
ND2X1 gate5469(.O (I5242), .I1 (g3242), .I2 (g3247));
ND2X1 gate5470(.O (I7529), .I1 (g5662), .I2 (I7527));
ND2X1 gate5471(.O (g1822), .I1 (g1070), .I2 (g1084));
ND2X1 gate5472(.O (I3876), .I1 (g2397), .I2 (I3874));
ND2X1 gate5473(.O (I2091), .I1 (g29), .I2 (key_out_23));
ND2X1 gate5474(.O (I3915), .I1 (g287), .I2 (I3914));
ND2X1 gate5475(.O (I9051), .I1 (g6832), .I2 (I9050));
ND2X1 gate5476(.O (I2767), .I1 (g749), .I2 (I2766));
ND2X1 gate5477(.O (I1979), .I1 (g512), .I2 (I1978));
ND2X1 gate5478(.O (g3597), .I1 (I4783), .I2 (I4784));
ND3X1 gate5479(.O (g2831), .I1 (g2007), .I2 (g862), .I3 (g1784));
ND2X1 gate5480(.O (g5683), .I1 (I7433), .I2 (I7434));
ND2X1 gate5481(.O (g5778), .I1 (I7542), .I2 (I7543));
ND2X1 gate5482(.O (I2015), .I1 (g260), .I2 (I2013));
ND2X1 gate5483(.O (g930), .I1 (I1970), .I2 (I1971));
ND2X1 gate5484(.O (g5782), .I1 (I7570), .I2 (I7571));
ND2X1 gate5485(.O (g4002), .I1 (I5293), .I2 (I5294));
ND2X1 gate5486(.O (I2246), .I1 (g598), .I2 (I2244));
ND2X1 gate5487(.O (I6743), .I1 (g4708), .I2 (g582));
ND2X1 gate5488(.O (I7549), .I1 (g64), .I2 (I7548));
ND2X1 gate5489(.O (g2947), .I1 (g1411), .I2 (g2026));
ND2X1 gate5490(.O (g4762), .I1 (I6391), .I2 (key_out_58));
ND3X1 gate5491(.O (g2095), .I1 (g1584), .I2 (g749), .I3 (g736));
ND2X1 gate5492(.O (g944), .I1 (I2004), .I2 (I2005));
ND2X1 gate5493(.O (I6474), .I1 (g4541), .I2 (I6473));
ND2X1 gate5494(.O (I7232), .I1 (g5372), .I2 (I7230));
ND2X1 gate5495(.O (I1953), .I1 (g248), .I2 (I1951));
ND2X1 gate5496(.O (g2719), .I1 (I3875), .I2 (I3876));
ND2X1 gate5497(.O (I8203), .I1 (g6192), .I2 (I8201));
ND2X1 gate5498(.O (I4008), .I1 (g292), .I2 (g2568));
ND2X1 gate5499(.O (g4237), .I1 (g4049), .I2 (g4017));
ND2X1 gate5500(.O (g1829), .I1 (I2898), .I2 (I2899));
ND2X1 gate5501(.O (g901), .I1 (g314), .I2 (g310));
ND2X1 gate5502(.O (g941), .I1 (I1995), .I2 (I1996));
ND2X1 gate5503(.O (I7570), .I1 (g79), .I2 (I7569));
ND2X1 gate5504(.O (I2108), .I1 (g602), .I2 (g610));
ND2X1 gate5505(.O (g1540), .I1 (I2507), .I2 (I2508));
ND4X1 gate5506(.O (g4814), .I1 (g4550), .I2 (g1575), .I3 (g1550), .I4 (g2073));
ND2X1 gate5507(.O (I7311), .I1 (g5364), .I2 (g590));
ND2X1 gate5508(.O (I5270), .I1 (g3705), .I2 (key_out_22));
ND2X1 gate5509(.O (g2745), .I1 (I3915), .I2 (I3916));
ND3X1 gate5510(.O (g1797), .I1 (g98), .I2 (g1064), .I3 (g1070));
ND2X1 gate5511(.O (g2791), .I1 (I3989), .I2 (I3990));
ND2X1 gate5512(.O (I7239), .I1 (g5374), .I2 (I7237));
ND4X1 gate5513(.O (g3526), .I1 (g3196), .I2 (g3023), .I3 (g2197), .I4 (g2981));
ND3X1 gate5514(.O (g6741), .I1 (g6705), .I2 (g6461), .I3 (g4941));
ND2X1 gate5515(.O (I8196), .I1 (g6188), .I2 (I8194));
ND2X1 gate5516(.O (I3895), .I1 (g2422), .I2 (I3893));
ND2X1 gate5517(.O (I4783), .I1 (g2846), .I2 (I4782));
ND2X1 gate5518(.O (I2021), .I1 (g528), .I2 (g254));
ND2X1 gate5519(.O (g905), .I1 (g301), .I2 (g319));
ND2X1 gate5520(.O (g3276), .I1 (I4546), .I2 (I4547));
ND2X1 gate5521(.O (g6774), .I1 (g6754), .I2 (g6750));
ND2X1 gate5522(.O (I5207), .I1 (key_out_2), .I2 (key_out_5));
ND2X1 gate5523(.O (I2301), .I1 (g341), .I2 (I2299));
ND2X1 gate5524(.O (I5259), .I1 (g3719), .I2 (key_out_27));
ND2X1 gate5525(.O (I7440), .I1 (g5515), .I2 (I7439));
ND2X1 gate5526(.O (I7528), .I1 (g49), .I2 (I7527));
ND2X1 gate5527(.O (g4640), .I1 (g4402), .I2 (g1056));
ND4X1 gate5528(.O (g4812), .I1 (g4550), .I2 (g1560), .I3 (g1559), .I4 (g2073));
ND2X1 gate5529(.O (g1845), .I1 (I2934), .I2 (I2935));
ND2X1 gate5530(.O (g6397), .I1 (I8202), .I2 (I8203));
ND2X1 gate5531(.O (I5768), .I1 (g3957), .I2 (key_out_34));
ND2X1 gate5532(.O (I1978), .I1 (g512), .I2 (g230));
ND2X1 gate5533(.O (g4610), .I1 (key_out_75), .I2 (key_out_73));
ND2X1 gate5534(.O (I5228), .I1 (g3263), .I2 (key_out_29));
ND2X1 gate5535(.O (I2074), .I1 (g11), .I2 (key_out_25));
ND3X1 gate5536(.O (g3140), .I1 (g2409), .I2 (g1060), .I3 (g1620));
ND2X1 gate5537(.O (I6390), .I1 (g4504), .I2 (g4610));
ND2X1 gate5538(.O (I3177), .I1 (g1706), .I2 (g736));
ND2X1 gate5539(.O (I4152), .I1 (g139), .I2 (I4150));
ND2X1 gate5540(.O (I6501), .I1 (g3541), .I2 (key_out_91));
ND2X1 gate5541(.O (I7548), .I1 (g64), .I2 (g5672));
ND2X1 gate5542(.O (g1815), .I1 (g102), .I2 (g1070));
ND2X1 gate5543(.O (I7555), .I1 (g69), .I2 (g5674));
ND4X1 gate5544(.O (g3517), .I1 (g3173), .I2 (g3002), .I3 (g2976), .I4 (g2179));
ND2X1 gate5545(.O (I2080), .I1 (g25), .I2 (g19));
ND2X1 gate5546(.O (I4211), .I1 (g2294), .I2 (I4210));
ND2X1 gate5547(.O (I3399), .I1 (g1826), .I2 (I3398));
ND2X1 gate5548(.O (I5195), .I1 (key_out_7), .I2 (key_out_4));
ND2X1 gate5549(.O (I7313), .I1 (g590), .I2 (I7311));
ND2X1 gate5550(.O (g2582), .I1 (I3698), .I2 (I3699));
ND2X1 gate5551(.O (I4939), .I1 (g3437), .I2 (g357));
ND2X1 gate5552(.O (g950), .I1 (I2022), .I2 (I2023));
ND2X1 gate5553(.O (g4819), .I1 (I6500), .I2 (key_out_90));
ND2X1 gate5554(.O (I7521), .I1 (g361), .I2 (I7520));
ND2X1 gate5555(.O (I2023), .I1 (g254), .I2 (I2021));
ND2X1 gate5556(.O (I4446), .I1 (g606), .I2 (I4444));
ND2X1 gate5557(.O (I5783), .I1 (g3810), .I2 (I5782));
ND2X1 gate5558(.O (g2940), .I1 (g197), .I2 (g2381));
ND2X1 gate5559(.O (g4825), .I1 (g4472), .I2 (g4465));
ND2X1 gate5560(.O (I5293), .I1 (g3421), .I2 (I5292));
ND2X1 gate5561(.O (I5761), .I1 (g3503), .I2 (I5759));
ND2X1 gate5562(.O (I1971), .I1 (g236), .I2 (I1969));
ND2X1 gate5563(.O (I3972), .I1 (g2518), .I2 (I3970));
ND2X1 gate5564(.O (I4159), .I1 (g2015), .I2 (g619));
ND2X1 gate5565(.O (I6661), .I1 (g3541), .I2 (key_out_33));
ND2X1 gate5566(.O (g1398), .I1 (g306), .I2 (g889));
ND2X1 gate5567(.O (I6475), .I1 (g578), .I2 (I6473));
ND2X1 gate5568(.O (I3934), .I1 (g288), .I2 (I3933));
ND2X1 gate5569(.O (I7541), .I1 (g59), .I2 (g5669));
ND2X1 gate5570(.O (I2508), .I1 (key_out_106), .I2 (I2506));
ND4X1 gate5571(.O (g5854), .I1 (g5638), .I2 (g1683), .I3 (g1552), .I4 (g2062));
ND2X1 gate5572(.O (g4465), .I1 (g319), .I2 (g4253));
ND2X1 gate5573(.O (I2072), .I1 (g15), .I2 (g11));
ND2X1 gate5574(.O (I7238), .I1 (g179), .I2 (I7237));
ND2X1 gate5575(.O (g3955), .I1 (key_out_60), .I2 (I5189));
ND2X1 gate5576(.O (I7209), .I1 (g143), .I2 (I7208));
ND2X1 gate5577(.O (g5431), .I1 (I7098), .I2 (I7099));
ND2X1 gate5578(.O (I2681), .I1 (g918), .I2 (g613));
ND2X1 gate5579(.O (I2013), .I1 (g532), .I2 (g260));
ND2X1 gate5580(.O (I4234), .I1 (g2267), .I2 (I4233));
ND2X1 gate5581(.O (g2780), .I1 (I3971), .I2 (I3972));
ND2X1 gate5582(.O (g2067), .I1 (I3178), .I2 (I3179));
ND2X1 gate5583(.O (I1962), .I1 (g520), .I2 (I1961));
ND2X1 gate5584(.O (I5258), .I1 (g3714), .I2 (key_out_27));
ND3X1 gate5585(.O (g1387), .I1 (g862), .I2 (g314), .I3 (g301));
ND2X1 gate5586(.O (I2060), .I1 (g7), .I2 (g3));
ND2X1 gate5587(.O (g5781), .I1 (I7563), .I2 (I7564));
ND2X1 gate5588(.O (g2263), .I1 (I3399), .I2 (I3400));
ND2X1 gate5589(.O (g4221), .I1 (I5648), .I2 (I5649));
ND2X1 gate5590(.O (g1359), .I1 (g866), .I2 (g306));
ND2X1 gate5591(.O (I7231), .I1 (g170), .I2 (I7230));
ND2X1 gate5592(.O (I3953), .I1 (g289), .I2 (I3952));
ND2X1 gate5593(.O (I5187), .I1 (key_out_8), .I2 (key_out_6));
ND3X1 gate5594(.O (g5852), .I1 (g5638), .I2 (g2053), .I3 (g1661));
ND4X1 gate5595(.O (g3520), .I1 (g3183), .I2 (g3002), .I3 (g2197), .I4 (g2968));
ND2X1 gate5596(.O (g1047), .I1 (I2090), .I2 (I2091));
ND2X1 gate5597(.O (I7099), .I1 (g574), .I2 (I7097));
ND2X1 gate5598(.O (I3848), .I1 (g2370), .I2 (I3846));
ND2X1 gate5599(.O (I3699), .I1 (g642), .I2 (I3697));
ND2X1 gate5600(.O (I3398), .I1 (g1826), .I2 (g135));
ND2X1 gate5601(.O (I1969), .I1 (g516), .I2 (g236));
ND2X1 gate5602(.O (I5307), .I1 (g478), .I2 (g3512));
ND2X1 gate5603(.O (g3974), .I1 (I5243), .I2 (I5244));
ND2X1 gate5604(.O (I5536), .I1 (g3907), .I2 (I5535));
ND2X1 gate5605(.O (g1417), .I1 (g873), .I2 (g889));
ND2X1 gate5606(.O (I7543), .I1 (g5669), .I2 (I7541));
ND2X1 gate5607(.O (g5943), .I1 (g5818), .I2 (g2940));
ND2X1 gate5608(.O (I7534), .I1 (g54), .I2 (g5666));
ND2X1 gate5609(.O (g4319), .I1 (I5783), .I2 (I5784));
ND2X1 gate5610(.O (I3893), .I1 (g286), .I2 (g2422));
ND2X1 gate5611(.O (g2080), .I1 (I3189), .I2 (I3190));
ND2X1 gate5612(.O (I2683), .I1 (g613), .I2 (I2681));
ND2X1 gate5613(.O (I5537), .I1 (g654), .I2 (I5535));
ND2X1 gate5614(.O (I3170), .I1 (g1534), .I2 (I3168));
ND2X1 gate5615(.O (I3125), .I1 (g1279), .I2 (g1276));
ND2X1 gate5616(.O (I5243), .I1 (g3242), .I2 (key_out_28));
ND2X1 gate5617(.O (I1988), .I1 (g224), .I2 (I1986));
ND2X1 gate5618(.O (I6194), .I1 (g4199), .I2 (g631));
ND2X1 gate5619(.O (g3207), .I1 (I4445), .I2 (I4446));
ND2X1 gate5620(.O (I2526), .I1 (g766), .I2 (g719));
ND2X1 gate5621(.O (g6929), .I1 (g4536), .I2 (g6927));
ND2X1 gate5622(.O (g3215), .I1 (g2340), .I2 (g1402));
ND2X1 gate5623(.O (I3446), .I1 (g1689), .I2 (I3445));
ND2X1 gate5624(.O (I7208), .I1 (g143), .I2 (g5367));
ND2X1 gate5625(.O (g5783), .I1 (I7577), .I2 (I7578));
ND2X1 gate5626(.O (I4545), .I1 (g2853), .I2 (g353));
ND2X1 gate5627(.O (I2004), .I1 (g500), .I2 (I2003));
ND2X1 gate5628(.O (I2527), .I1 (g766), .I2 (I2526));
ND2X1 gate5629(.O (I5649), .I1 (key_out_110), .I2 (I5647));
ND2X1 gate5630(.O (g6778), .I1 (g6762), .I2 (g6758));
ND2X1 gate5631(.O (g1686), .I1 (I2675), .I2 (I2676));
ND2X1 gate5632(.O (g4223), .I1 (I5658), .I2 (I5659));
ND2X1 gate5633(.O (I1996), .I1 (g218), .I2 (I1994));
ND2X1 gate5634(.O (I3447), .I1 (g729), .I2 (I3445));
ND2X1 gate5635(.O (I4204), .I1 (g2255), .I2 (I4203));
ND2X1 gate5636(.O (I3874), .I1 (g285), .I2 (g2397));
ND2X1 gate5637(.O (g2944), .I1 (g269), .I2 (g2381));
ND2X1 gate5638(.O (g1253), .I1 (I2245), .I2 (I2246));
ND3X1 gate5639(.O (g2434), .I1 (g1064), .I2 (g1070), .I3 (g1620));
ND2X1 gate5640(.O (I2299), .I1 (g830), .I2 (g341));
ND3X1 gate5641(.O (g5866), .I1 (g5649), .I2 (g1529), .I3 (g2081));
ND2X1 gate5642(.O (g1687), .I1 (I2682), .I2 (I2683));
ND2X1 gate5643(.O (I3935), .I1 (g2473), .I2 (I3933));
ND2X1 gate5644(.O (g4017), .I1 (g107), .I2 (g3425));
ND2X1 gate5645(.O (I4528), .I1 (g646), .I2 (I4526));
ND2X1 gate5646(.O (I2244), .I1 (key_out_32), .I2 (g598));
ND2X1 gate5647(.O (I4151), .I1 (g2551), .I2 (I4150));
ND2X1 gate5648(.O (I6392), .I1 (g4610), .I2 (key_out_59));
ND2X1 gate5649(.O (I4010), .I1 (g2568), .I2 (I4008));
ND2X1 gate5650(.O (I2082), .I1 (g19), .I2 (key_out_24));
ND4X1 gate5651(.O (g5818), .I1 (g5638), .I2 (g2056), .I3 (g1666), .I4 (g1661));
ND2X1 gate5652(.O (g3979), .I1 (I5258), .I2 (I5259));
ND2X1 gate5653(.O (I6176), .I1 (g4236), .I2 (I6175));
ND2X1 gate5654(.O (I4235), .I1 (g798), .I2 (I4233));
ND2X1 gate5655(.O (I2110), .I1 (g610), .I2 (I2108));
ND2X1 gate5656(.O (I7098), .I1 (g5194), .I2 (I7097));
ND2X1 gate5657(.O (I3456), .I1 (g1691), .I2 (I3455));
ND4X1 gate5658(.O (g5821), .I1 (g5638), .I2 (g2056), .I3 (g1076), .I4 (g1666));
ND2X1 gate5659(.O (I3698), .I1 (g1570), .I2 (I3697));
ND2X1 gate5660(.O (g2995), .I1 (I4183), .I2 (I4184));
ND2X1 gate5661(.O (I6473), .I1 (g4541), .I2 (g578));
ND2X1 gate5662(.O (I5659), .I1 (key_out_104), .I2 (I5657));
ND2X1 gate5663(.O (g5636), .I1 (g5564), .I2 (g4769));
ND2X1 gate5664(.O (I6177), .I1 (g571), .I2 (I6175));
ND2X1 gate5665(.O (I2899), .I1 (g634), .I2 (I2897));
ND2X1 gate5666(.O (I3457), .I1 (g784), .I2 (I3455));
ND2X1 gate5667(.O (I3989), .I1 (g291), .I2 (I3988));
ND2X1 gate5668(.O (I3971), .I1 (g290), .I2 (I3970));
ND2X1 gate5669(.O (I4160), .I1 (g2015), .I2 (I4159));
ND2X1 gate5670(.O (I2089), .I1 (g33), .I2 (g29));
ND2X1 gate5671(.O (g4670), .I1 (g4611), .I2 (g3528));
ND4X1 gate5672(.O (g4813), .I1 (g4550), .I2 (g965), .I3 (g1560), .I4 (g2073));
ND2X1 gate5673(.O (I3740), .I1 (g2021), .I2 (I3739));
ND2X1 gate5674(.O (I8194), .I1 (g471), .I2 (g6188));
ND2X1 gate5675(.O (I5300), .I1 (g471), .I2 (g3505));
ND3X1 gate5676(.O (g3893), .I1 (g3664), .I2 (g3656), .I3 (g3647));
ND2X1 gate5677(.O (g6928), .I1 (g4532), .I2 (g6926));
ND2X1 gate5678(.O (I7578), .I1 (g5680), .I2 (I7576));
ND2X1 gate5679(.O (I7535), .I1 (g54), .I2 (I7534));
ND2X1 gate5680(.O (I1961), .I1 (g520), .I2 (g242));
ND4X1 gate5681(.O (g3544), .I1 (g2594), .I2 (g2215), .I3 (g2197), .I4 (g2179));
ND2X1 gate5682(.O (g6394), .I1 (I8195), .I2 (I8196));
ND2X1 gate5683(.O (I5648), .I1 (key_out_111), .I2 (I5647));
ND2X1 gate5684(.O (I7246), .I1 (g5377), .I2 (I7244));
ND2X1 gate5685(.O (g3756), .I1 (I4940), .I2 (I4941));
ND2X1 gate5686(.O (I2062), .I1 (g3), .I2 (key_out_26));
ND2X1 gate5687(.O (I6195), .I1 (g4199), .I2 (I6194));
ND2X1 gate5688(.O (I7216), .I1 (g152), .I2 (g5368));
ND4X1 gate5689(.O (g3536), .I1 (g3219), .I2 (g2215), .I3 (g3007), .I4 (g2179));
ND2X1 gate5690(.O (I7564), .I1 (g5676), .I2 (I7562));
ND2X1 gate5691(.O (g4300), .I1 (I5760), .I2 (I5761));
ND2X1 gate5692(.O (I4184), .I1 (g749), .I2 (I4182));
ND2X1 gate5693(.O (I2005), .I1 (g212), .I2 (I2003));
ND2X1 gate5694(.O (g5318), .I1 (key_out_112), .I2 (g5060));
ND4X1 gate5695(.O (g5872), .I1 (g5649), .I2 (g1557), .I3 (g1564), .I4 (g2113));
NR2X1 gate5696(.O (g5552), .I1 (g5354), .I2 (g5356));
NR2X1 gate5697(.O (g4235), .I1 (g3780), .I2 (g3362));
NR2X1 gate5698(.O (g6073), .I1 (g197), .I2 (g5862));
NR2X1 gate5699(.O (g4776), .I1 (g4449), .I2 (g4453));
NR2X1 gate5700(.O (g4777), .I1 (g4457), .I2 (g4459));
NR2X1 gate5701(.O (g4238), .I1 (g3755), .I2 (g3279));
NR4X1 gate5702(.O (g6433), .I1 (g6385), .I2 (g3733), .I3 (g4092), .I4 (g4314));
NR2X1 gate5703(.O (g6496), .I1 (g952), .I2 (g6354));
NR2X1 gate5704(.O (g1422), .I1 (g1039), .I2 (g913));
NR2X1 gate5705(.O (g3931), .I1 (g3353), .I2 (g3361));
NR2X1 gate5706(.O (g1560), .I1 (g996), .I2 (g980));
NR2X1 gate5707(.O (g3905), .I1 (g3512), .I2 (g478));
NR2X1 gate5708(.O (g5094), .I1 (g4685), .I2 (g4686));
NR2X1 gate5709(.O (g3973), .I1 (g3368), .I2 (g3374));
NR2X1 gate5710(.O (g3528), .I1 (g1802), .I2 (g3167));
NR2X1 gate5711(.O (g5541), .I1 (g5388), .I2 (g1880));
NR2X1 gate5712(.O (g3621), .I1 (g1407), .I2 (g2842));
NR2X1 gate5713(.O (g1449), .I1 (g489), .I2 (g1048));
NR2X1 gate5714(.O (g3965), .I1 (g3359), .I2 (g3367));
NR2X1 gate5715(.O (g3933), .I1 (g3327), .I2 (g3336));
NR4X1 gate5716(.O (g6280), .I1 (I7978), .I2 (I7979), .I3 (I7980), .I4 (I7981));
NR2X1 gate5717(.O (g2433), .I1 (g1418), .I2 (g1449));
NR3X1 gate5718(.O (g1470), .I1 (g937), .I2 (g930), .I3 (g928));
NR4X1 gate5719(.O (g6427), .I1 (g6376), .I2 (g4086), .I3 (g4074), .I4 (g4068));
NR4X1 gate5720(.O (g6446), .I1 (g6385), .I2 (g4334), .I3 (g4092), .I4 (g4314));
NR4X1 gate5721(.O (g6359), .I1 (I8135), .I2 (I8136), .I3 (I8137), .I4 (I8138));
NR3X1 gate5722(.O (g1459), .I1 (g926), .I2 (g950), .I3 (g948));
NR2X1 gate5723(.O (g4584), .I1 (g4164), .I2 (g4168));
NR2X1 gate5724(.O (g3926), .I1 (g3338), .I2 (g3350));
NR4X1 gate5725(.O (g6279), .I1 (I7969), .I2 (I7970), .I3 (I7971), .I4 (I7972));
NR2X1 gate5726(.O (g5265), .I1 (g4863), .I2 (g4865));
NR2X1 gate5727(.O (g3927), .I1 (g3382), .I2 (g3383));
NR2X1 gate5728(.O (g3903), .I1 (g3505), .I2 (g471));
NR2X1 gate5729(.O (g1418), .I1 (g486), .I2 (g943));
NR2X1 gate5730(.O (g4578), .I1 (g4234), .I2 (g3928));
NR2X1 gate5731(.O (g4261), .I1 (g3762), .I2 (g3295));
NR4X1 gate5732(.O (g6358), .I1 (I8126), .I2 (I8127), .I3 (I8128), .I4 (I8129));
NR2X1 gate5733(.O (g4589), .I1 (g4180), .I2 (g4183));
NR2X1 gate5734(.O (g1474), .I1 (g760), .I2 (g754));
NR2X1 gate5735(.O (g3956), .I1 (g3337), .I2 (g3349));
NR2X1 gate5736(.O (g4774), .I1 (g4442), .I2 (g4445));
NR2X1 gate5737(.O (g5091), .I1 (g4698), .I2 (g4701));
NR2X1 gate5738(.O (g4950), .I1 (g1472), .I2 (g4680));
NR2X1 gate5739(.O (g5227), .I1 (g5019), .I2 (key_out_9));
NR2X1 gate5740(.O (g4585), .I1 (g4171), .I2 (g4177));
NR2X1 gate5741(.O (g6494), .I1 (g952), .I2 (g6348));
NR3X1 gate5742(.O (g5048), .I1 (g4819), .I2 (key_out_10), .I3 (key_out_9));
NR3X1 gate5743(.O (g3664), .I1 (g2804), .I2 (g2791), .I3 (g2780));
NR2X1 gate5744(.O (g4000), .I1 (g1250), .I2 (g3425));
NR2X1 gate5745(.O (g5418), .I1 (g5162), .I2 (g5169));
NR2X1 gate5746(.O (g5093), .I1 (g4683), .I2 (g4684));
NR2X1 gate5747(.O (g4779), .I1 (g4461), .I2 (g4464));
NR2X1 gate5748(.O (g6492), .I1 (g6348), .I2 (g1734));
NR3X1 gate5749(.O (g4240), .I1 (g1589), .I2 (g1879), .I3 (g3793));
NR2X1 gate5750(.O (g4596), .I1 (g4184), .I2 (g4186));
NR2X1 gate5751(.O (g1603), .I1 (g1039), .I2 (g658));
NR3X1 gate5752(.O (g2908), .I1 (g536), .I2 (g2010), .I3 (g541));
NR2X1 gate5753(.O (g4581), .I1 (g4156), .I2 (g4160));
NR2X1 gate5754(.O (g5423), .I1 (g5170), .I2 (g5175));
NR2X1 gate5755(.O (g4432), .I1 (g923), .I2 (g4253));
NR4X1 gate5756(.O (g6436), .I1 (g6385), .I2 (g3733), .I3 (g4328), .I4 (g4080));
NR2X1 gate5757(.O (g4568), .I1 (g4233), .I2 (g3924));
NR4X1 gate5758(.O (g6335), .I1 (I8079), .I2 (I8080), .I3 (I8081), .I4 (I8082));
NR2X1 gate5759(.O (g5753), .I1 (g1477), .I2 (g5688));
NR2X1 gate5760(.O (g6495), .I1 (g6354), .I2 (g1775));
NR4X1 gate5761(.O (g6442), .I1 (g6376), .I2 (g4323), .I3 (g4074), .I4 (g4302));
NR4X1 gate5762(.O (g6429), .I1 (g6376), .I2 (g4086), .I3 (g4074), .I4 (g4302));
NR4X1 gate5763(.O (g6281), .I1 (I7987), .I2 (I7988), .I3 (I7989), .I4 (I7990));
NR4X1 gate5764(.O (g6449), .I1 (g6385), .I2 (g4334), .I3 (g4328), .I4 (g4080));
NR2X1 gate5765(.O (g4590), .I1 (g4169), .I2 (g4172));
NR2X1 gate5766(.O (g4877), .I1 (g952), .I2 (g4680));
NR4X1 gate5767(.O (g6445), .I1 (g6376), .I2 (g4323), .I3 (g4309), .I4 (g4068));
NR4X1 gate5768(.O (g5561), .I1 (g5391), .I2 (g1589), .I3 (g3793), .I4 (g1880));
NR2X1 gate5769(.O (g3929), .I1 (g3373), .I2 (g3376));
NR3X1 gate5770(.O (g1473), .I1 (g944), .I2 (g941), .I3 (g939));
NR2X1 gate5771(.O (g4967), .I1 (g4674), .I2 (g952));
NR4X1 gate5772(.O (g6430), .I1 (g6385), .I2 (g3733), .I3 (g4092), .I4 (g4080));
NR2X1 gate5773(.O (g4993), .I1 (g4674), .I2 (g1477));
NR4X1 gate5774(.O (g6448), .I1 (g6376), .I2 (g4323), .I3 (g4309), .I4 (g4302));
NR3X1 gate5775(.O (g3647), .I1 (g2731), .I2 (g2719), .I3 (g2698));
NR2X1 gate5776(.O (g3925), .I1 (g3303), .I2 (g3315));
NR2X1 gate5777(.O (g5731), .I1 (g952), .I2 (g5688));
NR2X1 gate5778(.O (g3959), .I1 (g3352), .I2 (g3360));
NR2X1 gate5779(.O (g1481), .I1 (g815), .I2 (g809));
NR3X1 gate5780(.O (g3656), .I1 (g2769), .I2 (g2757), .I3 (g2745));
NR2X1 gate5781(.O (g4245), .I1 (g3759), .I2 (g3288));
NR2X1 gate5782(.O (g3930), .I1 (g3317), .I2 (g3328));
NR2X1 gate5783(.O (g5249), .I1 (g4868), .I2 (g4870));
NR2X1 gate5784(.O (g3966), .I1 (g3329), .I2 (g3339));
NR4X1 gate5785(.O (g6400), .I1 (I8208), .I2 (I8209), .I3 (I8210), .I4 (I8211));
NR2X1 gate5786(.O (g4266), .I1 (g3757), .I2 (g3283));
NR4X1 gate5787(.O (g6451), .I1 (g6385), .I2 (g4334), .I3 (g4328), .I4 (g4314));
NR3X1 gate5788(.O (g5324), .I1 (g5069), .I2 (g4410), .I3 (g766));
NR4X1 gate5789(.O (g6443), .I1 (g6385), .I2 (g4334), .I3 (g4092), .I4 (g4080));
NR2X1 gate5790(.O (g5088), .I1 (g4691), .I2 (g4697));
NR2X1 gate5791(.O (g3958), .I1 (g3316), .I2 (g3326));
NR2X1 gate5792(.O (g4241), .I1 (g3774), .I2 (g3341));
NR4X1 gate5793(.O (g6432), .I1 (g6376), .I2 (g4086), .I3 (g4309), .I4 (g4068));
NR4X1 gate5794(.O (g6357), .I1 (I8117), .I2 (I8118), .I3 (I8119), .I4 (I8120));
NR2X1 gate5795(.O (g3923), .I1 (g3378), .I2 (g3381));
NR2X1 gate5796(.O (g6075), .I1 (g269), .I2 (g5863));
NR2X1 gate5797(.O (g3934), .I1 (g3377), .I2 (g3379));
NR4X1 gate5798(.O (g6439), .I1 (g6385), .I2 (g3733), .I3 (g4328), .I4 (g4314));
NR2X1 gate5799(.O (g4272), .I1 (g3767), .I2 (g3319));
NR2X1 gate5800(.O (g1879), .I1 (g1603), .I2 (g1416));
NR3X1 gate5801(.O (g5325), .I1 (g5077), .I2 (g4416), .I3 (g821));
NR4X1 gate5802(.O (g6435), .I1 (g6376), .I2 (g4086), .I3 (g4309), .I4 (g4302));
NR2X1 gate5803(.O (g4586), .I1 (g4161), .I2 (g4165));
NR2X1 gate5804(.O (g3939), .I1 (g3340), .I2 (g3351));
NR4X1 gate5805(.O (g6438), .I1 (g6376), .I2 (g4323), .I3 (g4074), .I4 (g4068));
NR2X1 gate5806(.O (g1518), .I1 (g980), .I2 (g965));
NR2X1 gate5807(.O (g4239), .I1 (g3763), .I2 (g3296));
NR2X1 gate5808(.O (g4591), .I1 (g4178), .I2 (g4181));
endmodule