
module s5378_0 ( clk, n3065gat, n3066gat, n3067gat, n3068gat, n3069gat, 
        n3070gat, n3071gat, n3072gat, n3073gat, n3074gat, n3075gat, n3076gat, 
        n3077gat, n3078gat, n3079gat, n3080gat, n3081gat, n3082gat, n3083gat, 
        n3084gat, n3085gat, n3086gat, n3087gat, n3088gat, n3089gat, n3090gat, 
        n3091gat, n3092gat, n3093gat, n3094gat, n3095gat, n3097gat, n3098gat, 
        n3099gat, n3100gat, n3104gat, n3105gat, n3106gat, n3107gat, n3108gat, 
        n3109gat, n3110gat, n3111gat, n3112gat, n3113gat, n3114gat, n3115gat, 
        n3116gat, n3117gat, n3118gat, n3119gat, n3120gat, n3121gat, n3122gat, 
        n3123gat, n3124gat, n3125gat, n3126gat, n3127gat, n3128gat, n3129gat, 
        n3130gat, n3131gat, n3132gat, n3133gat, n3134gat, n3135gat, n3136gat, 
        n3137gat, n3138gat, n3139gat, n3140gat, n3141gat, n3142gat, n3143gat, 
        n3144gat, n3145gat, n3146gat, n3147gat, n3148gat, n3149gat, n3150gat, 
        n3151gat, n3152gat, test_si, test_so, test_se );
  input clk, n3065gat, n3066gat, n3067gat, n3068gat, n3069gat, n3070gat,
         n3071gat, n3072gat, n3073gat, n3074gat, n3075gat, n3076gat, n3077gat,
         n3078gat, n3079gat, n3080gat, n3081gat, n3082gat, n3083gat, n3084gat,
         n3085gat, n3086gat, n3087gat, n3088gat, n3089gat, n3090gat, n3091gat,
         n3092gat, n3093gat, n3094gat, n3095gat, n3097gat, n3098gat, n3099gat,
         n3100gat, test_si, test_se;
  output n3104gat, n3105gat, n3106gat, n3107gat, n3108gat, n3109gat, n3110gat,
         n3111gat, n3112gat, n3113gat, n3114gat, n3115gat, n3116gat, n3117gat,
         n3118gat, n3119gat, n3120gat, n3121gat, n3122gat, n3123gat, n3124gat,
         n3125gat, n3126gat, n3127gat, n3128gat, n3129gat, n3130gat, n3131gat,
         n3132gat, n3133gat, n3134gat, n3135gat, n3136gat, n3137gat, n3138gat,
         n3139gat, n3140gat, n3141gat, n3142gat, n3143gat, n3144gat, n3145gat,
         n3146gat, n3147gat, n3148gat, n3149gat, n3150gat, n3151gat, n3152gat,
         test_so;
  wire   n2522gat, n1821gat, n2476gat, n2468gat, n2526gat, n2464gat, n2102gat,
         n1763gat, n1197gat, n667gat, n1834gat, n1767gat, n2021gat, n2182gat,
         n2040gat, n2266gat, n1975gat, n470gat, n148gat, n1771gat, n1525gat,
         n2897gat, n748gat, n43gat, n55gat, n2914gat, n2928gat, n2927gat,
         n2896gat, n2922gat, n2894gat, n2921gat, n2895gat, n933gat, n504gat,
         n2913gat, n2920gat, n2905gat, n2898gat, n567gat, n2989gat, n2918gat,
         n2952gat, n2919gat, n2910gat, n2907gat, n2911gat, n2912gat, n2909gat,
         n2908gat, n2971gat, n2904gat, n2891gat, n2903gat, n2915gat, n2901gat,
         n2890gat, n2888gat, n2887gat, n2886gat, n3010gat, n3016gat, n2579gat,
         n2613gat, n2983gat, n2917gat, n2892gat, n2900gat, n2929gat, n2925gat,
         n2916gat, n2899gat, n2926gat, n2924gat, n2923gat, n3147gat, n3142gat,
         n1620gat, n1827gat, n1606gat, n1610gat, n1793gat, n1516gat, n1565gat,
         n1696gat, n2009gat, n1636gat, n2163gat, n2015gat, n2017gat, n2194gat,
         n2057gat, n2556gat, n2436gat, n2387gat, n2330gat, n2396gat, n2198gat,
         n2197gat, n2196gat, n1882gat, n1613gat, n1391gat, n1927gat, n1567gat,
         n1564gat, n1915gat, n1800gat, n1593gat, n185, n186, n188, n189, n190,
         n195, n196, n197, n231, n232, n244, n568, n569, n572, n576, n587,
         n588, n606, n608, n651, n657, n667, n3139gat, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n699, n700, n704, n705, n706, n707, n708, n709, n711,
         n712, n713, n715, n717, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248;
  assign n3152gat = n3147gat;
  assign n3112gat = n3147gat;
  assign n3115gat = n3147gat;
  assign n3148gat = n3147gat;
  assign n3141gat = n3142gat;
  assign n3140gat = n3139gat;

  DFZX1 gate1 ( .D(n2897gat), .TD(test_si), .SEL(test_se), .CK(clk), .Q(n1248), 
        .QB(n737) );
  DFZX1 gate2 ( .D(n3069gat), .TD(n1248), .SEL(test_se), .CK(clk), .Q(n1160)
         );
  DFZX1 gate3 ( .D(n3070gat), .TD(n1160), .SEL(test_se), .CK(clk), .Q(n1146), 
        .QB(n751) );
  DFZX1 gate4 ( .D(n3072gat), .TD(n1146), .SEL(test_se), .CK(clk), .Q(n1144)
         );
  DFZX1 gate5 ( .D(n3071gat), .TD(n1144), .SEL(test_se), .CK(clk), .Q(n1145)
         );
  DFZX1 gate6 ( .D(n3069gat), .TD(n1145), .SEL(test_se), .CK(clk), .Q(n1159), 
        .QB(n731) );
  DFZX1 gate7 ( .D(n3070gat), .TD(n1159), .SEL(test_se), .CK(clk), .Q(n1161), 
        .QB(n747) );
  DFZX1 gate8 ( .D(n3072gat), .TD(n1161), .SEL(test_se), .CK(clk), .Q(n1162), 
        .QB(n746) );
  DFZX1 gate9 ( .D(n3071gat), .TD(n1162), .SEL(test_se), .CK(clk), .Q(n1163), 
        .QB(n736) );
  DFZX1 gate10 ( .D(n748gat), .TD(n1163), .SEL(test_se), .CK(clk), .Q(n1247), 
        .QB(n657) );
  DFZX1 gate11 ( .D(n3065gat), .TD(n1247), .SEL(test_se), .CK(clk), .Q(n1143), 
        .QB(n757) );
  DFZX1 gate12 ( .D(n3067gat), .TD(n1143), .SEL(test_se), .CK(clk), .Q(n1123)
         );
  DFZX1 gate13 ( .D(n3066gat), .TD(n1123), .SEL(test_se), .CK(clk), .Q(n1125)
         );
  DFZX1 gate14 ( .D(n3073gat), .TD(n1125), .SEL(test_se), .CK(clk), .Q(n1164), 
        .QB(n753) );
  DFZX1 gate15 ( .D(n3068gat), .TD(n1164), .SEL(test_se), .CK(clk), .Q(n1122)
         );
  DFZX1 gate16 ( .D(n43gat), .TD(n1122), .SEL(test_se), .CK(clk), .Q(n2522gat)
         );
  DFZX1 gate17 ( .D(n1620gat), .TD(n2522gat), .SEL(test_se), .CK(clk), .Q(
        n1140), .QB(n675) );
  DFZX1 gate18 ( .D(n675), .TD(n1140), .SEL(test_se), .CK(clk), .Q(n1246), 
        .QB(n651) );
  DFZX1 gate19 ( .D(n1827gat), .TD(n1246), .SEL(test_se), .CK(clk), .Q(
        n1821gat) );
  DFZX1 gate20 ( .D(n1827gat), .TD(n1821gat), .SEL(test_se), .CK(clk), .Q(
        n1142), .QB(n758) );
  DFZX1 gate21 ( .D(n676), .TD(n1142), .SEL(test_se), .CK(clk), .Q(n1245), 
        .QB(n677) );
  DFZX1 gate22 ( .D(n677), .TD(n1245), .SEL(test_se), .CK(clk), .Q(n1141) );
  DFZX1 gate23 ( .D(n3065gat), .TD(n1141), .SEL(test_se), .CK(clk), .Q(n1244), 
        .QB(n732) );
  DFZX1 gate24 ( .D(n3067gat), .TD(n1244), .SEL(test_se), .CK(clk), .Q(n1105), 
        .QB(n756) );
  DFZX1 gate25 ( .D(n3066gat), .TD(n1105), .SEL(test_se), .CK(clk), .Q(n1165)
         );
  DFZX1 gate26 ( .D(n3073gat), .TD(n1165), .SEL(test_se), .CK(clk), .Q(n1101)
         );
  DFZX1 gate27 ( .D(n3068gat), .TD(n1101), .SEL(test_se), .CK(clk), .Q(n1166)
         );
  DFZX1 gate28 ( .D(n55gat), .TD(n1166), .SEL(test_se), .CK(clk), .Q(n2476gat)
         );
  DFZX1 gate29 ( .D(n2914gat), .TD(n2476gat), .SEL(test_se), .CK(clk), .Q(
        n1211), .QB(n740) );
  DFZX1 gate30 ( .D(n2928gat), .TD(n1211), .SEL(test_se), .CK(clk), .Q(n1108), 
        .QB(n755) );
  DFZX1 gate31 ( .D(n2927gat), .TD(n1108), .SEL(test_se), .CK(clk), .Q(n1167)
         );
  DFZX1 gate32 ( .D(n2896gat), .TD(n1167), .SEL(test_se), .CK(clk), .Q(n1212)
         );
  DFZX1 gate33 ( .D(n2922gat), .TD(n1212), .SEL(test_se), .CK(clk), .Q(n1213)
         );
  DFZX1 gate34 ( .D(n2897gat), .TD(n1213), .SEL(test_se), .CK(clk), .Q(n1111)
         );
  DFZX1 gate35 ( .D(n2894gat), .TD(n1111), .SEL(test_se), .CK(clk), .Q(n1168)
         );
  DFZX1 gate36 ( .D(n2921gat), .TD(n1168), .SEL(test_se), .CK(clk), .Q(n1169)
         );
  DFZX1 gate37 ( .D(n2895gat), .TD(n1169), .SEL(test_se), .CK(clk), .Q(n1109), 
        .QB(n739) );
  DFZX1 gate38 ( .D(n933gat), .TD(n1109), .SEL(test_se), .CK(clk), .Q(n2468gat) );
  DFZX1 gate39 ( .D(n3070gat), .TD(n2468gat), .SEL(test_se), .CK(clk), .Q(
        n1205) );
  DFZX1 gate40 ( .D(n3069gat), .TD(n1205), .SEL(test_se), .CK(clk), .Q(n1206)
         );
  DFZX1 gate41 ( .D(n3071gat), .TD(n1206), .SEL(test_se), .CK(clk), .Q(n1207)
         );
  DFZX1 gate42 ( .D(n3072gat), .TD(n1207), .SEL(test_se), .CK(clk), .Q(n1100)
         );
  DFZX1 gate43 ( .D(n2923gat), .TD(n1100), .SEL(test_se), .CK(clk), .Q(n1106), 
        .QB(n678) );
  DFZX1 gate44 ( .D(n2917gat), .TD(n1106), .SEL(test_se), .CK(clk), .Q(n1104), 
        .QB(n679) );
  DFZX1 gate45 ( .D(n2924gat), .TD(n1104), .SEL(test_se), .CK(clk), .Q(n1170), 
        .QB(n680) );
  DFZX1 gate46 ( .D(n2926gat), .TD(n1170), .SEL(test_se), .CK(clk), .Q(n1099), 
        .QB(n681) );
  DFZX1 gate47 ( .D(n2892gat), .TD(n1099), .SEL(test_se), .CK(clk), .Q(n1171), 
        .QB(n682) );
  DFZX1 gate48 ( .D(n504gat), .TD(n1171), .SEL(test_se), .CK(clk), .Q(n2526gat) );
  DFZX1 gate49 ( .D(n2913gat), .TD(n2526gat), .SEL(test_se), .CK(clk), .Q(
        n1208), .QB(n754) );
  DFZX1 gate50 ( .D(n2920gat), .TD(n1208), .SEL(test_se), .CK(clk), .Q(n1107), 
        .QB(n738) );
  DFZX1 gate51 ( .D(n2905gat), .TD(n1107), .SEL(test_se), .CK(clk), .Q(n1172)
         );
  DFZX1 gate52 ( .D(n2900gat), .TD(n1172), .SEL(test_se), .CK(clk), .Q(n1209), 
        .QB(n683) );
  DFZX1 gate53 ( .D(n2925gat), .TD(n1209), .SEL(test_se), .CK(clk), .Q(n1210), 
        .QB(n684) );
  DFZX1 gate54 ( .D(n2929gat), .TD(n1210), .SEL(test_se), .CK(clk), .Q(n1112), 
        .QB(n685) );
  DFZX1 gate55 ( .D(n2898gat), .TD(n1112), .SEL(test_se), .CK(clk), .Q(n1173)
         );
  DFZX1 gate56 ( .D(n2916gat), .TD(n1173), .SEL(test_se), .CK(clk), .Q(n1174), 
        .QB(n686) );
  DFZX1 gate57 ( .D(n2899gat), .TD(n1174), .SEL(test_se), .CK(clk), .Q(n1110), 
        .QB(n687) );
  DFZX1 gate58 ( .D(n567gat), .TD(n1110), .SEL(test_se), .CK(clk), .Q(n2464gat) );
  DFZX1 gate59 ( .D(n2396gat), .TD(n2464gat), .SEL(test_se), .CK(clk), .Q(
        n1175), .QB(n688) );
  DFZX1 gate60 ( .D(n2198gat), .TD(n1175), .SEL(test_se), .CK(clk), .Q(n1176), 
        .QB(n689) );
  DFZX1 gate61 ( .D(n2196gat), .TD(n1176), .SEL(test_se), .CK(clk), .Q(n1177), 
        .QB(n690) );
  DFZX1 gate62 ( .D(n196), .TD(n1177), .SEL(test_se), .CK(clk), .Q(n1178), 
        .QB(n691) );
  DFZX1 gate63 ( .D(n2197gat), .TD(n1178), .SEL(test_se), .CK(clk), .Q(n1179), 
        .QB(n692) );
  DFZX1 gate64 ( .D(n195), .TD(n1179), .SEL(test_se), .CK(clk), .Q(n1151), 
        .QB(n693) );
  DFZX1 gate65 ( .D(n2330gat), .TD(n1151), .SEL(test_se), .CK(clk), .Q(n1180), 
        .QB(n694) );
  DFZX1 gate66 ( .D(n2387gat), .TD(n1180), .SEL(test_se), .CK(clk), .Q(n1181), 
        .QB(n695) );
  DFZX1 gate67 ( .D(n2556gat), .TD(n1181), .SEL(test_se), .CK(clk), .Q(n1214), 
        .QB(n696) );
  DFZX1 gate68 ( .D(n2436gat), .TD(n1214), .SEL(test_se), .CK(clk), .Q(n1215), 
        .QB(n697) );
  DFZX1 gate69 ( .D(n1606gat), .TD(n1215), .SEL(test_se), .CK(clk), .Q(
        n2102gat) );
  DFZX1 gate70 ( .D(n1882gat), .TD(n2102gat), .SEL(test_se), .CK(clk), .Q(
        n1182) );
  DFZX1 gate71 ( .D(n1610gat), .TD(n1182), .SEL(test_se), .CK(clk), .Q(
        n1763gat) );
  DFZX1 gate72 ( .D(n2989gat), .TD(n1763gat), .SEL(test_se), .CK(clk), .Q(
        n1183) );
  DFZX1 gate73 ( .D(n2918gat), .TD(n1183), .SEL(test_se), .CK(clk), .Q(n1184), 
        .QB(n752) );
  DFZX1 gate74 ( .D(n2952gat), .TD(n1184), .SEL(test_se), .CK(clk), .Q(n1156)
         );
  DFZX1 gate75 ( .D(n2919gat), .TD(n1156), .SEL(test_se), .CK(clk), .Q(n1157)
         );
  DFZX1 gate76 ( .D(n2910gat), .TD(n1157), .SEL(test_se), .CK(clk), .Q(n1158)
         );
  DFZX1 gate77 ( .D(n2907gat), .TD(n1158), .SEL(test_se), .CK(clk), .Q(n1154)
         );
  DFZX1 gate78 ( .D(n2911gat), .TD(n1154), .SEL(test_se), .CK(clk), .Q(n1155)
         );
  DFZX1 gate79 ( .D(n2912gat), .TD(n1155), .SEL(test_se), .CK(clk), .Q(n1152)
         );
  DFZX1 gate80 ( .D(n2909gat), .TD(n1152), .SEL(test_se), .CK(clk), .Q(n1153)
         );
  DFZX1 gate81 ( .D(n2908gat), .TD(n1153), .SEL(test_se), .CK(clk), .Q(
        n1197gat) );
  DFZX1 gate82 ( .D(n2971gat), .TD(n1197gat), .SEL(test_se), .CK(clk), .Q(
        n1243), .QB(n1090) );
  DFZX1 gate83 ( .D(n2904gat), .TD(n1243), .SEL(test_se), .CK(clk), .Q(n667gat) );
  DFZX1 gate84 ( .D(n2891gat), .TD(n667gat), .SEL(test_se), .CK(clk), .Q(n1185) );
  DFZX1 gate85 ( .D(n2903gat), .TD(n1185), .SEL(test_se), .CK(clk), .Q(n1120)
         );
  DFZX1 gate86 ( .D(n2915gat), .TD(n1120), .SEL(test_se), .CK(clk), .Q(n1124)
         );
  DFZX1 gate87 ( .D(n2901gat), .TD(n1124), .SEL(test_se), .CK(clk), .Q(n1121)
         );
  DFZX1 gate88 ( .D(n2890gat), .TD(n1121), .SEL(test_se), .CK(clk), .Q(n1118), 
        .QB(n759) );
  DFZX1 gate89 ( .D(n2888gat), .TD(n1118), .SEL(test_se), .CK(clk), .Q(n1119)
         );
  DFZX1 gate90 ( .D(n2887gat), .TD(n1119), .SEL(test_se), .CK(clk), .Q(n1116)
         );
  DFZX1 gate91 ( .D(n2886gat), .TD(n1116), .SEL(test_se), .CK(clk), .Q(n1117)
         );
  DFZX1 gate92 ( .D(n3010gat), .TD(n1117), .SEL(test_se), .CK(clk), .Q(n1089)
         );
  DFZX1 gate93 ( .D(n3016gat), .TD(n1089), .SEL(test_se), .CK(clk), .Q(n1242), 
        .QB(n608) );
  DFZX1 gate94 ( .D(n672), .TD(n1242), .SEL(test_se), .CK(clk), .Q(n1129), 
        .QB(n699) );
  DFZX1 gate95 ( .D(n2579gat), .TD(n1129), .SEL(test_se), .CK(clk), .Q(n1241), 
        .QB(n1137) );
  DFZX1 gate96 ( .D(n674), .TD(n1241), .SEL(test_se), .CK(clk), .Q(n1127), 
        .QB(n700) );
  DFZX1 gate97 ( .D(n197), .TD(n1127), .SEL(test_se), .CK(clk), .Q(n1126), 
        .QB(n3128gat) );
  DFZX1 gate98 ( .D(n2194gat), .TD(n1126), .SEL(test_se), .CK(clk), .Q(n1128), 
        .QB(n3127gat) );
  DFZX1 gate99 ( .D(n2057gat), .TD(n1128), .SEL(test_se), .CK(clk), .Q(n1240), 
        .QB(n3126gat) );
  DFZX1 gate100 ( .D(n231), .TD(n1240), .SEL(test_se), .CK(clk), .Q(n1138) );
  DFZX1 gate101 ( .D(n673), .TD(n1138), .SEL(test_se), .CK(clk), .Q(n1239), 
        .QB(n704) );
  DFZX1 gate102 ( .D(n2613gat), .TD(n1239), .SEL(test_se), .CK(clk), .Q(n1238), 
        .QB(n606) );
  DFZX1 gate103 ( .D(n188), .TD(n1238), .SEL(test_se), .CK(clk), .Q(n1834gat)
         );
  DFZX1 gate104 ( .D(n189), .TD(n1834gat), .SEL(test_se), .CK(clk), .Q(
        n1767gat) );
  DFZX1 gate105 ( .D(n3149gat), .TD(n1767gat), .SEL(test_se), .CK(clk), .Q(
        n1103) );
  DFZX1 gate106 ( .D(n697), .TD(n1103), .SEL(test_se), .CK(clk), .Q(n1147), 
        .QB(n744) );
  DFZX1 gate107 ( .D(n695), .TD(n1147), .SEL(test_se), .CK(clk), .Q(n1186), 
        .QB(n748) );
  DFZX1 gate108 ( .D(n694), .TD(n1186), .SEL(test_se), .CK(clk), .Q(n1150), 
        .QB(n734) );
  DFZX1 gate109 ( .D(n693), .TD(n1150), .SEL(test_se), .CK(clk), .Q(n1148), 
        .QB(n741) );
  DFZX1 gate110 ( .D(n696), .TD(n1148), .SEL(test_se), .CK(clk), .Q(n1149), 
        .QB(n735) );
  DFZX1 gate111 ( .D(n688), .TD(n1149), .SEL(test_se), .CK(clk), .Q(n1187), 
        .QB(n743) );
  DFZX1 gate112 ( .D(n689), .TD(n1187), .SEL(test_se), .CK(clk), .Q(n1188), 
        .QB(n745) );
  DFZX1 gate113 ( .D(n691), .TD(n1188), .SEL(test_se), .CK(clk), .Q(n1189), 
        .QB(n730) );
  DFZX1 gate114 ( .D(n692), .TD(n1189), .SEL(test_se), .CK(clk), .Q(n1190), 
        .QB(n742) );
  DFZX1 gate115 ( .D(n690), .TD(n1190), .SEL(test_se), .CK(clk), .Q(n1191), 
        .QB(n733) );
  DFZX1 gate116 ( .D(n1793gat), .TD(n1191), .SEL(test_se), .CK(clk), .Q(n1237), 
        .QB(n1102) );
  DFZX1 gate117 ( .D(n670), .TD(n1237), .SEL(test_se), .CK(clk), .Q(n2021gat)
         );
  DFZX1 gate118 ( .D(n1516gat), .TD(n2021gat), .SEL(test_se), .CK(clk), .Q(
        n1113), .QB(n708) );
  DFZX1 gate119 ( .D(n708), .TD(n1113), .SEL(test_se), .CK(clk), .Q(n1131) );
  DFZX1 gate120 ( .D(n186), .TD(n1131), .SEL(test_se), .CK(clk), .Q(n1130) );
  DFZX1 gate121 ( .D(n1565gat), .TD(n1130), .SEL(test_se), .CK(clk), .Q(n1236), 
        .QB(n709) );
  DFZX1 gate122 ( .D(n709), .TD(n1236), .SEL(test_se), .CK(clk), .Q(n1192) );
  DFZX1 gate123 ( .D(n190), .TD(n1192), .SEL(test_se), .CK(clk), .Q(n1235), 
        .QB(n1091) );
  DFZX1 gate124 ( .D(n3127gat), .TD(n1235), .SEL(test_se), .CK(clk), .Q(n1193)
         );
  DFZX1 gate125 ( .D(n3126gat), .TD(n1193), .SEL(test_se), .CK(clk), .Q(n1133)
         );
  DFZX1 gate126 ( .D(n3128gat), .TD(n1133), .SEL(test_se), .CK(clk), .Q(n1134)
         );
  DFZX1 gate127 ( .D(n667), .TD(n1134), .SEL(test_se), .CK(clk), .Q(n2182gat)
         );
  DFZX1 gate128 ( .D(n2983gat), .TD(n2182gat), .SEL(test_se), .CK(clk), .Q(
        n1234), .QB(n711) );
  DFZX1 gate129 ( .D(n711), .TD(n1234), .SEL(test_se), .CK(clk), .Q(n1135), 
        .QB(n712) );
  DFZX1 gate130 ( .D(n712), .TD(n1135), .SEL(test_se), .CK(clk), .Q(n1233), 
        .QB(n713) );
  DFZX1 gate131 ( .D(n713), .TD(n1233), .SEL(test_se), .CK(clk), .Q(n1194) );
  DFZX1 gate132 ( .D(n1696gat), .TD(n1194), .SEL(test_se), .CK(clk), .Q(n1195), 
        .QB(n715) );
  DFZX1 gate133 ( .D(n2009gat), .TD(n1195), .SEL(test_se), .CK(clk), .Q(n1196), 
        .QB(n3106gat) );
  DFZX1 gate134 ( .D(n715), .TD(n1196), .SEL(test_se), .CK(clk), .Q(n1232), 
        .QB(n717) );
  DFZX1 gate135 ( .D(n1636gat), .TD(n1232), .SEL(test_se), .CK(clk), .Q(n1115)
         );
  DFZX1 gate136 ( .D(n232), .TD(n1115), .SEL(test_se), .CK(clk), .Q(n1114) );
  DFZX1 gate140 ( .D(n244), .TD(n1114), .SEL(test_se), .CK(clk), .Q(n1136), 
        .QB(n720) );
  DFZX1 gate141 ( .D(n720), .TD(n1136), .SEL(test_se), .CK(clk), .Q(n1087), 
        .QB(n721) );
  DFZX1 gate142 ( .D(n721), .TD(n1087), .SEL(test_se), .CK(clk), .Q(n1132) );
  DFZX1 gate143 ( .D(n2163gat), .TD(n1132), .SEL(test_se), .CK(clk), .Q(n1197)
         );
  DFZX1 gate144 ( .D(n185), .TD(n1197), .SEL(test_se), .CK(clk), .Q(n2040gat)
         );
  DFZX1 gate145 ( .D(n2015gat), .TD(n2040gat), .SEL(test_se), .CK(clk), .Q(
        n1231), .QB(n722) );
  DFZX1 gate146 ( .D(n722), .TD(n1231), .SEL(test_se), .CK(clk), .Q(n1230), 
        .QB(n723) );
  DFZX1 gate147 ( .D(n2017gat), .TD(n1230), .SEL(test_se), .CK(clk), .Q(n1229), 
        .QB(n724) );
  DFZX1 gate148 ( .D(n724), .TD(n1229), .SEL(test_se), .CK(clk), .Q(n1228), 
        .QB(n588) );
  DFZX1 gate149 ( .D(n700), .TD(n1228), .SEL(test_se), .CK(clk), .Q(n2266gat)
         );
  DFZX1 gate150 ( .D(n723), .TD(n2266gat), .SEL(test_se), .CK(clk), .Q(n1088), 
        .QB(n725) );
  DFZX1 gate151 ( .D(n725), .TD(n1088), .SEL(test_se), .CK(clk), .Q(n1227), 
        .QB(n726) );
  DFZX1 gate152 ( .D(n726), .TD(n1227), .SEL(test_se), .CK(clk), .Q(n1139), 
        .QB(n727) );
  DFZX1 gate153 ( .D(n727), .TD(n1139), .SEL(test_se), .CK(clk), .Q(n1226), 
        .QB(n728) );
  DFZX1 gate154 ( .D(n728), .TD(n1226), .SEL(test_se), .CK(clk), .Q(n1225), 
        .QB(n587) );
  DFZX1 gate155 ( .D(n704), .TD(n1225), .SEL(test_se), .CK(clk), .Q(n1975gat)
         );
  DFZX1 gate156 ( .D(n699), .TD(n1975gat), .SEL(test_se), .CK(clk), .Q(n1086)
         );
  DFZX1 gate157 ( .D(n682), .TD(n1086), .SEL(test_se), .CK(clk), .Q(n1198) );
  DFZX1 gate158 ( .D(n679), .TD(n1198), .SEL(test_se), .CK(clk), .Q(n1095), 
        .QB(n749) );
  DFZX1 gate159 ( .D(n683), .TD(n1095), .SEL(test_se), .CK(clk), .Q(n1199), 
        .QB(n750) );
  DFZX1 gate160 ( .D(n685), .TD(n1199), .SEL(test_se), .CK(clk), .Q(n1098) );
  DFZX1 gate161 ( .D(n684), .TD(n1098), .SEL(test_se), .CK(clk), .Q(n1094) );
  DFZX1 gate162 ( .D(n686), .TD(n1094), .SEL(test_se), .CK(clk), .Q(n1097) );
  DFZX1 gate163 ( .D(n687), .TD(n1097), .SEL(test_se), .CK(clk), .Q(n1096) );
  DFZX1 gate164 ( .D(n680), .TD(n1096), .SEL(test_se), .CK(clk), .Q(n1200) );
  DFZX1 gate165 ( .D(n681), .TD(n1200), .SEL(test_se), .CK(clk), .Q(n470gat)
         );
  DFZX1 gate166 ( .D(n678), .TD(n470gat), .SEL(test_se), .CK(clk), .Q(n148gat)
         );
  DFZX1 gate167 ( .D(n717), .TD(n148gat), .SEL(test_se), .CK(clk), .Q(n1224), 
        .QB(n729) );
  DFZX1 gate168 ( .D(n729), .TD(n1224), .SEL(test_se), .CK(clk), .Q(n1201) );
  DFZX1 gate169 ( .D(n1613gat), .TD(n1201), .SEL(test_se), .CK(clk), .Q(
        n1771gat) );
  DFZX1 gate170 ( .D(n1391gat), .TD(n1771gat), .SEL(test_se), .CK(clk), .Q(
        n1223), .QB(n576) );
  DFZX1 gate171 ( .D(n1927gat), .TD(n1223), .SEL(test_se), .CK(clk), .Q(n1222), 
        .QB(n1093) );
  DFZX1 gate172 ( .D(n707), .TD(n1222), .SEL(test_se), .CK(clk), .Q(n1221), 
        .QB(n1092) );
  DFZX1 gate173 ( .D(n705), .TD(n1221), .SEL(test_se), .CK(clk), .Q(n1220), 
        .QB(n568) );
  DFZX1 gate174 ( .D(n1567gat), .TD(n1220), .SEL(test_se), .CK(clk), .Q(n1202)
         );
  DFZX1 gate175 ( .D(n1564gat), .TD(n1202), .SEL(test_se), .CK(clk), .Q(n1219), 
        .QB(n569) );
  DFZX1 gate176 ( .D(n706), .TD(n1219), .SEL(test_se), .CK(clk), .Q(n1525gat)
         );
  DFZX1 gate177 ( .D(n1915gat), .TD(n1525gat), .SEL(test_se), .CK(clk), .Q(
        n1203), .QB(n760) );
  DFZX1 gate178 ( .D(n1800gat), .TD(n1203), .SEL(test_se), .CK(clk), .Q(n1204)
         );
  DFZX1 gate179 ( .D(n1593gat), .TD(n1204), .SEL(test_se), .CK(clk), .Q(
        test_so), .QB(n572) );
  INVCKX2 U521 ( .I(n1044), .O(n1057) );
  OAI12X1 U522 ( .B1(n671), .B2(n1216), .A1(n1044), .O(n1037) );
  TIE0X1 U523 ( .O(n1216) );
  TIE1X1 U524 ( .O(n3147gat) );
  AN3B2X1 U525 ( .I1(n761), .B1(n741), .B2(n762), .O(n706) );
  ND2X1 U526 ( .I1(n197), .I2(n763), .O(n674) );
  XOR2X1 U527 ( .I1(n2266gat), .I2(n764), .O(n763) );
  OR2B1XLP U528 ( .I1(n1134), .B1(n1193), .O(n764) );
  ND2X1 U529 ( .I1(n195), .I2(n765), .O(n673) );
  XOR2X1 U530 ( .I1(n1975gat), .I2(n766), .O(n765) );
  ND3X1 U531 ( .I1(n767), .I2(n741), .I3(n762), .O(n766) );
  ND2X1 U532 ( .I1(n768), .I2(n196), .O(n672) );
  XOR2X1 U533 ( .I1(n769), .I2(n1086), .O(n768) );
  ND3X1 U534 ( .I1(n770), .I2(n730), .I3(n771), .O(n769) );
  ND3X1 U535 ( .I1(n772), .I2(n773), .I3(n774), .O(n670) );
  AN4B1XLP U536 ( .I1(n1088), .I2(n1087), .I3(n775), .B1(n726), .O(n3146gat)
         );
  AOI112X1 U537 ( .C1(n1196), .C2(n776), .A1(n777), .B1(n723), .O(n775) );
  ND2X1 U538 ( .I1(n1132), .I2(n1136), .O(n777) );
  NR2X1 U539 ( .I1(n185), .I2(n776), .O(n3145gat) );
  AN2X1 U540 ( .I1(n1201), .I2(n778), .O(n776) );
  ND2X1 U541 ( .I1(n779), .I2(n780), .O(n3139gat) );
  OAI112X1 U542 ( .C1(n781), .C2(n758), .A1(n1196), .B1(n782), .O(n780) );
  OA112X1 U543 ( .C1(n676), .C2(n1141), .A1(n715), .B1(n783), .O(n782) );
  INVCKX1 U544 ( .I(n3098gat), .O(n783) );
  AN2X1 U545 ( .I1(n3097gat), .I2(n784), .O(n781) );
  MXL2XLP U546 ( .A(n785), .B(n786), .S(n787), .OB(n779) );
  OAI13X1 U547 ( .B1(n1525gat), .B2(n1113), .B3(n788), .A1(n789), .O(n786) );
  MXL2XLP U548 ( .A(n790), .B(n572), .S(n1204), .OB(n789) );
  AOI12X1 U549 ( .B1(n708), .B2(n791), .A1(n1114), .O(n790) );
  OAI22X1 U550 ( .A1(n1114), .A2(n760), .B1(n1115), .B2(n792), .O(n785) );
  INVCKX1 U551 ( .I(n793), .O(n792) );
  OAI33X1 U552 ( .A1(n794), .A2(n1202), .A3(n795), .B1(n796), .B2(n1203), .B3(
        n708), .O(n793) );
  ND2X1 U553 ( .I1(n797), .I2(n798), .O(n3016gat) );
  AN4B1XLP U554 ( .I1(n2522gat), .I2(n2526gat), .I3(n2464gat), .B1(n1090), .O(
        n798) );
  AN4B1XLP U555 ( .I1(n2476gat), .I2(n2468gat), .I3(n1089), .B1(n3090gat), .O(
        n797) );
  AOI112X1 U556 ( .C1(n2182gat), .C2(n799), .A1(n800), .B1(n801), .O(n2983gat)
         );
  ND2X1 U557 ( .I1(n1091), .I2(n802), .O(n799) );
  MXL2XLP U558 ( .A(n803), .B(n804), .S(n787), .OB(n3142gat) );
  AOI23X1 U559 ( .B1(n186), .B2(n708), .B3(n1092), .A1(n1093), .A2(n805), .O(
        n804) );
  OAI112X1 U560 ( .C1(n788), .C2(n576), .A1(n791), .B1(n796), .O(n805) );
  AOI22X1 U561 ( .A1(n806), .A2(n569), .B1(n1202), .B2(n568), .O(n803) );
  OAI12X1 U562 ( .B1(n1202), .B2(n795), .A1(n796), .O(n806) );
  AN2X1 U563 ( .I1(n791), .I2(n788), .O(n795) );
  OAI22X1 U564 ( .A1(n807), .A2(n808), .B1(n809), .B2(n810), .O(n3133gat) );
  OA222X1 U565 ( .A1(n811), .A2(n1166), .B1(n812), .B2(n1155), .C1(n813), .C2(
        n1171), .O(n810) );
  OAI22X1 U566 ( .A1(n814), .A2(n808), .B1(n809), .B2(n815), .O(n3130gat) );
  AOI222X1 U567 ( .A1(n816), .A2(n732), .B1(n817), .B2(n752), .C1(n818), .C2(
        n678), .O(n815) );
  OAI12X1 U568 ( .B1(n819), .B2(n820), .A1(n821), .O(n2952gat) );
  OAI22X1 U569 ( .A1(n822), .A2(n808), .B1(n809), .B2(n823), .O(n3129gat) );
  OA222X1 U570 ( .A1(n811), .A2(n1101), .B1(n812), .B2(n824), .C1(n813), .C2(
        n1099), .O(n823) );
  INVCKX1 U571 ( .I(n3116gat), .O(n824) );
  OAI22X1 U572 ( .A1(n825), .A2(n808), .B1(n809), .B2(n826), .O(n3136gat) );
  OA222X1 U573 ( .A1(n811), .A2(n1145), .B1(n812), .B2(n1158), .C1(n813), .C2(
        n1207), .O(n826) );
  OAI22X1 U574 ( .A1(n827), .A2(n808), .B1(n809), .B2(n828), .O(n3137gat) );
  OA222X1 U575 ( .A1(n811), .A2(n1144), .B1(n812), .B2(n1154), .C1(n813), .C2(
        n1100), .O(n828) );
  OAI22X1 U576 ( .A1(n829), .A2(n808), .B1(n809), .B2(n830), .O(n3132gat) );
  OA222X1 U577 ( .A1(n811), .A2(n1105), .B1(n812), .B2(n1156), .C1(n813), .C2(
        n1104), .O(n830) );
  OAI22X1 U578 ( .A1(n831), .A2(n808), .B1(n809), .B2(n832), .O(n3134gat) );
  OA222X1 U579 ( .A1(n811), .A2(n1160), .B1(n812), .B2(n1153), .C1(n813), .C2(
        n1206), .O(n832) );
  OAI22X1 U580 ( .A1(n833), .A2(n808), .B1(n809), .B2(n834), .O(n3131gat) );
  OA222X1 U581 ( .A1(n811), .A2(n1165), .B1(n812), .B2(n1157), .C1(n813), .C2(
        n1170), .O(n834) );
  OAI22X1 U582 ( .A1(n835), .A2(n808), .B1(n809), .B2(n836), .O(n3135gat) );
  OA222X1 U583 ( .A1(n811), .A2(n1146), .B1(n812), .B2(n1152), .C1(n813), .C2(
        n1205), .O(n836) );
  OA12X1 U584 ( .B1(n837), .B2(n838), .A1(n839), .O(n809) );
  MXL2XLP U585 ( .A(n840), .B(n841), .S(n3088gat), .OB(n808) );
  AN4B1XLP U586 ( .I1(n842), .I2(n843), .I3(n844), .B1(n3085gat), .O(n841) );
  INVCKX1 U587 ( .I(n838), .O(n840) );
  OAI12X1 U588 ( .B1(n845), .B2(n846), .A1(n842), .O(n838) );
  OAI222X1 U589 ( .A1(n847), .A2(n848), .B1(n849), .B2(n850), .C1(n851), .C2(
        n852), .O(n2929gat) );
  XNR2X1 U590 ( .I1(n1098), .I2(n853), .O(n850) );
  MXL2XLP U591 ( .A(n854), .B(n855), .S(n856), .OB(n2926gat) );
  XOR2X1 U592 ( .I1(n470gat), .I2(n857), .O(n855) );
  NR2X1 U593 ( .I1(n858), .I2(n859), .O(n857) );
  AOI12X1 U594 ( .B1(n1200), .B2(n749), .A1(n1198), .O(n858) );
  OAI222X1 U595 ( .A1(n847), .A2(n854), .B1(n849), .B2(n860), .C1(n851), .C2(
        n861), .O(n2925gat) );
  XOR2X1 U596 ( .I1(n1094), .I2(n862), .O(n860) );
  NR2X1 U597 ( .I1(n863), .I2(n853), .O(n862) );
  AOI12X1 U598 ( .B1(n1097), .B2(n750), .A1(n1098), .O(n863) );
  MXL2XLP U599 ( .A(n864), .B(n865), .S(n856), .OB(n2924gat) );
  XNR2X1 U600 ( .I1(n1200), .I2(n866), .O(n865) );
  MXL2XLP U601 ( .A(n867), .B(n868), .S(n856), .OB(n2923gat) );
  XOR2X1 U602 ( .I1(n148gat), .I2(n869), .O(n868) );
  NR2X1 U603 ( .I1(n1200), .I2(n866), .O(n869) );
  ND2X1 U604 ( .I1(n870), .I2(n749), .O(n866) );
  OAI22X1 U605 ( .A1(n851), .A2(n871), .B1(n820), .B2(n847), .O(n2920gat) );
  OAI12X1 U606 ( .B1(n819), .B2(n864), .A1(n821), .O(n2919gat) );
  OAI12X1 U607 ( .B1(n819), .B2(n867), .A1(n821), .O(n2918gat) );
  MXL2XLP U608 ( .A(n820), .B(n872), .S(n856), .OB(n2917gat) );
  XOR2X1 U609 ( .I1(n1095), .I2(n870), .O(n872) );
  NR2X1 U610 ( .I1(n859), .I2(n1198), .O(n870) );
  OAI222X1 U611 ( .A1(n847), .A2(n873), .B1(n849), .B2(n874), .C1(n851), .C2(
        n875), .O(n2916gat) );
  XNR2X1 U612 ( .I1(n1097), .I2(n876), .O(n874) );
  OR2B1XLP U613 ( .I1(n2927gat), .B1(n821), .O(n2915gat) );
  OAI22X1 U614 ( .A1(n877), .A2(n878), .B1(n879), .B2(n864), .O(n2927gat) );
  OAI22X1 U615 ( .A1(n851), .A2(n880), .B1(n847), .B2(n867), .O(n2913gat) );
  OAI12X1 U616 ( .B1(n819), .B2(n873), .A1(n821), .O(n2912gat) );
  OAI12X1 U617 ( .B1(n819), .B2(n881), .A1(n821), .O(n2911gat) );
  OAI12X1 U618 ( .B1(n819), .B2(n882), .A1(n821), .O(n2910gat) );
  OAI12X1 U619 ( .B1(n819), .B2(n883), .A1(n821), .O(n2909gat) );
  OAI12X1 U620 ( .B1(n819), .B2(n854), .A1(n821), .O(n2908gat) );
  OAI12X1 U621 ( .B1(n819), .B2(n848), .A1(n821), .O(n2907gat) );
  AOI33X1 U622 ( .A1(n884), .A2(n3086gat), .A3(n885), .B1(n886), .B2(n837), 
        .B3(n887), .O(n819) );
  OAI22X1 U623 ( .A1(n851), .A2(n878), .B1(n847), .B2(n864), .O(n2905gat) );
  INVCKX1 U624 ( .I(n3066gat), .O(n864) );
  INVCKX1 U625 ( .I(n3075gat), .O(n878) );
  OR2B1XLP U626 ( .I1(n2922gat), .B1(n821), .O(n2904gat) );
  OAI22X1 U627 ( .A1(n877), .A2(n861), .B1(n879), .B2(n854), .O(n2922gat) );
  INVCKX1 U628 ( .I(n3073gat), .O(n854) );
  INVCKX1 U629 ( .I(n3082gat), .O(n861) );
  OR2B1XLP U630 ( .I1(n2928gat), .B1(n821), .O(n2903gat) );
  OAI22X1 U631 ( .A1(n877), .A2(n871), .B1(n879), .B2(n820), .O(n2928gat) );
  INVCKX1 U632 ( .I(n3067gat), .O(n820) );
  INVCKX1 U633 ( .I(n3076gat), .O(n871) );
  OR2B1XLP U634 ( .I1(n2896gat), .B1(n821), .O(n2901gat) );
  OAI222X1 U635 ( .A1(n847), .A2(n882), .B1(n849), .B2(n888), .C1(n851), .C2(
        n889), .O(n2900gat) );
  XOR2X1 U636 ( .I1(n1199), .I2(n890), .O(n888) );
  OAI222X1 U637 ( .A1(n847), .A2(n883), .B1(n849), .B2(n891), .C1(n851), .C2(
        n892), .O(n2899gat) );
  XOR2X1 U638 ( .I1(n1096), .I2(n893), .O(n891) );
  NR2X1 U639 ( .I1(n1097), .I2(n876), .O(n893) );
  ND2X1 U640 ( .I1(n890), .I2(n750), .O(n876) );
  NR2X1 U641 ( .I1(n853), .I2(n1098), .O(n890) );
  ND2X1 U642 ( .I1(n851), .I2(n847), .O(n849) );
  OAI22X1 U643 ( .A1(n851), .A2(n894), .B1(n847), .B2(n881), .O(n2898gat) );
  OR4B2XLP U644 ( .I1(n3088gat), .I2(n3086gat), .B1(n3093gat), .B2(n895), .O(
        n847) );
  OAI22X1 U645 ( .A1(n877), .A2(n889), .B1(n879), .B2(n882), .O(n2896gat) );
  INVCKX1 U646 ( .I(n3071gat), .O(n882) );
  INVCKX1 U647 ( .I(n3080gat), .O(n889) );
  MXL2XLP U648 ( .A(n881), .B(n896), .S(n856), .OB(n2892gat) );
  AN2X1 U649 ( .I1(n851), .I2(n897), .O(n856) );
  OR4B2XLP U650 ( .I1(n3086gat), .I2(n898), .B1(n885), .B2(n899), .O(n897) );
  ND3X1 U651 ( .I1(n3088gat), .I2(n900), .I3(n886), .O(n851) );
  XNR2X1 U652 ( .I1(n1198), .I2(n859), .O(n896) );
  OR2B1XLP U653 ( .I1(n2914gat), .B1(n821), .O(n2891gat) );
  OAI22X1 U654 ( .A1(n877), .A2(n880), .B1(n879), .B2(n867), .O(n2914gat) );
  INVCKX1 U655 ( .I(n3065gat), .O(n867) );
  INVCKX1 U656 ( .I(n3074gat), .O(n880) );
  OR2B1XLP U657 ( .I1(n2897gat), .B1(n821), .O(n2890gat) );
  OAI22X1 U658 ( .A1(n877), .A2(n852), .B1(n879), .B2(n848), .O(n2897gat) );
  INVCKX1 U659 ( .I(n3072gat), .O(n848) );
  INVCKX1 U660 ( .I(n3081gat), .O(n852) );
  OR2B1XLP U661 ( .I1(n2894gat), .B1(n821), .O(n2888gat) );
  OAI22X1 U662 ( .A1(n877), .A2(n894), .B1(n879), .B2(n881), .O(n2894gat) );
  INVCKX1 U663 ( .I(n3068gat), .O(n881) );
  INVCKX1 U664 ( .I(n3077gat), .O(n894) );
  OR2B1XLP U665 ( .I1(n2921gat), .B1(n821), .O(n2887gat) );
  OAI22X1 U666 ( .A1(n877), .A2(n875), .B1(n879), .B2(n873), .O(n2921gat) );
  INVCKX1 U667 ( .I(n3070gat), .O(n873) );
  INVCKX1 U668 ( .I(n3079gat), .O(n875) );
  OR2B1XLP U669 ( .I1(n2895gat), .B1(n821), .O(n2886gat) );
  OR4B2XLP U670 ( .I1(n1179), .I2(n788), .B1(n695), .B2(n901), .O(n821) );
  AOI112X1 U671 ( .C1(n902), .C2(n690), .A1(n903), .B1(n794), .O(n901) );
  NR3X1 U672 ( .I1(n904), .I2(n905), .I3(n691), .O(n794) );
  MXL2XLP U673 ( .A(n906), .B(n907), .S(n1183), .OB(n903) );
  AN4B2X1 U674 ( .I1(n1151), .I2(n1214), .B1(n1180), .B2(n1215), .O(n906) );
  INVCKX1 U675 ( .I(n186), .O(n788) );
  OAI22X1 U676 ( .A1(n877), .A2(n892), .B1(n879), .B2(n883), .O(n2895gat) );
  INVCKX1 U677 ( .I(n3069gat), .O(n883) );
  INVCKX1 U678 ( .I(n3078gat), .O(n892) );
  OAI112X1 U679 ( .C1(n908), .C2(n909), .A1(n910), .B1(n911), .O(n3104gat) );
  OR4B2XLP U680 ( .I1(n3088gat), .I2(n900), .B1(n912), .B2(n3094gat), .O(n910)
         );
  ND2X1 U681 ( .I1(n913), .I2(n914), .O(n3105gat) );
  AOI33X1 U682 ( .A1(n885), .A2(n915), .A3(n884), .B1(n900), .B2(n837), .B3(
        n886), .O(n913) );
  ND2X1 U683 ( .I1(n916), .I2(n2613gat), .O(n3143gat) );
  ND2X1 U684 ( .I1(n1157), .I2(n917), .O(n3109gat) );
  ND2X1 U685 ( .I1(n1184), .I2(n918), .O(n3108gat) );
  OAI12X1 U686 ( .B1(n822), .B2(n839), .A1(n231), .O(n3125gat) );
  INVCKX1 U687 ( .I(n919), .O(n822) );
  OAI122X1 U688 ( .B1(n1164), .B2(n920), .C1(n1213), .C2(n811), .A1(n921), .O(
        n919) );
  AOI122X1 U689 ( .B1(n818), .B2(n684), .C1(n817), .C2(n922), .A1(n923), .O(
        n921) );
  AOI112X1 U690 ( .C1(n737), .C2(n924), .A1(n925), .B1(n926), .O(n923) );
  INVCKX1 U691 ( .I(n927), .O(n924) );
  OAI12X1 U692 ( .B1(n827), .B2(n839), .A1(n2971gat), .O(n3124gat) );
  XNR2X1 U693 ( .I1(n1197gat), .I2(n3116gat), .O(n2971gat) );
  OA112X1 U694 ( .C1(n1112), .C2(n813), .A1(n928), .B1(n929), .O(n827) );
  OA22X1 U695 ( .A1(n920), .A2(n1162), .B1(n811), .B2(n1111), .O(n929) );
  AOI23X1 U696 ( .B1(n930), .B2(n737), .B3(n931), .A1(n817), .A2(n759), .O(
        n928) );
  INVCKX1 U697 ( .I(n812), .O(n817) );
  OAI12X1 U698 ( .B1(n825), .B2(n839), .A1(n3010gat), .O(n3123gat) );
  XOR2X1 U699 ( .I1(n667gat), .I2(n932), .O(n3010gat) );
  INVCKX1 U700 ( .I(n933), .O(n825) );
  OAI122X1 U701 ( .B1(n1163), .B2(n920), .C1(n1212), .C2(n811), .A1(n934), .O(
        n933) );
  OA22X1 U702 ( .A1(n812), .A2(n1121), .B1(n813), .B2(n1209), .O(n934) );
  OAI12X1 U703 ( .B1(n835), .B2(n839), .A1(n504gat), .O(n3122gat) );
  XOR3X1 U704 ( .I1(n935), .I2(n936), .I3(n1104), .O(n504gat) );
  XOR4XLP U705 ( .I1(n1206), .I2(n1207), .I3(n1171), .I4(n1205), .O(n936) );
  XOR4XLP U706 ( .I1(n1106), .I2(n1170), .I3(n1099), .I4(n1100), .O(n935) );
  INVCKX1 U707 ( .I(n937), .O(n835) );
  OAI122X1 U708 ( .B1(n1161), .B2(n920), .C1(n1169), .C2(n811), .A1(n938), .O(
        n937) );
  OA22X1 U709 ( .A1(n812), .A2(n1116), .B1(n813), .B2(n1174), .O(n938) );
  OAI12X1 U710 ( .B1(n831), .B2(n839), .A1(n567gat), .O(n3121gat) );
  XOR3X1 U711 ( .I1(n939), .I2(n940), .I3(n1107), .O(n567gat) );
  XOR4XLP U712 ( .I1(n1209), .I2(n1210), .I3(n1174), .I4(n1208), .O(n940) );
  XOR4XLP U713 ( .I1(n1172), .I2(n1173), .I3(n1110), .I4(n1112), .O(n939) );
  AOI122X1 U714 ( .B1(n731), .B2(n941), .C1(n739), .C2(n816), .A1(n942), .O(
        n831) );
  OAI22X1 U715 ( .A1(n812), .A2(n1117), .B1(n813), .B2(n1110), .O(n942) );
  OAI12X1 U716 ( .B1(n807), .B2(n839), .A1(n55gat), .O(n3120gat) );
  XNR2X1 U717 ( .I1(n943), .I2(n944), .O(n55gat) );
  XOR4XLP U718 ( .I1(n1145), .I2(n1165), .I3(n1166), .I4(n945), .O(n944) );
  OAI12X1 U719 ( .B1(n1160), .B2(n751), .A1(n946), .O(n945) );
  XOR4XLP U720 ( .I1(n1101), .I2(n1105), .I3(n1144), .I4(n732), .O(n943) );
  INVCKX1 U721 ( .I(n947), .O(n807) );
  OAI122X1 U722 ( .B1(n1122), .B2(n920), .C1(n1168), .C2(n811), .A1(n948), .O(
        n947) );
  OA22X1 U723 ( .A1(n812), .A2(n1119), .B1(n813), .B2(n1173), .O(n948) );
  OAI12X1 U724 ( .B1(n829), .B2(n839), .A1(n933gat), .O(n3119gat) );
  XOR3X1 U725 ( .I1(n949), .I2(n950), .I3(n1108), .O(n933gat) );
  XOR4XLP U726 ( .I1(n1212), .I2(n1213), .I3(n1169), .I4(n1211), .O(n950) );
  XOR4XLP U727 ( .I1(n1167), .I2(n1168), .I3(n1109), .I4(n1111), .O(n949) );
  INVCKX1 U728 ( .I(n951), .O(n829) );
  OAI122X1 U729 ( .B1(n1123), .B2(n920), .C1(n1108), .C2(n811), .A1(n952), .O(
        n951) );
  MAOI1X1 U730 ( .A1(n818), .A2(n738), .B1(n812), .B2(n1120), .O(n952) );
  INVCKX1 U731 ( .I(n813), .O(n818) );
  ND2X1 U732 ( .I1(n2579gat), .I2(n916), .O(n3144gat) );
  INVCKX1 U733 ( .I(n953), .O(n916) );
  OAI122X1 U734 ( .B1(n954), .B2(n791), .C1(n1102), .C2(n955), .A1(n956), .O(
        n953) );
  AOI33X1 U735 ( .A1(n3149gat), .A2(n708), .A3(n957), .B1(n737), .B2(n717), 
        .B3(n1196), .O(n956) );
  MXL2XLP U736 ( .A(n1115), .B(n1114), .S(n787), .OB(n957) );
  AOI22X1 U737 ( .A1(n958), .A2(n959), .B1(n960), .B2(n961), .O(n955) );
  OAI122X1 U738 ( .B1(n962), .B2(n904), .C1(n963), .C2(n964), .A1(n965), .O(
        n961) );
  AOI22X1 U739 ( .A1(n966), .A2(n967), .B1(n968), .B2(n969), .O(n965) );
  OAI22X1 U740 ( .A1(n1112), .A2(n970), .B1(n1111), .B2(n971), .O(n969) );
  MXL2XLP U741 ( .A(n1212), .B(n1209), .S(n796), .OB(n966) );
  AOI122X1 U742 ( .B1(n972), .B2(n756), .C1(n973), .C2(n679), .A1(n974), .O(
        n963) );
  OAI22X1 U743 ( .A1(n1171), .A2(n970), .B1(n1166), .B2(n971), .O(n974) );
  AOI122X1 U744 ( .B1(n972), .B2(n732), .C1(n973), .C2(n678), .A1(n975), .O(
        n962) );
  OAI22X1 U745 ( .A1(n1170), .A2(n970), .B1(n1165), .B2(n971), .O(n975) );
  OAI122X1 U746 ( .B1(n976), .B2(n904), .C1(n977), .C2(n964), .A1(n978), .O(
        n959) );
  AOI222X1 U747 ( .A1(n979), .A2(n980), .B1(n967), .B2(n981), .C1(n902), .C2(
        n982), .O(n978) );
  ND2X1 U748 ( .I1(n1103), .I2(n983), .O(n981) );
  OAI122X1 U749 ( .B1(n1169), .B2(n971), .C1(n1174), .C2(n970), .A1(n984), .O(
        n980) );
  AOI22X1 U750 ( .A1(n972), .A2(n739), .B1(n973), .B2(n687), .O(n984) );
  INVCKX1 U751 ( .I(n985), .O(n979) );
  AOI122X1 U752 ( .B1(n972), .B2(n755), .C1(n973), .C2(n738), .A1(n986), .O(
        n977) );
  OAI22X1 U753 ( .A1(n1173), .A2(n970), .B1(n1168), .B2(n971), .O(n986) );
  AOI122X1 U754 ( .B1(n972), .B2(n740), .C1(n973), .C2(n754), .A1(n987), .O(
        n976) );
  OAI22X1 U755 ( .A1(n1172), .A2(n970), .B1(n1167), .B2(n971), .O(n987) );
  ND2X1 U756 ( .I1(n691), .I2(n3149gat), .O(n971) );
  ND2X1 U757 ( .I1(n796), .I2(n691), .O(n970) );
  NR2X1 U758 ( .I1(n691), .I2(n3149gat), .O(n973) );
  NR2X1 U759 ( .I1(n691), .I2(n796), .O(n972) );
  INVCKX1 U760 ( .I(n3149gat), .O(n796) );
  INVCKX1 U761 ( .I(n988), .O(n958) );
  AOI23X1 U762 ( .B1(n989), .B2(n990), .B3(n967), .A1(n991), .A2(n992), .O(
        n954) );
  OAI12X1 U763 ( .B1(n1185), .B2(n993), .A1(n994), .O(n992) );
  MXL2XLP U764 ( .A(n995), .B(n996), .S(n1178), .OB(n994) );
  OAI222X1 U765 ( .A1(n1120), .A2(n904), .B1(n1121), .B2(n985), .C1(n1117), 
        .C2(n964), .O(n996) );
  OAI122X1 U766 ( .B1(n1116), .B2(n964), .C1(n1124), .C2(n997), .A1(n998), .O(
        n995) );
  OA22X1 U767 ( .A1(n985), .A2(n1118), .B1(n904), .B2(n1119), .O(n998) );
  ND2X1 U768 ( .I1(n1175), .I2(n689), .O(n904) );
  ND2X1 U769 ( .I1(n689), .I2(n688), .O(n985) );
  ND2X1 U770 ( .I1(n1176), .I2(n688), .O(n964) );
  INVCKX1 U771 ( .I(n993), .O(n967) );
  XOR2X1 U772 ( .I1(n1162), .I2(n932), .O(n990) );
  INVCKX1 U773 ( .I(n922), .O(n932) );
  XNR2X1 U774 ( .I1(n999), .I2(n1000), .O(n922) );
  XOR4XLP U775 ( .I1(n1118), .I2(n1119), .I3(n1116), .I4(n1117), .O(n1000) );
  XOR4XLP U776 ( .I1(n1120), .I2(n1121), .I3(n1185), .I4(n1124), .O(n999) );
  OAI12X1 U777 ( .B1(n833), .B2(n839), .A1(n43gat), .O(n3118gat) );
  XOR4XLP U778 ( .I1(n1159), .I2(n1161), .I3(n1001), .I4(n1002), .O(n43gat) );
  XOR4XLP U779 ( .I1(n1125), .I2(n1143), .I3(n1122), .I4(n1123), .O(n1002) );
  OAI12X1 U780 ( .B1(n1003), .B2(n753), .A1(n1004), .O(n1001) );
  MXL2XLP U781 ( .A(n1005), .B(n1006), .S(n1162), .OB(n1004) );
  NR2X1 U782 ( .I1(n1163), .I2(n1164), .O(n1006) );
  XOR2X1 U783 ( .I1(n1163), .I2(n1164), .O(n1005) );
  INVCKX1 U784 ( .I(n1007), .O(n833) );
  OAI122X1 U785 ( .B1(n1125), .B2(n920), .C1(n1167), .C2(n811), .A1(n1008), 
        .O(n1007) );
  OA22X1 U786 ( .A1(n812), .A2(n1124), .B1(n813), .B2(n1172), .O(n1008) );
  OAI12X1 U787 ( .B1(n814), .B2(n839), .A1(n748gat), .O(n3117gat) );
  XOR4XLP U788 ( .I1(n3086gat), .I2(n1009), .I3(n898), .I4(n1010), .O(n748gat)
         );
  XOR2X1 U789 ( .I1(n3089gat), .I2(n3088gat), .O(n1010) );
  MXL2XLP U790 ( .A(n1011), .B(n1012), .S(n3085gat), .OB(n1009) );
  AOI12X1 U791 ( .B1(n3083gat), .B2(n3084gat), .A1(n842), .O(n1012) );
  XNR2X1 U792 ( .I1(n3083gat), .I2(n3084gat), .O(n1011) );
  OAI112X1 U793 ( .C1(n843), .C2(n844), .A1(n1013), .B1(n842), .O(n839) );
  AOI122X1 U794 ( .B1(n757), .B2(n941), .C1(n740), .C2(n816), .A1(n1014), .O(
        n814) );
  OAI22X1 U795 ( .A1(n812), .A2(n1185), .B1(n813), .B2(n1208), .O(n1014) );
  ND2X1 U796 ( .I1(n927), .I2(n925), .O(n813) );
  ND2X1 U797 ( .I1(n926), .I2(n930), .O(n812) );
  INVCKX1 U798 ( .I(n925), .O(n930) );
  INVCKX1 U799 ( .I(n811), .O(n816) );
  ND2X1 U800 ( .I1(n931), .I2(n925), .O(n811) );
  INVCKX1 U801 ( .I(n920), .O(n941) );
  ND2X1 U802 ( .I1(n926), .I2(n925), .O(n920) );
  OAI22X1 U803 ( .A1(n837), .A2(n877), .B1(n898), .B2(n879), .O(n925) );
  NR2X1 U804 ( .I1(n927), .I2(n931), .O(n926) );
  NR2X1 U805 ( .I1(n844), .I2(n845), .O(n931) );
  NR2X1 U806 ( .I1(n879), .I2(n1013), .O(n845) );
  NR2X1 U807 ( .I1(n846), .I2(n843), .O(n927) );
  ND2X1 U808 ( .I1(n1015), .I2(n1155), .O(n3111gat) );
  ND2X1 U809 ( .I1(n1156), .I2(n1016), .O(n3110gat) );
  OAI112X1 U810 ( .C1(n900), .C2(n1017), .A1(n909), .B1(n1018), .O(n3151gat)
         );
  ND3X1 U811 ( .I1(n3086gat), .I2(n1013), .I3(n884), .O(n909) );
  AN2X1 U812 ( .I1(n899), .I2(n898), .O(n884) );
  AN4B1XLP U813 ( .I1(n842), .I2(n1196), .I3(n3088gat), .B1(n879), .O(n899) );
  ND2X1 U814 ( .I1(n912), .I2(n837), .O(n1017) );
  INVCKX1 U815 ( .I(n3088gat), .O(n837) );
  ND2X1 U816 ( .I1(n1152), .I2(n1019), .O(n3113gat) );
  ND2X1 U817 ( .I1(n1020), .I2(n1158), .O(n3114gat) );
  OAI12X1 U818 ( .B1(n1125), .B2(n1197), .A1(n1021), .O(n3150gat) );
  XOR4XLP U819 ( .I1(n1214), .I2(n1215), .I3(n704), .I4(n1022), .O(n2613gat)
         );
  XOR3X1 U820 ( .I1(n1151), .I2(n1180), .I3(n1181), .O(n1022) );
  XOR4XLP U821 ( .I1(n1178), .I2(n1023), .I3(n689), .I4(n1129), .O(n2579gat)
         );
  MXL2XLP U822 ( .A(n1024), .B(n1025), .S(n1175), .OB(n1023) );
  OR2X1 U823 ( .I1(n991), .I2(n960), .O(n1025) );
  AN2B1XLP U824 ( .I1(n1179), .B1(n1177), .O(n960) );
  ND2X1 U825 ( .I1(n905), .I2(n988), .O(n1024) );
  ND2X1 U826 ( .I1(n1179), .I2(n1177), .O(n988) );
  NR2X1 U827 ( .I1(n911), .I2(n1026), .O(n2556gat) );
  AOI12X1 U828 ( .B1(n767), .B2(n735), .A1(n705), .O(n911) );
  MXL2XLP U829 ( .A(n1027), .B(n1028), .S(n3088gat), .OB(n244) );
  ND2X1 U830 ( .I1(n886), .I2(n887), .O(n1028) );
  INVCKX1 U831 ( .I(n900), .O(n887) );
  ND2X1 U832 ( .I1(n1029), .I2(n843), .O(n900) );
  NR2X1 U833 ( .I1(n877), .I2(n898), .O(n843) );
  AN2B1XLP U834 ( .I1(n3094gat), .B1(n912), .O(n886) );
  ND2X1 U835 ( .I1(n1029), .I2(n844), .O(n912) );
  NR2X1 U836 ( .I1(n877), .I2(n915), .O(n844) );
  INVCKX1 U837 ( .I(n3095gat), .O(n877) );
  AN3X1 U838 ( .I1(n1196), .I2(n1013), .I3(n842), .O(n1029) );
  ND2X1 U839 ( .I1(n846), .I2(n895), .O(n1027) );
  AN4B1XLP U840 ( .I1(n885), .I2(n1196), .I3(n842), .B1(n898), .O(n895) );
  INVCKX1 U841 ( .I(n3087gat), .O(n898) );
  NR2X1 U842 ( .I1(n3083gat), .I2(n3084gat), .O(n842) );
  NR2X1 U843 ( .I1(n1013), .I2(n908), .O(n885) );
  NR2X1 U844 ( .I1(n3091gat), .I2(n3092gat), .O(n908) );
  INVCKX1 U845 ( .I(n3085gat), .O(n1013) );
  NR2X1 U846 ( .I1(n879), .I2(n915), .O(n846) );
  INVCKX1 U847 ( .I(n3086gat), .O(n915) );
  INVCKX1 U848 ( .I(n3093gat), .O(n879) );
  NR2X1 U849 ( .I1(n1026), .I2(n914), .O(n2436gat) );
  XOR2X1 U850 ( .I1(n1147), .I2(n1030), .O(n914) );
  NR2X1 U851 ( .I1(n1031), .I2(n1016), .O(n2396gat) );
  XOR2X1 U852 ( .I1(n1187), .I2(n1032), .O(n1016) );
  NR2X1 U853 ( .I1(n1026), .I2(n1021), .O(n2387gat) );
  AO112X1 U854 ( .C1(n1186), .C2(n1148), .A1(n1033), .B1(n1030), .O(n1021) );
  NR2X1 U855 ( .I1(n1018), .I2(n1026), .O(n2330gat) );
  INVCKX1 U856 ( .I(n1034), .O(n232) );
  XOR4XLP U857 ( .I1(n1126), .I2(n1127), .I3(n3126gat), .I4(n1128), .O(n231)
         );
  NR2X1 U858 ( .I1(n1015), .I2(n1031), .O(n2198gat) );
  NR2X1 U859 ( .I1(n1031), .I2(n918), .O(n2197gat) );
  XOR2X1 U860 ( .I1(n770), .I2(n742), .O(n918) );
  NR2X1 U861 ( .I1(n1031), .I2(n917), .O(n2196gat) );
  ND2X1 U862 ( .I1(n770), .I2(n1035), .O(n917) );
  AO12X1 U863 ( .B1(n743), .B2(n1032), .A1(n733), .O(n1035) );
  ND3X1 U864 ( .I1(n733), .I2(n743), .I3(n1032), .O(n770) );
  NR2X1 U865 ( .I1(n1020), .I2(n1036), .O(n2194gat) );
  AN2X1 U866 ( .I1(n1134), .I2(n1193), .O(n1020) );
  AN4B2X1 U867 ( .I1(n1194), .I2(n1037), .B1(n1038), .B2(n1132), .O(n2163gat)
         );
  NR2X1 U868 ( .I1(n1036), .I2(n1019), .O(n2057gat) );
  OR2B1XLP U869 ( .I1(n802), .B1(n1039), .O(n1019) );
  OAI12X1 U870 ( .B1(n1193), .B2(n1134), .A1(n1133), .O(n1039) );
  NR3X1 U871 ( .I1(n1134), .I2(n1133), .I3(n1193), .O(n802) );
  NR3X1 U872 ( .I1(n2040gat), .I2(n1135), .I3(n1195), .O(n2015gat) );
  OA112X1 U873 ( .C1(n715), .C2(n1194), .A1(n2017gat), .B1(n1037), .O(n2009gat) );
  NR2X1 U874 ( .I1(n784), .I2(n1038), .O(n2017gat) );
  INVCKX1 U875 ( .I(n1031), .O(n196) );
  ND2X1 U876 ( .I1(n197), .I2(n800), .O(n1031) );
  MXL2XLP U877 ( .A(n1040), .B(n1041), .S(n2989gat), .OB(n800) );
  AN4B1XLP U878 ( .I1(n733), .I2(n742), .I3(n730), .B1(n1042), .O(n1040) );
  ND2X1 U879 ( .I1(n1187), .I2(n1188), .O(n1042) );
  INVCKX1 U880 ( .I(n1026), .O(n195) );
  ND2X1 U881 ( .I1(n801), .I2(n197), .O(n1026) );
  INVCKX1 U882 ( .I(n1036), .O(n197) );
  OAI112X1 U883 ( .C1(n784), .C2(n588), .A1(n1037), .B1(n1043), .O(n1036) );
  AN2B1XLP U884 ( .I1(n1136), .B1(n723), .O(n1043) );
  OR4B2XLP U885 ( .I1(n608), .I2(n657), .B1(n1045), .B2(n1138), .O(n671) );
  NR2X1 U886 ( .I1(n1137), .I2(n606), .O(n1045) );
  AN2X1 U887 ( .I1(n1182), .I2(n2021gat), .O(n784) );
  AN2X1 U888 ( .I1(n1046), .I2(n1047), .O(n801) );
  MXL2XLP U889 ( .A(n1048), .B(n1049), .S(n1192), .OB(n1047) );
  NR2X1 U890 ( .I1(n787), .I2(n1050), .O(n1049) );
  INVCKX1 U891 ( .I(n2989gat), .O(n787) );
  MXL2XLP U892 ( .A(n1051), .B(n1052), .S(n1053), .OB(n1046) );
  NR2X1 U893 ( .I1(n1131), .I2(n1130), .O(n1053) );
  AN2B1XLP U894 ( .I1(n707), .B1(n2989gat), .O(n1052) );
  NR3X1 U895 ( .I1(n1054), .I2(n1186), .I3(n734), .O(n707) );
  NR2X1 U896 ( .I1(n2989gat), .I2(n1055), .O(n1051) );
  NR2X1 U897 ( .I1(n1038), .I2(n1055), .O(n1927gat) );
  NR2X1 U898 ( .I1(n1050), .I2(n1056), .O(n1915gat) );
  INVCKX1 U899 ( .I(n705), .O(n1050) );
  NR2X1 U900 ( .I1(n767), .I2(n735), .O(n705) );
  ND2X1 U901 ( .I1(n1030), .I2(n744), .O(n767) );
  INVCKX1 U902 ( .I(n774), .O(n189) );
  AN3B2X1 U903 ( .I1(n1057), .B1(n587), .B2(n1139), .O(n1882gat) );
  INVCKX1 U904 ( .I(n772), .O(n188) );
  OR3B2X1 U905 ( .I1(n190), .B1(n983), .B2(n1058), .O(n186) );
  INVCKX1 U906 ( .I(n773), .O(n185) );
  NR2X1 U907 ( .I1(n190), .I2(n667), .O(n773) );
  OR2B1XLP U908 ( .I1(n982), .B1(n1058), .O(n667) );
  OR4B2XLP U909 ( .I1(n747), .I2(n1162), .B1(n1163), .B2(n1059), .O(n1058) );
  ND2X1 U910 ( .I1(n791), .I2(n983), .O(n982) );
  OR4B2XLP U911 ( .I1(n1003), .I2(n1197), .B1(n1161), .B2(n731), .O(n983) );
  ND3X1 U912 ( .I1(n1059), .I2(n736), .I3(n1161), .O(n791) );
  NR2X1 U913 ( .I1(n3099gat), .I2(n651), .O(n1827gat) );
  NR2X1 U914 ( .I1(n1055), .I2(n1056), .O(n1800gat) );
  OR4B2XLP U915 ( .I1(n1187), .I2(n1060), .B1(n733), .B2(n730), .O(n1056) );
  ND2X1 U916 ( .I1(n1190), .I2(n1188), .O(n1060) );
  AN2B1XLP U917 ( .I1(n1061), .B1(n1062), .O(n1793gat) );
  AN2B1XLP U918 ( .I1(n1196), .B1(n778), .O(n3107gat) );
  AN2B1XLP U919 ( .I1(n1771gat), .B1(n715), .O(n778) );
  AN4B1XLP U920 ( .I1(n190), .I2(n902), .I3(n1063), .B1(n905), .O(n3138gat) );
  INVCKX1 U921 ( .I(n989), .O(n905) );
  NR2X1 U922 ( .I1(n1177), .I2(n1179), .O(n989) );
  AN2B1XLP U923 ( .I1(n907), .B1(n695), .O(n1063) );
  NR2X1 U924 ( .I1(n997), .I2(n1178), .O(n902) );
  ND2X1 U925 ( .I1(n859), .I2(n853), .O(n190) );
  OR2B1XLP U926 ( .I1(n1003), .B1(n1064), .O(n853) );
  ND3X1 U927 ( .I1(n1163), .I2(n746), .I3(n1064), .O(n859) );
  NR2X1 U928 ( .I1(n1065), .I2(n774), .O(n1696gat) );
  ND3X1 U929 ( .I1(n1162), .I2(n736), .I3(n1064), .O(n774) );
  NR3X1 U930 ( .I1(n1066), .I2(n1147), .I3(n735), .O(n1636gat) );
  NR3X1 U931 ( .I1(n747), .I2(n731), .I3(n1003), .O(n1620gat) );
  ND2X1 U932 ( .I1(n1162), .I2(n1163), .O(n1003) );
  NR2X1 U933 ( .I1(n1065), .I2(n772), .O(n1613gat) );
  ND3X1 U934 ( .I1(n736), .I2(n746), .I3(n1064), .O(n772) );
  AN2B1XLP U935 ( .I1(n1059), .B1(n1161), .O(n1064) );
  NR2X1 U936 ( .I1(n731), .I2(n1197), .O(n1059) );
  AN2B1XLP U937 ( .I1(n1606gat), .B1(n1065), .O(n1610gat) );
  OAI112X1 U938 ( .C1(n1141), .C2(n676), .A1(n1057), .B1(n1140), .O(n1065) );
  INVCKX1 U939 ( .I(n3100gat), .O(n1044) );
  ND2X1 U940 ( .I1(n1142), .I2(n1821gat), .O(n676) );
  NR2X1 U941 ( .I1(n1197), .I2(n1143), .O(n1606gat) );
  AN3B1X1 U942 ( .I1(n1194), .I2(n1033), .B1(n1054), .O(n1593gat) );
  NR2X1 U943 ( .I1(n1062), .I2(n1034), .O(n1567gat) );
  ND3X1 U944 ( .I1(n761), .I2(n748), .I3(n1018), .O(n1034) );
  NR2X1 U945 ( .I1(n741), .I2(n734), .O(n1018) );
  NR3X1 U946 ( .I1(n1062), .I2(n1054), .I3(n762), .O(n1565gat) );
  ND2X1 U947 ( .I1(n1186), .I2(n734), .O(n762) );
  OR4B2XLP U948 ( .I1(n1187), .I2(n1067), .B1(n733), .B2(n745), .O(n1062) );
  ND2X1 U949 ( .I1(n1190), .I2(n1189), .O(n1067) );
  NR3X1 U950 ( .I1(n1068), .I2(n1038), .I3(n1041), .O(n1564gat) );
  AN4B1XLP U951 ( .I1(n733), .I2(n742), .I3(n1189), .B1(n771), .O(n1041) );
  ND2X1 U952 ( .I1(n1187), .I2(n745), .O(n771) );
  AN4B1XLP U953 ( .I1(n1069), .I2(n1061), .I3(n3149gat), .B1(n1190), .O(n1038)
         );
  ND3X1 U954 ( .I1(n1834gat), .I2(n1767gat), .I3(n1182), .O(n3149gat) );
  OAI12X1 U955 ( .B1(n2989gat), .B2(n1055), .A1(n1068), .O(n1061) );
  ND2X1 U956 ( .I1(n1030), .I2(n761), .O(n1055) );
  NR3X1 U957 ( .I1(n1150), .I2(n1148), .I3(n1186), .O(n1030) );
  MXL2XLP U958 ( .A(n1070), .B(n1071), .S(n1191), .OB(n1069) );
  AOI23X1 U959 ( .B1(n1072), .B2(n1073), .B3(n1074), .A1(n1075), .A2(n1076), 
        .O(n1071) );
  XOR2X1 U960 ( .I1(n743), .I2(n946), .O(n1076) );
  MXL2XLP U961 ( .A(n1077), .B(n1078), .S(n1073), .OB(n1075) );
  OR3B2X1 U962 ( .I1(n1072), .B1(n1188), .B2(n730), .O(n1078) );
  MXL2XLP U963 ( .A(n1032), .B(n1079), .S(n1072), .OB(n1077) );
  NR2X1 U964 ( .I1(n1188), .I2(n730), .O(n1079) );
  NR2X1 U965 ( .I1(n1188), .I2(n1189), .O(n1032) );
  MUXB2X1 U966 ( .EB(n1080), .A(n1081), .B(n1082), .S(n1187), .O(n1074) );
  AN2X1 U967 ( .I1(n1160), .I2(n946), .O(n1082) );
  INVCKX1 U968 ( .I(n946), .O(n1081) );
  ND2X1 U969 ( .I1(n1160), .I2(n751), .O(n946) );
  OR2B1XLP U970 ( .I1(n1145), .B1(n1160), .O(n1073) );
  OR2B1XLP U971 ( .I1(n1144), .B1(n1160), .O(n1072) );
  ND2X1 U972 ( .I1(n1015), .I2(n1187), .O(n1070) );
  INVCKX1 U973 ( .I(n1048), .O(n1068) );
  NR3X1 U974 ( .I1(n744), .I2(n1149), .I3(n1066), .O(n1048) );
  ND3X1 U975 ( .I1(n2989gat), .I2(n741), .I3(n1033), .O(n1066) );
  OAI12X1 U976 ( .B1(n1182), .B2(n1763gat), .A1(n2102gat), .O(n2989gat) );
  AN4B1XLP U977 ( .I1(n1191), .I2(n1187), .I3(n1015), .B1(n1083), .O(n1516gat)
         );
  OR3B2X1 U978 ( .I1(n1054), .B1(n742), .B2(n1033), .O(n1083) );
  NR2X1 U979 ( .I1(n748), .I2(n734), .O(n1033) );
  ND2X1 U980 ( .I1(n761), .I2(n741), .O(n1054) );
  NR2X1 U981 ( .I1(n744), .I2(n735), .O(n761) );
  INVCKX1 U982 ( .I(n1080), .O(n1015) );
  ND2X1 U983 ( .I1(n1189), .I2(n1188), .O(n1080) );
  AN4B1XLP U984 ( .I1(n907), .I2(n1181), .I3(n991), .B1(n993), .O(n1391gat) );
  ND2X1 U985 ( .I1(n968), .I2(n1178), .O(n993) );
  INVCKX1 U986 ( .I(n997), .O(n968) );
  ND2X1 U987 ( .I1(n1176), .I2(n1175), .O(n997) );
  NR2X1 U988 ( .I1(n690), .I2(n1179), .O(n991) );
  AN4B1XLP U989 ( .I1(n1215), .I2(n1214), .I3(n1180), .B1(n1151), .O(n907) );
  XOR2X1 U990 ( .I1(n1084), .I2(n1085), .O(n3116gat) );
  XOR4XLP U991 ( .I1(n1154), .I2(n1155), .I3(n1152), .I4(n1153), .O(n1085) );
  XOR4XLP U992 ( .I1(n1156), .I2(n1157), .I3(n752), .I4(n1158), .O(n1084) );
endmodule

