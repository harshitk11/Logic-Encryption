
module s15850 ( clk, g18, g27, g109, g741, g742, g743, g744, g872, g873, g877, 
        g881, g1712, g1960, g1961, g1696, g750, g85, g42, g1700, g102, g104, 
        g101, g29, g28, g103, g83, g23, g87, g922, g892, g84, g919, g1182, 
        g925, g48, g895, g889, g1185, g41, g43, g99, g1173, g1203, g1188, 
        g1197, g46, g31, g45, g92, g89, g898, g91, g93, g913, g82, g88, g1194, 
        g47, g96, g910, g95, g904, g1176, g901, g44, g916, g100, g886, g30, 
        g86, g1170, g1200, g1191, g907, g90, g94, g1179, g2355, g2601, g2602, 
        g2603, g2604, g2605, g2606, g2607, g2608, g2609, g2610, g2611, g2612, 
        g2648, g2986, g3007, g3069, g4172, g4173, g4174, g4175, g4176, g4177, 
        g4178, g4179, g4180, g4181, g4887, g4888, g5101, g5105, g5658, g5659, 
        g5816, g6920, g6926, g6932, g6942, g6949, g6955, g7744, g8061, g8062, 
        g8271, g8313, g8316, g8318, g8323, g8328, g8331, g8335, g8340, g8347, 
        g8349, g8352, g8561, g8562, g8563, g8564, g8565, g8566, g8976, g8977, 
        g8978, g8979, g8980, g8981, g8982, g8983, g8984, g8985, g8986, g9451, 
        g9961, g10377, g10379, g10455, g10457, g10459, g10461, g10463, g10465, 
        g10628, g10801, g11163, g11206, g11489, g6842, g4171, g6267, g6257, 
        g1957, g6282, g6284, g6281, g6253, g6285, g6283, g6265, g3327, g6269, 
        g4204, g4193, g6266, g4203, g4212, g4196, g6263, g4194, g4192, g4213, 
        g6256, g6258, g6279, g4209, g4208, g4214, g4206, g6261, g6255, g6260, 
        g6274, g6271, g4195, g6273, g6275, g4201, g6264, g6270, g4216, g6262, 
        g6278, g4200, g6277, g4198, g4210, g4197, g6259, g4202, g6280, g4191, 
        g6254, g6268, g4205, g4207, g4215, g4199, g6272, g6276, g4211, test_si, 
        test_se );
  input clk, g18, g27, g109, g741, g742, g743, g744, g872, g873, g877, g881,
         g1712, g1960, g1961, g1696, g750, g85, g42, g1700, g102, g104, g101,
         g29, g28, g103, g83, g23, g87, g922, g892, g84, g919, g1182, g925,
         g48, g895, g889, g1185, g41, g43, g99, g1173, g1203, g1188, g1197,
         g46, g31, g45, g92, g89, g898, g91, g93, g913, g82, g88, g1194, g47,
         g96, g910, g95, g904, g1176, g901, g44, g916, g100, g886, g30, g86,
         g1170, g1200, g1191, g907, g90, g94, g1179, test_si, test_se;
  output g2355, g2601, g2602, g2603, g2604, g2605, g2606, g2607, g2608, g2609,
         g2610, g2611, g2612, g2648, g2986, g3007, g3069, g4172, g4173, g4174,
         g4175, g4176, g4177, g4178, g4179, g4180, g4181, g4887, g4888, g5101,
         g5105, g5658, g5659, g5816, g6920, g6926, g6932, g6942, g6949, g6955,
         g7744, g8061, g8062, g8271, g8313, g8316, g8318, g8323, g8328, g8331,
         g8335, g8340, g8347, g8349, g8352, g8561, g8562, g8563, g8564, g8565,
         g8566, g8976, g8977, g8978, g8979, g8980, g8981, g8982, g8983, g8984,
         g8985, g8986, g9451, g9961, g10377, g10379, g10455, g10457, g10459,
         g10461, g10463, g10465, g10628, g10801, g11163, g11206, g11489, g6842,
         g4171, g6267, g6257, g1957, g6282, g6284, g6281, g6253, g6285, g6283,
         g6265, g3327, g6269, g4204, g4193, g6266, g4203, g4212, g4196, g6263,
         g4194, g4192, g4213, g6256, g6258, g6279, g4209, g4208, g4214, g4206,
         g6261, g6255, g6260, g6274, g6271, g4195, g6273, g6275, g4201, g6264,
         g6270, g4216, g6262, g6278, g4200, g6277, g4198, g4210, g4197, g6259,
         g4202, g6280, g4191, g6254, g6268, g4205, g4207, g4215, g4199, g6272,
         g6276, g4211;
  wire   g18, g27, g872, g873, g1960, g1961, g85, g42, g102, g104, g101, g29,
         g28, g103, g83, g87, g922, g892, g84, g919, g1182, g925, g48, g895,
         g889, g1185, g41, g43, g99, g1173, g1203, g1188, g1197, g46, g31, g45,
         g92, g89, g898, g91, g93, g913, g82, g88, g1194, g47, g96, g910, g95,
         g904, g1176, g901, g44, g916, g100, g886, g30, g86, g1170, g1200,
         g1191, g907, g90, g94, g1179, g1736, g1737, g1956, g113, g745, g822,
         g632, g16, g806, g1217, g756, g1713, g814, g259, g1317, g262, g1356,
         g794, g261, g254, g1850, g17, g8, g255, g1955, g746, g1854, g1958,
         g1765, g826, g257, g874, g636, g818, g802, g810, g253, g875, g798,
         g114, g260, g258, g755, g256, g1360, g8244, g6829, g4334, g6733,
         g9266, g6819, g10782, g6215, g8254, g3506, g8769, g4500, g4477, g6828,
         g6830, g8765, g6198, g6747, g4903, g8245, g9272, g6821, g8768, g11639,
         g6841, g11391, g6757, g11340, g4338, g5543, g6234, g4498, g11372,
         g6823, g11320, g6193, g7581, g6834, g5770, g11641, g11292, g7032,
         g6525, g8046, g4940, g8047, g9555, g6180, g6832, g6123, g5755, g5445,
         g5173, g6839, g8260, g10785, g6334, g6621, g7709, g11640, g4890,
         g4480, g6179, g7590, g11380, g7930, g10784, g6332, g7705, g9269,
         g5421, g8040, g6838, g6795, g6205, g3381, g6983, g5126, g8050, g6679,
         g6831, g6653, g11393, g6786, g4484, g7137, g5390, g8384, g6759, g8024,
         g6833, g4892, g9721, g4340, g8044, g6728, g11392, g6331, g4471, g8042,
         g8054, g6502, g6216, g6826, g7191, g6638, g6827, g6333, g8049, g8019,
         g8052, g5194, g4473, g8766, g5918, g8045, g8173, g11349, g7843, g6531,
         g8059, g8767, g4114, g11636, g7586, g4465, g6126, g4891, g10780,
         g4342, g8048, g8055, g6508, g6820, g8041, g6840, g7134, g8772, g4893,
         g8505, g6163, g7202, g4325, g11514, g4904, g11291, g6627, g7541,
         g6526, g8051, g6439, g9110, g8043, g4330, g8147, g6224, g4902, g4490,
         g6516, g8820, g8775, g5083, g8060, g6244, g9150, g6656, g5536, g6824,
         g8250, g8053, g4506, g6471, g7632, g11290, g8039, g5529, g5148, g9124,
         g6822, g4905, g11376, g6895, g7189, g7297, g8771, g11625, g8945,
         g11338, g8435, g6911, g10865, g6469, g11257, g6898, g6900, g4264,
         g6088, g6923, g8194, g11256, g11300, g4238, g8773, g10864, g6934,
         g6096, g11314, g8921, g11269, g11268, g6481, g11335, g11487, g8941,
         g11443, g4231, g8431, g7133, g11306, g5996, g8286, g7290, g6068,
         g6468, g11478, g11486, g8287, g6524, g7257, g7301, g11334, g8923,
         g7441, g6026, g10799, g10798, g8943, g11293, g11265, g8887, g6514,
         g8433, g11579, g10771, g6522, g7183, g6537, g4309, g6243, g6542,
         g7303, g6902, g6529, g11264, g10795, g11607, g9961, g6926, g7294,
         g6909, g4283, g8939, g11327, g11606, g11303, g6506, g7626, g10770,
         g11483, g6545, g10767, g11326, g10898, g6507, g10718, g7292, g10861,
         g6515, g6528, g8649, g10776, g10859, g7299, g10858, g8193, g7244,
         g8563, g6908, g8938, g5910, g11482, g11647, g5396, g11331, g7295,
         g6541, g8284, g6901, g8559, g10860, g8973, g11310, g6500, g10855,
         g11603, g6672, g6523, g10707, g7298, g6551, g6099, g8282, g7219,
         g11298, g10866, g6534, g8776, g11261, g6513, g6916, g8777, g7291,
         g11330, g10773, g6042, g11259, g5914, g11258, g6054, g11602, g11337,
         g8889, g8285, g10791, g6049, g11336, g8926, g7293, g10800, g11308,
         g10936, g6470, g6897, g8885, g11260, g11488, g4556, g8288, g6755,
         g11610, g6045, g11270, g6059, g11267, g11294, g5404, g4089, g6015,
         g8770, g11266, g10863, g8429, g8281, g6910, g11305, g6538, g6093,
         g11485, g10797, g6949, g10711, g8283, g8920, g10862, g11333, g6080,
         g6480, g11484, g11609, g8940, g11312, g11608, g6000, g8428, g8430,
         g8566, g6924, g8883, g11329, g4255, g11328, g8774, g7204, g7300,
         g4293, g6533, g8564, g8631, g6922, g11263, g11332, g7143, g6479,
         g6501, g6920, g11605, g4274, g10717, g6912, g6929, g11325, g6894,
         g8779, g10793, g8944, g10765, g11604, g8434, g6546, g11262, g6906,
         g11324, g8922, g6478, g6907, g6035, g8937, g6915, g6002, g8432, g6928,
         g6930, g7660, g6071, g7302, g6038, g4239, g6918, g11481, g7296, g4117,
         g3524, g2478, g4076, g6155, g5556, g5392, g3462, n519, n523, n526,
         n527, n533, n540, n541, n546, n547, n552, n569, n577, n578, n592,
         n681, n1405, n1417, n1426, n1431, n1434, n1448, n1500, n1508, n1525,
         n1549, n1576, n1584, n1591, n1594, n1595, n1606, n1614, n1620, n1651,
         n1661, n1672, n1674, n1676, n1688, n1707, n1719, n1724, n1727, n1731,
         n1738, n1742, n1743, n1768, n1794, n1812, n1823, n1834, n1836, n1861,
         g8271, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323;
  assign g2355 = g18;
  assign g7744 = g27;
  assign g8061 = g872;
  assign g5101 = g872;
  assign g5105 = g873;
  assign g8062 = g873;
  assign g4888 = g1960;
  assign g4887 = g1961;
  assign g6267 = g85;
  assign g6257 = g42;
  assign g6282 = g102;
  assign g6284 = g104;
  assign g6281 = g101;
  assign g6253 = g29;
  assign g6285 = g28;
  assign g6283 = g103;
  assign g6265 = g83;
  assign g6269 = g87;
  assign g4204 = g922;
  assign g4193 = g892;
  assign g6266 = g84;
  assign g4203 = g919;
  assign g4212 = g1182;
  assign g4196 = g925;
  assign g6263 = g48;
  assign g4194 = g895;
  assign g4192 = g889;
  assign g4213 = g1185;
  assign g6256 = g41;
  assign g6258 = g43;
  assign g6279 = g99;
  assign g4209 = g1173;
  assign g4208 = g1203;
  assign g4214 = g1188;
  assign g4206 = g1197;
  assign g6261 = g46;
  assign g6255 = g31;
  assign g6260 = g45;
  assign g6274 = g92;
  assign g6271 = g89;
  assign g4195 = g898;
  assign g6273 = g91;
  assign g6275 = g93;
  assign g4201 = g913;
  assign g6264 = g82;
  assign g6270 = g88;
  assign g4216 = g1194;
  assign g6262 = g47;
  assign g6278 = g96;
  assign g4200 = g910;
  assign g6277 = g95;
  assign g4198 = g904;
  assign g4210 = g1176;
  assign g4197 = g901;
  assign g6259 = g44;
  assign g4202 = g916;
  assign g6280 = g100;
  assign g4191 = g886;
  assign g6254 = g30;
  assign g6268 = g86;
  assign g4205 = g1170;
  assign g4207 = g1200;
  assign g4215 = g1191;
  assign g4199 = g907;
  assign g6272 = g90;
  assign g6276 = g94;
  assign g4211 = g1179;
  assign g9451 = g9961;
  assign g8562 = g6926;
  assign g6932 = g8563;
  assign g8565 = g6949;
  assign g6955 = g8566;
  assign g6942 = g8564;
  assign g8561 = g6920;
  assign g5816 = g8271;

  DFZX1 gate1 ( .D(g4556), .TD(test_si), .SEL(test_se), .CK(clk), .Q(n2974) );
  DFZX1 gate2 ( .D(g8943), .TD(n2974), .SEL(test_se), .CK(clk), .Q(n3119), 
        .QB(n1878) );
  DFZX1 gate3 ( .D(g255), .TD(n3119), .SEL(test_se), .CK(clk), .Q(n3040) );
  DFZX1 gate4 ( .D(g11257), .TD(n3040), .SEL(test_se), .CK(clk), .Q(n3323), 
        .QB(n1915) );
  DFZX1 gate5 ( .D(g7032), .TD(n3323), .SEL(test_se), .CK(clk), .Q(n3105), 
        .QB(n2100) );
  DFZX1 gate6 ( .D(g6830), .TD(n3105), .SEL(test_se), .CK(clk), .Q(n3120), 
        .QB(n2061) );
  DFZX1 gate7 ( .D(g8920), .TD(n3120), .SEL(test_se), .CK(clk), .Q(n2889) );
  DFZX1 gate8 ( .D(g4340), .TD(n2889), .SEL(test_se), .CK(clk), .Q(n3121) );
  DFZX1 gate10 ( .D(g4239), .TD(n3121), .SEL(test_se), .CK(clk), .Q(n3103) );
  DFZX1 gate11 ( .D(g6538), .TD(n3103), .SEL(test_se), .CK(clk), .Q(n3322), 
        .QB(n1886) );
  DFZX1 gate12 ( .D(g8887), .TD(n3322), .SEL(test_se), .CK(clk), .Q(n3122) );
  DFZX1 gate13 ( .D(g11372), .TD(n3122), .SEL(test_se), .CK(clk), .Q(n3123), 
        .QB(n1873) );
  DFZX1 gate14 ( .D(g8260), .TD(n3123), .SEL(test_se), .CK(clk), .Q(n3124) );
  DFZX1 gate15 ( .D(g11391), .TD(n3124), .SEL(test_se), .CK(clk), .Q(n3125) );
  DFZX1 gate16 ( .D(g8432), .TD(n3125), .SEL(test_se), .CK(clk), .Q(n2893), 
        .QB(n2029) );
  DFZX1 gate17 ( .D(g6088), .TD(n2893), .SEL(test_se), .CK(clk), .Q(n2932) );
  DFZX1 gate18 ( .D(g6478), .TD(n2932), .SEL(test_se), .CK(clk), .Q(n3086) );
  DFZX1 gate19 ( .D(g6795), .TD(n3086), .SEL(test_se), .CK(clk), .Q(n2992) );
  DFZX1 gate20 ( .D(g11320), .TD(n2992), .SEL(test_se), .CK(clk), .Q(n3030) );
  DFZX1 gate21 ( .D(g6500), .TD(n3030), .SEL(test_se), .CK(clk), .Q(n3321), 
        .QB(n2057) );
  DFZX1 gate22 ( .D(g5392), .TD(n3321), .SEL(test_se), .CK(clk), .Q(g1736) );
  DFZX1 gate23 ( .D(n547), .TD(g1736), .SEL(test_se), .CK(clk), .Q(n3113) );
  DFZX1 gate24 ( .D(g10782), .TD(n3113), .SEL(test_se), .CK(clk), .Q(n3320), 
        .QB(n1952) );
  DFZX1 gate25 ( .D(g6216), .TD(n3320), .SEL(test_se), .CK(clk), .Q(n3319), 
        .QB(n2010) );
  DFZX1 gate26 ( .D(g1736), .TD(n3319), .SEL(test_se), .CK(clk), .Q(g1737) );
  DFZX1 gate27 ( .D(g10858), .TD(g1737), .SEL(test_se), .CK(clk), .Q(n3318), 
        .QB(n2052) );
  DFZX1 gate28 ( .D(g5914), .TD(n3318), .SEL(test_se), .CK(clk), .Q(n3317), 
        .QB(n1936) );
  DFZX1 gate29 ( .D(g7590), .TD(n3317), .SEL(test_se), .CK(clk), .Q(n2977) );
  DFZX1 gate30 ( .D(g6656), .TD(n2977), .SEL(test_se), .CK(clk), .Q(n3090), 
        .QB(n2101) );
  DFZX1 gate31 ( .D(g6728), .TD(n3090), .SEL(test_se), .CK(clk), .Q(g4177), 
        .QB(n1719) );
  DFZX1 gate32 ( .D(g5126), .TD(g4177), .SEL(test_se), .CK(clk), .Q(n3126), 
        .QB(n1893) );
  DFZX1 gate33 ( .D(g7290), .TD(n3126), .SEL(test_se), .CK(clk), .Q(n3316), 
        .QB(n1914) );
  DFZX1 gate34 ( .D(g6841), .TD(n3316), .SEL(test_se), .CK(clk), .Q(n3052) );
  DFZX1 gate35 ( .D(g8041), .TD(n3052), .SEL(test_se), .CK(clk), .Q(n2939) );
  DFZX1 gate37 ( .D(g8766), .TD(n2939), .SEL(test_se), .CK(clk), .Q(n2917), 
        .QB(n2034) );
  DFZX1 gate38 ( .D(n523), .TD(n2917), .SEL(test_se), .CK(clk), .Q(n3315), 
        .QB(n3062) );
  DFZX1 gate39 ( .D(g8019), .TD(n3315), .SEL(test_se), .CK(clk), .Q(g4180), 
        .QB(n1661) );
  DFZX1 gate40 ( .D(g6545), .TD(g4180), .SEL(test_se), .CK(clk), .Q(n3115) );
  DFZX1 gate42 ( .D(g256), .TD(n3115), .SEL(test_se), .CK(clk), .Q(n3029) );
  DFZX1 gate43 ( .D(g6533), .TD(n3029), .SEL(test_se), .CK(clk), .Q(n3079) );
  DFZX1 gate44 ( .D(g8820), .TD(n3079), .SEL(test_se), .CK(clk), .Q(n3127), 
        .QB(n1971) );
  DFZX1 gate45 ( .D(g8941), .TD(n3127), .SEL(test_se), .CK(clk), .Q(n2886) );
  DFZX1 gate46 ( .D(g10859), .TD(n2886), .SEL(test_se), .CK(clk), .Q(n3314), 
        .QB(n1940) );
  DFZX1 gate47 ( .D(g6922), .TD(n3314), .SEL(test_se), .CK(clk), .Q(n3070) );
  DFZX1 gate48 ( .D(g8772), .TD(n3070), .SEL(test_se), .CK(clk), .Q(n2919), 
        .QB(n1885) );
  DFZX1 gate49 ( .D(g8433), .TD(n2919), .SEL(test_se), .CK(clk), .Q(n3313), 
        .QB(n1882) );
  DFZX1 gate50 ( .D(g6526), .TD(n3313), .SEL(test_se), .CK(clk), .Q(g8985), 
        .QB(n2047) );
  DFZX1 gate51 ( .D(g10793), .TD(g8985), .SEL(test_se), .CK(clk), .Q(n3312), 
        .QB(n2020) );
  DFZX1 gate52 ( .D(g11333), .TD(n3312), .SEL(test_se), .CK(clk), .Q(n2991), 
        .QB(n1974) );
  DFZX1 gate53 ( .D(g11392), .TD(n2991), .SEL(test_se), .CK(clk), .Q(n3128), 
        .QB(n1969) );
  DFZX1 gate54 ( .D(g3506), .TD(n3128), .SEL(test_se), .CK(clk), .Q(g3007), 
        .QB(n3064) );
  DFZX1 gate55 ( .D(g1713), .TD(g3007), .SEL(test_se), .CK(clk), .Q(n2947) );
  DFZX1 gate56 ( .D(g794), .TD(n2947), .SEL(test_se), .CK(clk), .Q(n3027) );
  DFZX1 gate57 ( .D(g6093), .TD(n3027), .SEL(test_se), .CK(clk), .Q(n2931) );
  DFZX1 gate58 ( .D(g8889), .TD(n2931), .SEL(test_se), .CK(clk), .Q(n2891), 
        .QB(n1965) );
  DFZX1 gate59 ( .D(g7302), .TD(n2891), .SEL(test_se), .CK(clk), .Q(n3311), 
        .QB(n1879) );
  DFZX1 gate60 ( .D(g6525), .TD(n3311), .SEL(test_se), .CK(clk), .Q(n3187), 
        .QB(n1874) );
  DFZX1 gate61 ( .D(g8429), .TD(n3187), .SEL(test_se), .CK(clk), .Q(n3129), 
        .QB(n1927) );
  DFZX1 gate62 ( .D(g7292), .TD(n3129), .SEL(test_se), .CK(clk), .Q(n2980), 
        .QB(n1921) );
  DFZX1 gate63 ( .D(g104), .TD(n2980), .SEL(test_se), .CK(clk), .Q(g2602) );
  DFZX1 gate64 ( .D(g6621), .TD(g2602), .SEL(test_se), .CK(clk), .Q(g8977), 
        .QB(n2045) );
  DFZX1 gate65 ( .D(g7134), .TD(g8977), .SEL(test_se), .CK(clk), .Q(n3130) );
  DFZX1 gate66 ( .D(g260), .TD(n3130), .SEL(test_se), .CK(clk), .Q(n3043) );
  DFZX1 gate67 ( .D(g6333), .TD(n3043), .SEL(test_se), .CK(clk), .Q(n3131), 
        .QB(n2025) );
  DFZX1 gate68 ( .D(g6826), .TD(n3131), .SEL(test_se), .CK(clk), .Q(n3310), 
        .QB(n1944) );
  DFZX1 gate69 ( .D(g1955), .TD(n3310), .SEL(test_se), .CK(clk), .Q(g1956) );
  DFZX1 gate70 ( .D(g10860), .TD(g1956), .SEL(test_se), .CK(clk), .Q(n3309), 
        .QB(n2051) );
  DFZX1 gate71 ( .D(g11483), .TD(n3309), .SEL(test_se), .CK(clk), .Q(n2970), 
        .QB(n2088) );
  DFZX1 gate72 ( .D(n577), .TD(n2970), .SEL(test_se), .CK(clk), .Q(g113) );
  DFZX1 gate73 ( .D(g7626), .TD(g113), .SEL(test_se), .CK(clk), .Q(n3132) );
  DFZX1 gate74 ( .D(g10866), .TD(n3132), .SEL(test_se), .CK(clk), .Q(n3308), 
        .QB(n2048) );
  DFZX1 gate75 ( .D(g8193), .TD(n3308), .SEL(test_se), .CK(clk), .Q(n3307), 
        .QB(n2021) );
  DFZX1 gate76 ( .D(g6983), .TD(n3307), .SEL(test_se), .CK(clk), .Q(n2996), 
        .QB(n1920) );
  DFZX1 gate77 ( .D(g6839), .TD(n2996), .SEL(test_se), .CK(clk), .Q(n3012), 
        .QB(n1907) );
  DFZX1 gate78 ( .D(g4076), .TD(n3012), .SEL(test_se), .CK(clk), .Q(n2949) );
  DFZX1 gate79 ( .D(g4293), .TD(n2949), .SEL(test_se), .CK(clk), .Q(n3066) );
  DFZX1 gate80 ( .D(g11482), .TD(n3066), .SEL(test_se), .CK(clk), .Q(n2971), 
        .QB(n2089) );
  DFZX1 gate81 ( .D(g1956), .TD(n2971), .SEL(test_se), .CK(clk), .Q(g1957) );
  DFZX1 gate82 ( .D(g6507), .TD(g1957), .SEL(test_se), .CK(clk), .Q(n3306), 
        .QB(n1930) );
  DFZX1 gate83 ( .D(g6096), .TD(n3306), .SEL(test_se), .CK(clk), .Q(n2930) );
  DFZX1 gate84 ( .D(g8250), .TD(n2930), .SEL(test_se), .CK(clk), .Q(n3092) );
  DFZX1 gate86 ( .D(g8282), .TD(n3092), .SEL(test_se), .CK(clk), .Q(n2897), 
        .QB(n2005) );
  DFZX1 gate87 ( .D(g8435), .TD(n2897), .SEL(test_se), .CK(clk), .Q(n3133), 
        .QB(n2077) );
  DFZX1 gate88 ( .D(g6924), .TD(n3133), .SEL(test_se), .CK(clk), .Q(n3005) );
  DFZX1 gate89 ( .D(g6819), .TD(n3005), .SEL(test_se), .CK(clk), .Q(n3305), 
        .QB(n2064) );
  DFZX1 gate90 ( .D(g746), .TD(n3305), .SEL(test_se), .CK(clk), .Q(g745) );
  DFZX1 gate91 ( .D(g6244), .TD(g745), .SEL(test_se), .CK(clk), .Q(n2962) );
  DFZX1 gate92 ( .D(g6627), .TD(n2962), .SEL(test_se), .CK(clk), .Q(g8979), 
        .QB(n2044) );
  DFZX1 gate93 ( .D(n526), .TD(g8979), .SEL(test_se), .CK(clk), .Q(n3304), 
        .QB(n3056) );
  DFZX1 gate94 ( .D(g3007), .TD(n3304), .SEL(test_se), .CK(clk), .Q(n3063) );
  DFZX1 gate95 ( .D(g6071), .TD(n3063), .SEL(test_se), .CK(clk), .Q(n2934) );
  DFZX1 gate96 ( .D(g8046), .TD(n2934), .SEL(test_se), .CK(clk), .Q(n3303), 
        .QB(n1910) );
  DFZX1 gate97 ( .D(g10707), .TD(n3303), .SEL(test_se), .CK(clk), .Q(n3302), 
        .QB(n1950) );
  DFZX1 gate98 ( .D(g6198), .TD(n3302), .SEL(test_se), .CK(clk), .Q(n2928) );
  DFZX1 gate99 ( .D(g8051), .TD(n2928), .SEL(test_se), .CK(clk), .Q(n3301), 
        .QB(n1909) );
  DFZX1 gate100 ( .D(g8024), .TD(n3301), .SEL(test_se), .CK(clk), .Q(g822), 
        .QB(n1614) );
  DFZX1 gate101 ( .D(g29), .TD(g822), .SEL(test_se), .CK(clk), .Q(g2609) );
  DFZX1 gate102 ( .D(g10862), .TD(g2609), .SEL(test_se), .CK(clk), .Q(n3300), 
        .QB(n2050) );
  DFZX1 gate103 ( .D(g8050), .TD(n3300), .SEL(test_se), .CK(clk), .Q(n2902), 
        .QB(n2009) );
  DFZX1 gate104 ( .D(g7133), .TD(n2902), .SEL(test_se), .CK(clk), .Q(n2993), 
        .QB(n1901) );
  DFZX1 gate105 ( .D(g7930), .TD(n2993), .SEL(test_se), .CK(clk), .Q(n2995) );
  DFZX1 gate106 ( .D(g6832), .TD(n2995), .SEL(test_se), .CK(clk), .Q(n3019) );
  DFZX1 gate107 ( .D(g11308), .TD(n3019), .SEL(test_se), .CK(clk), .Q(n3083)
         );
  DFZX1 gate109 ( .D(g6918), .TD(n3083), .SEL(test_se), .CK(clk), .Q(n3008) );
  DFZX1 gate110 ( .D(g8769), .TD(n3008), .SEL(test_se), .CK(clk), .Q(n2927), 
        .QB(n2032) );
  DFZX1 gate112 ( .D(g6909), .TD(n2927), .SEL(test_se), .CK(clk), .Q(n3299), 
        .QB(n2002) );
  DFZX1 gate113 ( .D(g4940), .TD(n3299), .SEL(test_se), .CK(clk), .Q(g4173), 
        .QB(n1836) );
  DFZX1 gate114 ( .D(g5404), .TD(g4173), .SEL(test_se), .CK(clk), .Q(n3134), 
        .QB(n1958) );
  DFZX1 gate115 ( .D(g11265), .TD(n3134), .SEL(test_se), .CK(clk), .Q(n3298), 
        .QB(n1875) );
  DFZX1 gate116 ( .D(g6930), .TD(n3298), .SEL(test_se), .CK(clk), .Q(n3006) );
  DFZX1 gate117 ( .D(n552), .TD(n3006), .SEL(test_se), .CK(clk), .Q(n3068) );
  DFZX1 gate118 ( .D(g4891), .TD(n3068), .SEL(test_se), .CK(clk), .Q(g632) );
  DFZX1 gate119 ( .D(g6224), .TD(g632), .SEL(test_se), .CK(clk), .Q(n2964) );
  DFZX1 gate120 ( .D(g7586), .TD(n2964), .SEL(test_se), .CK(clk), .Q(n2976) );
  DFZX1 gate121 ( .D(g10770), .TD(n2976), .SEL(test_se), .CK(clk), .Q(n3297), 
        .QB(n2069) );
  DFZX1 gate122 ( .D(g2986), .TD(n3297), .SEL(test_se), .CK(clk), .Q(n3296), 
        .QB(n1834) );
  DFZX1 gate123 ( .D(g3524), .TD(n3296), .SEL(test_se), .CK(clk), .Q(g16) );
  DFZX1 gate124 ( .D(g6934), .TD(g16), .SEL(test_se), .CK(clk), .Q(n3109) );
  DFZX1 gate125 ( .D(g11256), .TD(n3109), .SEL(test_se), .CK(clk), .Q(n3295), 
        .QB(n1957) );
  DFZX1 gate126 ( .D(g6824), .TD(n3295), .SEL(test_se), .CK(clk), .Q(n3016), 
        .QB(n2070) );
  DFZX1 gate127 ( .D(g1360), .TD(n3016), .SEL(test_se), .CK(clk), .Q(n3294), 
        .QB(n1606) );
  DFZX1 gate128 ( .D(g6126), .TD(n3294), .SEL(test_se), .CK(clk), .Q(g806), 
        .QB(n1707) );
  DFZX1 gate129 ( .D(g8767), .TD(g806), .SEL(test_se), .CK(clk), .Q(n2915) );
  DFZX1 gate130 ( .D(g102), .TD(n2915), .SEL(test_se), .CK(clk), .Q(g2605) );
  DFZX1 gate131 ( .D(g6546), .TD(g2605), .SEL(test_se), .CK(clk), .Q(n3065) );
  DFZX1 gate132 ( .D(g4238), .TD(n3065), .SEL(test_se), .CK(clk), .Q(n3110), 
        .QB(n2095) );
  DFZX1 gate133 ( .D(g6823), .TD(n3110), .SEL(test_se), .CK(clk), .Q(n3014), 
        .QB(n1943) );
  DFZX1 gate134 ( .D(g6928), .TD(n3014), .SEL(test_se), .CK(clk), .Q(n3293), 
        .QB(n1933) );
  DFZX1 gate135 ( .D(g11602), .TD(n3293), .SEL(test_se), .CK(clk), .Q(n3135)
         );
  DFZX1 gate136 ( .D(g9721), .TD(n3135), .SEL(test_se), .CK(clk), .Q(n3136), 
        .QB(n1963) );
  DFZX1 gate137 ( .D(g4890), .TD(n3136), .SEL(test_se), .CK(clk), .Q(n3292), 
        .QB(n1508) );
  DFZX1 gate138 ( .D(n1867), .TD(n3292), .SEL(test_se), .CK(clk), .Q(g1217) );
  DFZX1 gate139 ( .D(g6524), .TD(g1217), .SEL(test_se), .CK(clk), .Q(n3111) );
  DFZX1 gate140 ( .D(g8045), .TD(n3111), .SEL(test_se), .CK(clk), .Q(n3291), 
        .QB(n1985) );
  DFZX1 gate141 ( .D(g6469), .TD(n3291), .SEL(test_se), .CK(clk), .Q(n3095) );
  DFZX1 gate142 ( .D(g6471), .TD(n3095), .SEL(test_se), .CK(clk), .Q(n3137) );
  DFZX1 gate143 ( .D(g6821), .TD(n3137), .SEL(test_se), .CK(clk), .Q(n3290), 
        .QB(n1888) );
  DFZX1 gate144 ( .D(g11514), .TD(n3290), .SEL(test_se), .CK(clk), .Q(n2961)
         );
  DFZX1 gate146 ( .D(g4480), .TD(n2961), .SEL(test_se), .CK(clk), .Q(n3184) );
  DFZX1 gate147 ( .D(g11610), .TD(n3184), .SEL(test_se), .CK(clk), .Q(n3138)
         );
  DFZX1 gate148 ( .D(g7843), .TD(n3138), .SEL(test_se), .CK(clk), .Q(n2924), 
        .QB(n1883) );
  DFZX1 gate149 ( .D(g11310), .TD(n2924), .SEL(test_se), .CK(clk), .Q(n3075), 
        .QB(n2081) );
  DFZX1 gate150 ( .D(g5536), .TD(n3075), .SEL(test_se), .CK(clk), .Q(g4175), 
        .QB(n1724) );
  DFZX1 gate151 ( .D(g28), .TD(g4175), .SEL(test_se), .CK(clk), .Q(g2603) );
  DFZX1 gate152 ( .D(g11331), .TD(g2603), .SEL(test_se), .CK(clk), .Q(n3289), 
        .QB(n1959) );
  DFZX1 gate153 ( .D(g11380), .TD(n3289), .SEL(test_se), .CK(clk), .Q(n3139), 
        .QB(n1955) );
  DFZX1 gate154 ( .D(g6838), .TD(n3139), .SEL(test_se), .CK(clk), .Q(n2945) );
  DFZX1 gate155 ( .D(g103), .TD(n2945), .SEL(test_se), .CK(clk), .Q(g2606) );
  DFZX1 gate156 ( .D(g8288), .TD(g2606), .SEL(test_se), .CK(clk), .Q(n3140), 
        .QB(n2006) );
  DFZX1 gate157 ( .D(g755), .TD(n3140), .SEL(test_se), .CK(clk), .Q(g756) );
  DFZX1 gate158 ( .D(g4892), .TD(g756), .SEL(test_se), .CK(clk), .Q(n3288), 
        .QB(n1525) );
  DFZX1 gate159 ( .D(g5390), .TD(n3288), .SEL(test_se), .CK(clk), .Q(n3141), 
        .QB(n1891) );
  DFZX1 gate160 ( .D(g10855), .TD(n3141), .SEL(test_se), .CK(clk), .Q(n3287), 
        .QB(n2053) );
  DFZX1 gate162 ( .D(g10898), .TD(n3287), .SEL(test_se), .CK(clk), .Q(n3059), 
        .QB(n2092) );
  DFZX1 gate163 ( .D(g10865), .TD(n3059), .SEL(test_se), .CK(clk), .Q(n3286), 
        .QB(n1937) );
  DFZX1 gate164 ( .D(g6822), .TD(n3286), .SEL(test_se), .CK(clk), .Q(n3285), 
        .QB(n1951) );
  DFZX1 gate165 ( .D(g6528), .TD(n3285), .SEL(test_se), .CK(clk), .Q(n3085) );
  DFZX1 gate166 ( .D(g6180), .TD(n3085), .SEL(test_se), .CK(clk), .Q(n2913) );
  DFZX1 gate167 ( .D(g10718), .TD(n2913), .SEL(test_se), .CK(clk), .Q(n3050), 
        .QB(n2094) );
  DFZX1 gate168 ( .D(g6912), .TD(n3050), .SEL(test_se), .CK(clk), .Q(n3007) );
  DFZX1 gate169 ( .D(n527), .TD(n3007), .SEL(test_se), .CK(clk), .Q(n3284), 
        .QB(n1431) );
  DFZX1 gate170 ( .D(g6234), .TD(n3284), .SEL(test_se), .CK(clk), .Q(n3283), 
        .QB(n1919) );
  DFZX1 gate171 ( .D(g6099), .TD(n3283), .SEL(test_se), .CK(clk), .Q(n2929) );
  DFZX1 gate172 ( .D(g11259), .TD(n2929), .SEL(test_se), .CK(clk), .Q(n3031), 
        .QB(n1926) );
  DFZX1 gate173 ( .D(g8039), .TD(n3031), .SEL(test_se), .CK(clk), .Q(n2916) );
  DFZX1 gate174 ( .D(g6059), .TD(n2916), .SEL(test_se), .CK(clk), .Q(n2936) );
  DFZX1 gate175 ( .D(g5396), .TD(n2936), .SEL(test_se), .CK(clk), .Q(g1713), 
        .QB(n1823) );
  DFZX1 gate176 ( .D(g262), .TD(g1713), .SEL(test_se), .CK(clk), .Q(n3042) );
  DFZX1 gate177 ( .D(g6906), .TD(n3042), .SEL(test_se), .CK(clk), .Q(n3282), 
        .QB(n1932) );
  DFZX1 gate178 ( .D(g11266), .TD(n3282), .SEL(test_se), .CK(clk), .Q(n3281), 
        .QB(n1899) );
  DFZX1 gate179 ( .D(g11294), .TD(n3281), .SEL(test_se), .CK(clk), .Q(n3142)
         );
  DFZX1 gate180 ( .D(g5421), .TD(n3142), .SEL(test_se), .CK(clk), .Q(n3084) );
  DFZX1 gate181 ( .D(g8649), .TD(n3084), .SEL(test_se), .CK(clk), .Q(n3280), 
        .QB(n1905) );
  DFZX1 gate182 ( .D(g11312), .TD(n3280), .SEL(test_se), .CK(clk), .Q(n3069)
         );
  DFZX1 gate183 ( .D(g6840), .TD(n3069), .SEL(test_se), .CK(clk), .Q(n3279), 
        .QB(n2067) );
  DFZX1 gate184 ( .D(g254), .TD(n3279), .SEL(test_se), .CK(clk), .Q(n3038) );
  DFZX1 gate185 ( .D(g7202), .TD(n3038), .SEL(test_se), .CK(clk), .Q(g814), 
        .QB(n1676) );
  DFZX1 gate186 ( .D(g6834), .TD(g814), .SEL(test_se), .CK(clk), .Q(n3049) );
  DFZX1 gate187 ( .D(g10795), .TD(n3049), .SEL(test_se), .CK(clk), .Q(n3278), 
        .QB(n2019) );
  DFZX1 gate188 ( .D(g103), .TD(n3278), .SEL(test_se), .CK(clk), .Q(g2612) );
  DFZX1 gate189 ( .D(g875), .TD(g2612), .SEL(test_se), .CK(clk), .Q(n3000) );
  DFZX1 gate190 ( .D(g6831), .TD(n3000), .SEL(test_se), .CK(clk), .Q(n3277), 
        .QB(n2074) );
  DFZX1 gate191 ( .D(g8060), .TD(n3277), .SEL(test_se), .CK(clk), .Q(n2906), 
        .QB(n2008) );
  DFZX1 gate192 ( .D(g4893), .TD(n2906), .SEL(test_se), .CK(clk), .Q(n3143), 
        .QB(n2004) );
  DFZX1 gate193 ( .D(g7244), .TD(n3143), .SEL(test_se), .CK(clk), .Q(n3001) );
  DFZX1 gate194 ( .D(g6026), .TD(n3001), .SEL(test_se), .CK(clk), .Q(g259) );
  DFZX1 gate195 ( .D(g3069), .TD(g259), .SEL(test_se), .CK(clk), .Q(n3060) );
  DFZX1 gate196 ( .D(g11608), .TD(n3060), .SEL(test_se), .CK(clk), .Q(n3144)
         );
  DFZX1 gate197 ( .D(g7660), .TD(n3144), .SEL(test_se), .CK(clk), .Q(n3276), 
        .QB(n2001) );
  DFZX1 gate198 ( .D(g6911), .TD(n3276), .SEL(test_se), .CK(clk), .Q(n3087), 
        .QB(n2096) );
  DFZX1 gate199 ( .D(g11640), .TD(n3087), .SEL(test_se), .CK(clk), .Q(n3192)
         );
  DFZX1 gate200 ( .D(g8777), .TD(n3192), .SEL(test_se), .CK(clk), .Q(n3051) );
  DFZX1 gate201 ( .D(g4274), .TD(n3051), .SEL(test_se), .CK(clk), .Q(n3275), 
        .QB(n2014) );
  DFZX1 gate202 ( .D(g6215), .TD(n3275), .SEL(test_se), .CK(clk), .Q(n3145) );
  DFZX1 gate203 ( .D(g7297), .TD(n3145), .SEL(test_se), .CK(clk), .Q(n3274), 
        .QB(n1877) );
  DFZX1 gate204 ( .D(g11326), .TD(n3274), .SEL(test_se), .CK(clk), .Q(n2989), 
        .QB(n2011) );
  DFZX1 gate205 ( .D(g11269), .TD(n2989), .SEL(test_se), .CK(clk), .Q(n3037), 
        .QB(n1973) );
  DFZX1 gate206 ( .D(g11325), .TD(n3037), .SEL(test_se), .CK(clk), .Q(n3273), 
        .QB(n1918) );
  DFZX1 gate207 ( .D(g10864), .TD(n3273), .SEL(test_se), .CK(clk), .Q(n3272), 
        .QB(n2049) );
  DFZX1 gate208 ( .D(g11290), .TD(n3272), .SEL(test_se), .CK(clk), .Q(n3146)
         );
  DFZX1 gate209 ( .D(g10798), .TD(n3146), .SEL(test_se), .CK(clk), .Q(n3271), 
        .QB(n2017) );
  DFZX1 gate210 ( .D(g8284), .TD(n3271), .SEL(test_se), .CK(clk), .Q(n2896), 
        .QB(n2028) );
  DFZX1 gate211 ( .D(g11328), .TD(n2896), .SEL(test_se), .CK(clk), .Q(n2988), 
        .QB(n2026) );
  DFZX1 gate212 ( .D(g10800), .TD(n2988), .SEL(test_se), .CK(clk), .Q(n3270), 
        .QB(n2054) );
  DFZX1 gate213 ( .D(g8944), .TD(n3270), .SEL(test_se), .CK(clk), .Q(n2885) );
  DFZX1 gate214 ( .D(g7183), .TD(n2885), .SEL(test_se), .CK(clk), .Q(g8978), 
        .QB(n2038) );
  DFZX1 gate215 ( .D(g4465), .TD(g8978), .SEL(test_se), .CK(clk), .Q(n3269), 
        .QB(n1913) );
  DFZX1 gate216 ( .D(g1356), .TD(n3269), .SEL(test_se), .CK(clk), .Q(g1317) );
  DFZX1 gate217 ( .D(g11484), .TD(g1317), .SEL(test_se), .CK(clk), .Q(n2969), 
        .QB(n2087) );
  DFZX1 gate218 ( .D(g11263), .TD(n2969), .SEL(test_se), .CK(clk), .Q(n3268), 
        .QB(n1895) );
  DFZX1 gate219 ( .D(g6501), .TD(n3268), .SEL(test_se), .CK(clk), .Q(n3078), 
        .QB(n2097) );
  DFZX1 gate221 ( .D(g6757), .TD(n3078), .SEL(test_se), .CK(clk), .Q(n2903) );
  DFZX1 gate222 ( .D(g11334), .TD(n2903), .SEL(test_se), .CK(clk), .Q(n3267), 
        .QB(n1868) );
  DFZX1 gate223 ( .D(g6042), .TD(n3267), .SEL(test_se), .CK(clk), .Q(g262) );
  DFZX1 gate224 ( .D(g8384), .TD(g262), .SEL(test_se), .CK(clk), .Q(n3147), 
        .QB(n1953) );
  DFZX1 gate225 ( .D(g6653), .TD(n3147), .SEL(test_se), .CK(clk), .Q(g8983), 
        .QB(n2042) );
  DFZX1 gate226 ( .D(g257), .TD(g8983), .SEL(test_se), .CK(clk), .Q(n3033) );
  DFZX1 gate227 ( .D(n592), .TD(n3033), .SEL(test_se), .CK(clk), .Q(g1356) );
  DFZX1 gate228 ( .D(n569), .TD(g1356), .SEL(test_se), .CK(clk), .Q(g794), 
        .QB(n1812) );
  DFZX1 gate229 ( .D(n533), .TD(g794), .SEL(test_se), .CK(clk), .Q(n3266), 
        .QB(n1417) );
  DFZX1 gate230 ( .D(g6929), .TD(n3266), .SEL(test_se), .CK(clk), .Q(n3071) );
  DFZX1 gate231 ( .D(g11488), .TD(n3071), .SEL(test_se), .CK(clk), .Q(n2965), 
        .QB(n2083) );
  DFZX1 gate232 ( .D(g7299), .TD(n2965), .SEL(test_se), .CK(clk), .Q(n3265), 
        .QB(n1869) );
  DFZX1 gate233 ( .D(g4330), .TD(n3265), .SEL(test_se), .CK(clk), .Q(n3264), 
        .QB(n1949) );
  DFZX1 gate234 ( .D(g1958), .TD(n3264), .SEL(test_se), .CK(clk), .Q(n3263), 
        .QB(g8271) );
  DFZX1 gate235 ( .D(g7257), .TD(n3263), .SEL(test_se), .CK(clk), .Q(n3262), 
        .QB(n2063) );
  DFZX1 gate236 ( .D(g8775), .TD(n3262), .SEL(test_se), .CK(clk), .Q(n2920) );
  DFZX1 gate238 ( .D(g5770), .TD(n2920), .SEL(test_se), .CK(clk), .Q(n2940), 
        .QB(n1987) );
  DFZX1 gate239 ( .D(g11486), .TD(n2940), .SEL(test_se), .CK(clk), .Q(n2967), 
        .QB(n2085) );
  DFZX1 gate240 ( .D(g261), .TD(n2967), .SEL(test_se), .CK(clk), .Q(n3045) );
  DFZX1 gate241 ( .D(g4338), .TD(n3045), .SEL(test_se), .CK(clk), .Q(n3261), 
        .QB(n2072) );
  DFZX1 gate242 ( .D(g4500), .TD(n3261), .SEL(test_se), .CK(clk), .Q(n3055) );
  DFZX1 gate243 ( .D(n541), .TD(n3055), .SEL(test_se), .CK(clk), .Q(n3260), 
        .QB(n1500) );
  DFZX1 gate244 ( .D(g8147), .TD(n3260), .SEL(test_se), .CK(clk), .Q(n3259), 
        .QB(n1979) );
  DFZX1 gate245 ( .D(g6038), .TD(n3259), .SEL(test_se), .CK(clk), .Q(g261) );
  DFZX1 gate246 ( .D(g11337), .TD(g261), .SEL(test_se), .CK(clk), .Q(n3258), 
        .QB(n1894) );
  DFZX1 gate247 ( .D(g6045), .TD(n3258), .SEL(test_se), .CK(clk), .Q(g254) );
  DFZX1 gate248 ( .D(g7191), .TD(g254), .SEL(test_se), .CK(clk), .Q(g4178), 
        .QB(n1620) );
  DFZX1 gate249 ( .D(g826), .TD(g4178), .SEL(test_se), .CK(clk), .Q(n3020) );
  DFZX1 gate250 ( .D(g8774), .TD(n3020), .SEL(test_se), .CK(clk), .Q(n3048) );
  DFZX1 gate251 ( .D(g7293), .TD(n3048), .SEL(test_se), .CK(clk), .Q(n3257), 
        .QB(n1988) );
  DFZX1 gate252 ( .D(g6907), .TD(n3257), .SEL(test_se), .CK(clk), .Q(n3096) );
  DFZX1 gate253 ( .D(g4903), .TD(n3096), .SEL(test_se), .CK(clk), .Q(g1850) );
  DFZX1 gate254 ( .D(g6123), .TD(g1850), .SEL(test_se), .CK(clk), .Q(g4176), 
        .QB(n1731) );
  DFZX1 gate255 ( .D(g6506), .TD(g4176), .SEL(test_se), .CK(clk), .Q(n3256), 
        .QB(n1929) );
  DFZX1 gate256 ( .D(g11376), .TD(n3256), .SEL(test_se), .CK(clk), .Q(n3148), 
        .QB(n1892) );
  DFZX1 gate257 ( .D(g6542), .TD(n3148), .SEL(test_se), .CK(clk), .Q(n3074) );
  DFZX1 gate259 ( .D(g6551), .TD(n3074), .SEL(test_se), .CK(clk), .Q(n3112) );
  DFZX1 gate260 ( .D(g6901), .TD(n3112), .SEL(test_se), .CK(clk), .Q(n3100) );
  DFZX1 gate261 ( .D(g10797), .TD(n3100), .SEL(test_se), .CK(clk), .Q(n3255), 
        .QB(n2018) );
  DFZX1 gate262 ( .D(g8505), .TD(n3255), .SEL(test_se), .CK(clk), .Q(n3149), 
        .QB(n1968) );
  DFZX1 gate263 ( .D(g4117), .TD(n3149), .SEL(test_se), .CK(clk), .Q(g17) );
  DFZX1 gate264 ( .D(g11647), .TD(g17), .SEL(test_se), .CK(clk), .Q(n2950), 
        .QB(n2082) );
  DFZX1 gate265 ( .D(g11340), .TD(n2950), .SEL(test_se), .CK(clk), .Q(n3150), 
        .QB(n1872) );
  DFZX1 gate266 ( .D(g253), .TD(n3150), .SEL(test_se), .CK(clk), .Q(n3254), 
        .QB(n1983) );
  DFZX1 gate267 ( .D(g11625), .TD(n3254), .SEL(test_se), .CK(clk), .Q(n3253), 
        .QB(n2040) );
  DFZX1 gate268 ( .D(g636), .TD(n3253), .SEL(test_se), .CK(clk), .Q(g8) );
  DFZX1 gate269 ( .D(g6502), .TD(g8), .SEL(test_se), .CK(clk), .Q(n3151) );
  DFZX1 gate270 ( .D(n1861), .TD(n3151), .SEL(test_se), .CK(clk), .Q(g2648) );
  DFZX1 gate271 ( .D(g6049), .TD(g2648), .SEL(test_se), .CK(clk), .Q(g255) );
  DFZX1 gate272 ( .D(g8945), .TD(g255), .SEL(test_se), .CK(clk), .Q(n3152) );
  DFZX1 gate273 ( .D(g4231), .TD(n3152), .SEL(test_se), .CK(clk), .Q(n3252), 
        .QB(n2060) );
  DFZX1 gate274 ( .D(g8040), .TD(n3252), .SEL(test_se), .CK(clk), .Q(n2911) );
  DFZX1 gate276 ( .D(n681), .TD(n2911), .SEL(test_se), .CK(clk), .Q(n3251), 
        .QB(n1595) );
  DFZX1 gate277 ( .D(g6155), .TD(n3251), .SEL(test_se), .CK(clk), .Q(n3153), 
        .QB(n1870) );
  DFZX1 gate278 ( .D(g8043), .TD(n3153), .SEL(test_se), .CK(clk), .Q(n2912) );
  DFZX1 gate279 ( .D(g5173), .TD(n2912), .SEL(test_se), .CK(clk), .Q(n2952), 
        .QB(n1964) );
  DFZX1 gate280 ( .D(g6916), .TD(n2952), .SEL(test_se), .CK(clk), .Q(n3250), 
        .QB(n2058) );
  DFZX1 gate281 ( .D(g10861), .TD(n3250), .SEL(test_se), .CK(clk), .Q(n3249), 
        .QB(n1939) );
  DFZX1 gate282 ( .D(g8431), .TD(n3249), .SEL(test_se), .CK(clk), .Q(n3248), 
        .QB(n1916) );
  DFZX1 gate283 ( .D(g4309), .TD(n3248), .SEL(test_se), .CK(clk), .Q(n3116) );
  DFZX1 gate284 ( .D(g11485), .TD(n3116), .SEL(test_se), .CK(clk), .Q(n2968), 
        .QB(n2086) );
  DFZX1 gate285 ( .D(g6334), .TD(n2968), .SEL(test_se), .CK(clk), .Q(n3247), 
        .QB(n1880) );
  DFZX1 gate286 ( .D(g10767), .TD(n3247), .SEL(test_se), .CK(clk), .Q(n3246), 
        .QB(n1941) );
  DFZX1 gate287 ( .D(g8923), .TD(n3246), .SEL(test_se), .CK(clk), .Q(n2888) );
  DFZX1 gate288 ( .D(g7189), .TD(n2888), .SEL(test_se), .CK(clk), .Q(g8980), 
        .QB(n2037) );
  DFZX1 gate289 ( .D(g10799), .TD(g8980), .SEL(test_se), .CK(clk), .Q(n3245), 
        .QB(n2016) );
  DFZX1 gate290 ( .D(g6747), .TD(n3245), .SEL(test_se), .CK(clk), .Q(n3244), 
        .QB(n2031) );
  DFZX1 gate291 ( .D(g6080), .TD(n3244), .SEL(test_se), .CK(clk), .Q(n2933) );
  DFZX1 gate292 ( .D(g3381), .TD(n2933), .SEL(test_se), .CK(clk), .Q(g2986) );
  DFZX1 gate293 ( .D(g5910), .TD(g2986), .SEL(test_se), .CK(clk), .Q(n2938) );
  DFZX1 gate294 ( .D(g11393), .TD(n2938), .SEL(test_se), .CK(clk), .Q(n3082)
         );
  DFZX1 gate295 ( .D(g11349), .TD(n3082), .SEL(test_se), .CK(clk), .Q(n3107)
         );
  DFZX1 gate296 ( .D(g83), .TD(n3107), .SEL(test_se), .CK(clk), .Q(g1955) );
  DFZX1 gate297 ( .D(g6439), .TD(g1955), .SEL(test_se), .CK(clk), .Q(n2925), 
        .QB(n1911) );
  DFZX1 gate298 ( .D(g9266), .TD(n2925), .SEL(test_se), .CK(clk), .Q(n3188), 
        .QB(n1871) );
  DFZX1 gate300 ( .D(g1217), .TD(n3188), .SEL(test_se), .CK(clk), .Q(n2951) );
  DFZX1 gate301 ( .D(g8940), .TD(n2951), .SEL(test_se), .CK(clk), .Q(n3154) );
  DFZX1 gate302 ( .D(g7705), .TD(n3154), .SEL(test_se), .CK(clk), .Q(g4179), 
        .QB(n1688) );
  DFZX1 gate303 ( .D(g9269), .TD(g4179), .SEL(test_se), .CK(clk), .Q(n3155), 
        .QB(n1890) );
  DFZX1 gate304 ( .D(g6820), .TD(n3155), .SEL(test_se), .CK(clk), .Q(n3054) );
  DFZX1 gate305 ( .D(g756), .TD(n3054), .SEL(test_se), .CK(clk), .Q(g746), 
        .QB(n1794) );
  DFZX1 gate307 ( .D(g8042), .TD(g746), .SEL(test_se), .CK(clk), .Q(n3243), 
        .QB(n1986) );
  DFZX1 gate308 ( .D(g6759), .TD(n3243), .SEL(test_se), .CK(clk), .Q(n2910) );
  DFZX1 gate309 ( .D(g11487), .TD(n2910), .SEL(test_se), .CK(clk), .Q(n2966), 
        .QB(n2084) );
  DFZX1 gate310 ( .D(g802), .TD(n2966), .SEL(test_se), .CK(clk), .Q(n3023) );
  DFZX1 gate311 ( .D(g9124), .TD(n3023), .SEL(test_se), .CK(clk), .Q(n3156), 
        .QB(n1954) );
  DFZX1 gate312 ( .D(g11293), .TD(n3156), .SEL(test_se), .CK(clk), .Q(g1854), 
        .QB(n2998) );
  DFZX1 gate313 ( .D(g11298), .TD(g1854), .SEL(test_se), .CK(clk), .Q(n3118)
         );
  DFZX1 gate314 ( .D(g8287), .TD(n3118), .SEL(test_se), .CK(clk), .Q(n3157), 
        .QB(n1923) );
  DFZX1 gate315 ( .D(g8047), .TD(n3157), .SEL(test_se), .CK(clk), .Q(n2901) );
  DFZX1 gate316 ( .D(g6205), .TD(n2901), .SEL(test_se), .CK(clk), .Q(n2926), 
        .QB(n2065) );
  DFZX1 gate317 ( .D(g8885), .TD(n2926), .SEL(test_se), .CK(clk), .Q(n3158) );
  DFZX1 gate318 ( .D(g11305), .TD(n3158), .SEL(test_se), .CK(clk), .Q(n3093)
         );
  DFZX1 gate319 ( .D(g5556), .TD(n3093), .SEL(test_se), .CK(clk), .Q(g1958) );
  DFZX1 gate320 ( .D(n578), .TD(g1958), .SEL(test_se), .CK(clk), .Q(n2098) );
  DFZX1 gate321 ( .D(g2478), .TD(n2098), .SEL(test_se), .CK(clk), .Q(g1765) );
  DFZX1 gate322 ( .D(g10711), .TD(g1765), .SEL(test_se), .CK(clk), .Q(n3242), 
        .QB(n2071) );
  DFZX1 gate323 ( .D(g7303), .TD(n3242), .SEL(test_se), .CK(clk), .Q(n2985), 
        .QB(n1978) );
  DFZX1 gate324 ( .D(g5194), .TD(n2985), .SEL(test_se), .CK(clk), .Q(n3159) );
  DFZX1 gate325 ( .D(g7541), .TD(n3159), .SEL(test_se), .CK(clk), .Q(n3186) );
  DFZX1 gate326 ( .D(g11607), .TD(n3186), .SEL(test_se), .CK(clk), .Q(n3081)
         );
  DFZX1 gate327 ( .D(g6541), .TD(n3081), .SEL(test_se), .CK(clk), .Q(n3241), 
        .QB(n2056) );
  DFZX1 gate328 ( .D(g6827), .TD(n3241), .SEL(test_se), .CK(clk), .Q(n2943) );
  DFZX1 gate329 ( .D(g4114), .TD(n2943), .SEL(test_se), .CK(clk), .Q(g3069), 
        .QB(n3061) );
  DFZX1 gate330 ( .D(g11332), .TD(g3069), .SEL(test_se), .CK(clk), .Q(n3240), 
        .QB(n1898) );
  DFZX1 gate331 ( .D(g4902), .TD(n3240), .SEL(test_se), .CK(clk), .Q(n3239), 
        .QB(n1405) );
  DFZX1 gate332 ( .D(g6828), .TD(n3239), .SEL(test_se), .CK(clk), .Q(n3018), 
        .QB(n2078) );
  DFZX1 gate333 ( .D(g6516), .TD(n3018), .SEL(test_se), .CK(clk), .Q(n3160), 
        .QB(n1992) );
  DFZX1 gate334 ( .D(g8938), .TD(n3160), .SEL(test_se), .CK(clk), .Q(n3161), 
        .QB(n1972) );
  DFZX1 gate335 ( .D(g7298), .TD(n3161), .SEL(test_se), .CK(clk), .Q(n2982), 
        .QB(n1977) );
  DFZX1 gate336 ( .D(n519), .TD(n2982), .SEL(test_se), .CK(clk), .Q(n2080), 
        .QB(n3058) );
  DFZX1 gate337 ( .D(g6672), .TD(n2080), .SEL(test_se), .CK(clk), .Q(n3238), 
        .QB(n1434) );
  DFZX1 gate338 ( .D(g8048), .TD(n3238), .SEL(test_se), .CK(clk), .Q(n2922), 
        .QB(n1981) );
  DFZX1 gate339 ( .D(g798), .TD(n2922), .SEL(test_se), .CK(clk), .Q(n3025) );
  DFZX1 gate340 ( .D(g8285), .TD(n3025), .SEL(test_se), .CK(clk), .Q(n2895), 
        .QB(n1928) );
  DFZX1 gate341 ( .D(g8254), .TD(n2895), .SEL(test_se), .CK(clk), .Q(n3162) );
  DFZX1 gate343 ( .D(g11604), .TD(n3162), .SEL(test_se), .CK(clk), .Q(n3237), 
        .QB(n1948) );
  DFZX1 gate344 ( .D(g814), .TD(n3237), .SEL(test_se), .CK(clk), .Q(n3026) );
  DFZX1 gate345 ( .D(g11636), .TD(n3026), .SEL(test_se), .CK(clk), .Q(n3163), 
        .QB(n2000) );
  DFZX1 gate346 ( .D(g6910), .TD(n3163), .SEL(test_se), .CK(clk), .Q(n3236), 
        .QB(n1931) );
  DFZX1 gate347 ( .D(g8173), .TD(n3236), .SEL(test_se), .CK(clk), .Q(n2997), 
        .QB(n1993) );
  DFZX1 gate348 ( .D(g8245), .TD(n2997), .SEL(test_se), .CK(clk), .Q(g826), 
        .QB(n1674) );
  DFZX1 gate350 ( .D(g8281), .TD(g826), .SEL(test_se), .CK(clk), .Q(n3164), 
        .QB(n1906) );
  DFZX1 gate351 ( .D(n546), .TD(n3164), .SEL(test_se), .CK(clk), .Q(n3235), 
        .QB(n1448) );
  DFZX1 gate352 ( .D(g11314), .TD(n3235), .SEL(test_se), .CK(clk), .Q(n3117)
         );
  DFZX1 gate353 ( .D(g4905), .TD(n3117), .SEL(test_se), .CK(clk), .Q(n3234), 
        .QB(n1970) );
  DFZX1 gate354 ( .D(g4484), .TD(n3234), .SEL(test_se), .CK(clk), .Q(n3233), 
        .QB(n1908) );
  DFZX1 gate355 ( .D(g8937), .TD(n3233), .SEL(test_se), .CK(clk), .Q(n3183) );
  DFZX1 gate356 ( .D(g7300), .TD(n3183), .SEL(test_se), .CK(clk), .Q(n2986), 
        .QB(n1980) );
  DFZX1 gate357 ( .D(g6002), .TD(n2986), .SEL(test_se), .CK(clk), .Q(g257) );
  DFZX1 gate358 ( .D(n1865), .TD(g257), .SEL(test_se), .CK(clk), .Q(g874) );
  DFZX1 gate359 ( .D(g9110), .TD(g874), .SEL(test_se), .CK(clk), .Q(n3165), 
        .QB(n1889) );
  DFZX1 gate360 ( .D(g8926), .TD(n3165), .SEL(test_se), .CK(clk), .Q(n3166) );
  DFZX1 gate361 ( .D(g8631), .TD(n3166), .SEL(test_se), .CK(clk), .Q(g636), 
        .QB(n2892) );
  DFZX1 gate362 ( .D(g7632), .TD(g636), .SEL(test_se), .CK(clk), .Q(n2978) );
  DFZX1 gate363 ( .D(g9150), .TD(n2978), .SEL(test_se), .CK(clk), .Q(n2948) );
  DFZX1 gate364 ( .D(g6531), .TD(n2948), .SEL(test_se), .CK(clk), .Q(g8986), 
        .QB(n2046) );
  DFZX1 gate365 ( .D(g6786), .TD(g8986), .SEL(test_se), .CK(clk), .Q(n2923), 
        .QB(n2073) );
  DFZX1 gate366 ( .D(g11303), .TD(n2923), .SEL(test_se), .CK(clk), .Q(n3106)
         );
  DFZX1 gate367 ( .D(g4477), .TD(n3106), .SEL(test_se), .CK(clk), .Q(n2960), 
        .QB(n1884) );
  DFZX1 gate368 ( .D(g822), .TD(n2960), .SEL(test_se), .CK(clk), .Q(n3024) );
  DFZX1 gate369 ( .D(g11258), .TD(n3024), .SEL(test_se), .CK(clk), .Q(n3032), 
        .QB(n2012) );
  DFZX1 gate370 ( .D(g9272), .TD(n3032), .SEL(test_se), .CK(clk), .Q(n3189), 
        .QB(n1961) );
  DFZX1 gate371 ( .D(g10773), .TD(n3189), .SEL(test_se), .CK(clk), .Q(n3232), 
        .QB(n2068) );
  DFZX1 gate372 ( .D(g6470), .TD(n3232), .SEL(test_se), .CK(clk), .Q(n3104) );
  DFZX1 gate373 ( .D(g5083), .TD(n3104), .SEL(test_se), .CK(clk), .Q(n3057) );
  DFZX1 gate374 ( .D(g8286), .TD(n3057), .SEL(test_se), .CK(clk), .Q(n3231), 
        .QB(n1989) );
  DFZX1 gate375 ( .D(g8773), .TD(n3231), .SEL(test_se), .CK(clk), .Q(n3013) );
  DFZX1 gate377 ( .D(g6054), .TD(n3013), .SEL(test_se), .CK(clk), .Q(n2937) );
  DFZX1 gate378 ( .D(g101), .TD(n2937), .SEL(test_se), .CK(clk), .Q(g2601) );
  DFZX1 gate379 ( .D(g11260), .TD(g2601), .SEL(test_se), .CK(clk), .Q(n3230), 
        .QB(n1991) );
  DFZX1 gate380 ( .D(g11338), .TD(n3230), .SEL(test_se), .CK(clk), .Q(n2990), 
        .QB(n1975) );
  DFZX1 gate381 ( .D(g5918), .TD(n2990), .SEL(test_se), .CK(clk), .Q(n3167), 
        .QB(n1997) );
  DFZX1 gate382 ( .D(g8922), .TD(n3167), .SEL(test_se), .CK(clk), .Q(n3168) );
  DFZX1 gate383 ( .D(g8049), .TD(n3168), .SEL(test_se), .CK(clk), .Q(n2905), 
        .QB(n1934) );
  DFZX1 gate384 ( .D(g4342), .TD(n2905), .SEL(test_se), .CK(clk), .Q(n3169) );
  DFZX1 gate385 ( .D(n540), .TD(n3169), .SEL(test_se), .CK(clk), .Q(n3229), 
        .QB(n3094) );
  DFZX1 gate386 ( .D(g6755), .TD(n3229), .SEL(test_se), .CK(clk), .Q(n3228), 
        .QB(n1549) );
  DFZX1 gate387 ( .D(g6897), .TD(n3228), .SEL(test_se), .CK(clk), .Q(n3099) );
  DFZX1 gate388 ( .D(g7709), .TD(n3099), .SEL(test_se), .CK(clk), .Q(g818), 
        .QB(n1738) );
  DFZX1 gate389 ( .D(g4255), .TD(g818), .SEL(test_se), .CK(clk), .Q(n3227), 
        .QB(n1947) );
  DFZX1 gate390 ( .D(g5543), .TD(n3227), .SEL(test_se), .CK(clk), .Q(g802), 
        .QB(n1727) );
  DFZX1 gate391 ( .D(g6915), .TD(g802), .SEL(test_se), .CK(clk), .Q(n3226), 
        .QB(n1945) );
  DFZX1 gate392 ( .D(g6513), .TD(n3226), .SEL(test_se), .CK(clk), .Q(n3098) );
  DFZX1 gate393 ( .D(g6480), .TD(n3098), .SEL(test_se), .CK(clk), .Q(n3080) );
  DFZX1 gate394 ( .D(g6733), .TD(n3080), .SEL(test_se), .CK(clk), .Q(g810), 
        .QB(n1672) );
  DFZX1 gate395 ( .D(g11264), .TD(g810), .SEL(test_se), .CK(clk), .Q(n3036), 
        .QB(n1995) );
  DFZX1 gate396 ( .D(g8973), .TD(n3036), .SEL(test_se), .CK(clk), .Q(n3170) );
  DFZX1 gate397 ( .D(g6833), .TD(n3170), .SEL(test_se), .CK(clk), .Q(n2942) );
  DFZX1 gate398 ( .D(g5996), .TD(n2942), .SEL(test_se), .CK(clk), .Q(g253) );
  DFZX1 gate399 ( .D(n1866), .TD(g253), .SEL(test_se), .CK(clk), .Q(g875) );
  DFZX1 gate400 ( .D(g4473), .TD(g875), .SEL(test_se), .CK(clk), .Q(n2959), 
        .QB(n2013) );
  DFZX1 gate401 ( .D(g5755), .TD(n2959), .SEL(test_se), .CK(clk), .Q(n3171), 
        .QB(n1999) );
  DFZX1 gate402 ( .D(g7295), .TD(n3171), .SEL(test_se), .CK(clk), .Q(n2979), 
        .QB(n2093) );
  DFZX1 gate403 ( .D(g6068), .TD(n2979), .SEL(test_se), .CK(clk), .Q(n2935) );
  DFZX1 gate404 ( .D(g7137), .TD(n2935), .SEL(test_se), .CK(clk), .Q(n2899) );
  DFZX1 gate405 ( .D(g8779), .TD(n2899), .SEL(test_se), .CK(clk), .Q(n3011) );
  DFZX1 gate406 ( .D(g818), .TD(n3011), .SEL(test_se), .CK(clk), .Q(n3028) );
  DFZX1 gate407 ( .D(g11270), .TD(n3028), .SEL(test_se), .CK(clk), .Q(n3039), 
        .QB(n1881) );
  DFZX1 gate408 ( .D(g5529), .TD(n3039), .SEL(test_se), .CK(clk), .Q(g4174), 
        .QB(n1742) );
  DFZX1 gate409 ( .D(g11306), .TD(g4174), .SEL(test_se), .CK(clk), .Q(n3172)
         );
  DFZX1 gate410 ( .D(g11291), .TD(n3172), .SEL(test_se), .CK(clk), .Q(n3173)
         );
  DFZX1 gate411 ( .D(g4283), .TD(n3173), .SEL(test_se), .CK(clk), .Q(n3077) );
  DFZX1 gate412 ( .D(g29), .TD(n3077), .SEL(test_se), .CK(clk), .Q(g2604) );
  DFZX1 gate413 ( .D(g806), .TD(g2604), .SEL(test_se), .CK(clk), .Q(n3022) );
  DFZX1 gate414 ( .D(g6894), .TD(n3022), .SEL(test_se), .CK(clk), .Q(n3002) );
  DFZX1 gate415 ( .D(g6902), .TD(n3002), .SEL(test_se), .CK(clk), .Q(n3009) );
  DFZX1 gate416 ( .D(g8765), .TD(n3009), .SEL(test_se), .CK(clk), .Q(n2921) );
  DFZX1 gate417 ( .D(g4498), .TD(n2921), .SEL(test_se), .CK(clk), .Q(n2958), 
        .QB(n1924) );
  DFZX1 gate418 ( .D(g5148), .TD(n2958), .SEL(test_se), .CK(clk), .Q(n2953), 
        .QB(n1966) );
  DFZX1 gate419 ( .D(g7581), .TD(n2953), .SEL(test_se), .CK(clk), .Q(n2975), 
        .QB(n1994) );
  DFZX1 gate420 ( .D(g11267), .TD(n2975), .SEL(test_se), .CK(clk), .Q(n3044), 
        .QB(n1976) );
  DFZX1 gate421 ( .D(g10936), .TD(n3044), .SEL(test_se), .CK(clk), .Q(n3225), 
        .QB(n2062) );
  DFZX1 gate422 ( .D(g10784), .TD(n3225), .SEL(test_se), .CK(clk), .Q(n3047)
         );
  DFZX1 gate424 ( .D(g10765), .TD(n3047), .SEL(test_se), .CK(clk), .Q(n3224), 
        .QB(n1942) );
  DFZX1 gate425 ( .D(g6332), .TD(n3224), .SEL(test_se), .CK(clk), .Q(n3223), 
        .QB(n1984) );
  DFZX1 gate426 ( .D(g6479), .TD(n3223), .SEL(test_se), .CK(clk), .Q(n3089), 
        .QB(n2079) );
  DFZX1 gate427 ( .D(g6537), .TD(n3089), .SEL(test_se), .CK(clk), .Q(n3072) );
  DFZX1 gate428 ( .D(g8434), .TD(n3072), .SEL(test_se), .CK(clk), .Q(n3174), 
        .QB(n1922) );
  DFZX1 gate429 ( .D(g6908), .TD(n3174), .SEL(test_se), .CK(clk), .Q(n3004) );
  DFZX1 gate430 ( .D(g6243), .TD(n3004), .SEL(test_se), .CK(clk), .Q(g798), 
        .QB(n1651) );
  DFZX1 gate431 ( .D(g11324), .TD(g798), .SEL(test_se), .CK(clk), .Q(n3222), 
        .QB(n1897) );
  DFZX1 gate432 ( .D(g3462), .TD(n3222), .SEL(test_se), .CK(clk), .Q(g4172), 
        .QB(n1768) );
  DFZX1 gate433 ( .D(g11609), .TD(g4172), .SEL(test_se), .CK(clk), .Q(n3175)
         );
  DFZX1 gate434 ( .D(g810), .TD(n3175), .SEL(test_se), .CK(clk), .Q(n3021) );
  DFZX1 gate435 ( .D(g8244), .TD(n3021), .SEL(test_se), .CK(clk), .Q(g4181), 
        .QB(n1743) );
  DFZX1 gate436 ( .D(g8194), .TD(g4181), .SEL(test_se), .CK(clk), .Q(n3221), 
        .QB(n2041) );
  DFZX1 gate437 ( .D(g113), .TD(n3221), .SEL(test_se), .CK(clk), .Q(g114) );
  DFZX1 gate438 ( .D(g8052), .TD(g114), .SEL(test_se), .CK(clk), .Q(n2914) );
  DFZX1 gate439 ( .D(g4325), .TD(n2914), .SEL(test_se), .CK(clk), .Q(n2954) );
  DFZX1 gate441 ( .D(g11481), .TD(n2954), .SEL(test_se), .CK(clk), .Q(n2972), 
        .QB(n2090) );
  DFZX1 gate442 ( .D(g874), .TD(n2972), .SEL(test_se), .CK(clk), .Q(n3220), 
        .QB(n1594) );
  DFZX1 gate443 ( .D(g7301), .TD(n3220), .SEL(test_se), .CK(clk), .Q(n2984), 
        .QB(n1903) );
  DFZX1 gate444 ( .D(g6035), .TD(n2984), .SEL(test_se), .CK(clk), .Q(g260) );
  DFZX1 gate445 ( .D(g8059), .TD(g260), .SEL(test_se), .CK(clk), .Q(n2908) );
  DFZX1 gate446 ( .D(g1854), .TD(n2908), .SEL(test_se), .CK(clk), .Q(n3219), 
        .QB(n3076) );
  DFZX1 gate447 ( .D(g6015), .TD(n3219), .SEL(test_se), .CK(clk), .Q(g258) );
  DFZX1 gate448 ( .D(g11330), .TD(g258), .SEL(test_se), .CK(clk), .Q(n3176) );
  DFZX1 gate449 ( .D(g11605), .TD(n3176), .SEL(test_se), .CK(clk), .Q(n3193)
         );
  DFZX1 gate450 ( .D(g8921), .TD(n3193), .SEL(test_se), .CK(clk), .Q(n3177), 
        .QB(n1967) );
  DFZX1 gate451 ( .D(g8883), .TD(n3177), .SEL(test_se), .CK(clk), .Q(n2890) );
  DFZX1 gate452 ( .D(g28), .TD(n2890), .SEL(test_se), .CK(clk), .Q(g2608) );
  DFZX1 gate453 ( .D(g6163), .TD(g2608), .SEL(test_se), .CK(clk), .Q(n3218), 
        .QB(n1584) );
  DFZX1 gate454 ( .D(g6523), .TD(n3218), .SEL(test_se), .CK(clk), .Q(n3102) );
  DFZX1 gate455 ( .D(g11300), .TD(n3102), .SEL(test_se), .CK(clk), .Q(n3108)
         );
  DFZX1 gate456 ( .D(g9555), .TD(n3108), .SEL(test_se), .CK(clk), .Q(n2999), 
        .QB(n1962) );
  DFZX1 gate457 ( .D(g6481), .TD(n2999), .SEL(test_se), .CK(clk), .Q(n3217), 
        .QB(n1946) );
  DFZX1 gate458 ( .D(g4471), .TD(n3217), .SEL(test_se), .CK(clk), .Q(n3216), 
        .QB(n1982) );
  DFZX1 gate459 ( .D(g11606), .TD(n3216), .SEL(test_se), .CK(clk), .Q(n3088)
         );
  DFZX1 gate460 ( .D(g11335), .TD(n3088), .SEL(test_se), .CK(clk), .Q(n3215), 
        .QB(n1960) );
  DFZX1 gate461 ( .D(g10791), .TD(n3215), .SEL(test_se), .CK(clk), .Q(n3214), 
        .QB(n2022) );
  DFZX1 gate462 ( .D(g8939), .TD(n3214), .SEL(test_se), .CK(clk), .Q(n2887) );
  DFZX1 gate463 ( .D(g83), .TD(n2887), .SEL(test_se), .CK(clk), .Q(g755) );
  DFZX1 gate464 ( .D(g6529), .TD(g755), .SEL(test_se), .CK(clk), .Q(n3213), 
        .QB(n2059) );
  DFZX1 gate465 ( .D(g101), .TD(n3213), .SEL(test_se), .CK(clk), .Q(g2610) );
  DFZX1 gate466 ( .D(g10776), .TD(g2610), .SEL(test_se), .CK(clk), .Q(n3212), 
        .QB(n2055) );
  DFZX1 gate467 ( .D(g6514), .TD(n3212), .SEL(test_se), .CK(clk), .Q(n3114) );
  DFZX1 gate468 ( .D(g259), .TD(n3114), .SEL(test_se), .CK(clk), .Q(n3034) );
  DFZX1 gate469 ( .D(g4490), .TD(n3034), .SEL(test_se), .CK(clk), .Q(n2957), 
        .QB(n2076) );
  DFZX1 gate471 ( .D(g11639), .TD(n2957), .SEL(test_se), .CK(clk), .Q(n3178)
         );
  DFZX1 gate472 ( .D(g4089), .TD(n3178), .SEL(test_se), .CK(clk), .Q(n3211), 
        .QB(n1426) );
  DFZX1 gate473 ( .D(g10785), .TD(n3211), .SEL(test_se), .CK(clk), .Q(n3046)
         );
  DFZX1 gate474 ( .D(g6179), .TD(n3046), .SEL(test_se), .CK(clk), .Q(n3179) );
  DFZX1 gate475 ( .D(g8053), .TD(n3179), .SEL(test_se), .CK(clk), .Q(n2907) );
  DFZX1 gate476 ( .D(g11329), .TD(n2907), .SEL(test_se), .CK(clk), .Q(n3185)
         );
  DFZX1 gate477 ( .D(g104), .TD(n3185), .SEL(test_se), .CK(clk), .Q(g2607) );
  DFZX1 gate478 ( .D(g6515), .TD(g2607), .SEL(test_se), .CK(clk), .Q(n3067) );
  DFZX1 gate479 ( .D(g258), .TD(n3067), .SEL(test_se), .CK(clk), .Q(n3035) );
  DFZX1 gate480 ( .D(g7204), .TD(n3035), .SEL(test_se), .CK(clk), .Q(g8982), 
        .QB(n2036) );
  DFZX1 gate481 ( .D(g11443), .TD(g8982), .SEL(test_se), .CK(clk), .Q(n3210), 
        .QB(n1896) );
  DFZX1 gate482 ( .D(g11603), .TD(n3210), .SEL(test_se), .CK(clk), .Q(n3180)
         );
  DFZX1 gate483 ( .D(g8770), .TD(n3180), .SEL(test_se), .CK(clk), .Q(n3017) );
  DFZX1 gate484 ( .D(g11292), .TD(n3017), .SEL(test_se), .CK(clk), .Q(n3209), 
        .QB(n2066) );
  DFZX1 gate485 ( .D(g6331), .TD(n3209), .SEL(test_se), .CK(clk), .Q(n2946) );
  DFZX1 gate486 ( .D(g6900), .TD(n2946), .SEL(test_se), .CK(clk), .Q(n3097) );
  DFZX1 gate487 ( .D(g7294), .TD(n3097), .SEL(test_se), .CK(clk), .Q(n3208), 
        .QB(n1900) );
  DFZX1 gate488 ( .D(g6829), .TD(n3208), .SEL(test_se), .CK(clk), .Q(n2944) );
  DFZX1 gate489 ( .D(g8428), .TD(n2944), .SEL(test_se), .CK(clk), .Q(n3181), 
        .QB(n2030) );
  DFZX1 gate490 ( .D(g4904), .TD(n3181), .SEL(test_se), .CK(clk), .Q(n3207), 
        .QB(n1576) );
  DFZX1 gate491 ( .D(g8054), .TD(n3207), .SEL(test_se), .CK(clk), .Q(n2904) );
  DFZX1 gate492 ( .D(g11268), .TD(n2904), .SEL(test_se), .CK(clk), .Q(n3041), 
        .QB(n1902) );
  DFZX1 gate493 ( .D(g11262), .TD(n3041), .SEL(test_se), .CK(clk), .Q(n3206), 
        .QB(n1990) );
  DFZX1 gate494 ( .D(g8283), .TD(n3206), .SEL(test_se), .CK(clk), .Q(n3205), 
        .QB(n1912) );
  DFZX1 gate495 ( .D(g6193), .TD(n3205), .SEL(test_se), .CK(clk), .Q(n2963), 
        .QB(n1917) );
  DFZX1 gate496 ( .D(g8776), .TD(n2963), .SEL(test_se), .CK(clk), .Q(n3053) );
  DFZX1 gate497 ( .D(g7143), .TD(n3053), .SEL(test_se), .CK(clk), .Q(g8976), 
        .QB(n2039) );
  DFZX1 gate498 ( .D(g6898), .TD(g8976), .SEL(test_se), .CK(clk), .Q(n3010) );
  DFZX1 gate499 ( .D(g7291), .TD(n3010), .SEL(test_se), .CK(clk), .Q(n2981), 
        .QB(n2007) );
  DFZX1 gate500 ( .D(g11478), .TD(n2981), .SEL(test_se), .CK(clk), .Q(n2973), 
        .QB(n2091) );
  DFZX1 gate501 ( .D(g6000), .TD(n2973), .SEL(test_se), .CK(clk), .Q(g256) );
  DFZX1 gate502 ( .D(g4264), .TD(g256), .SEL(test_se), .CK(clk), .Q(n3204), 
        .QB(n2015) );
  DFZX1 gate503 ( .D(g102), .TD(n3204), .SEL(test_se), .CK(clk), .Q(g2611) );
  DFZX1 gate504 ( .D(g8768), .TD(g2611), .SEL(test_se), .CK(clk), .Q(n2918) );
  DFZX1 gate505 ( .D(g10863), .TD(n2918), .SEL(test_se), .CK(clk), .Q(n3203), 
        .QB(n1938) );
  DFZX1 gate506 ( .D(g6522), .TD(n3203), .SEL(test_se), .CK(clk), .Q(n3182) );
  DFZX1 gate507 ( .D(g11641), .TD(n3182), .SEL(test_se), .CK(clk), .Q(n3190)
         );
  DFZX1 gate508 ( .D(g10780), .TD(n3190), .SEL(test_se), .CK(clk), .Q(n3202), 
        .QB(n2075) );
  DFZX1 gate509 ( .D(g8044), .TD(n3202), .SEL(test_se), .CK(clk), .Q(n2909) );
  DFZX1 gate510 ( .D(g11579), .TD(n2909), .SEL(test_se), .CK(clk), .Q(n3201), 
        .QB(n2023) );
  DFZX1 gate511 ( .D(g7296), .TD(n3201), .SEL(test_se), .CK(clk), .Q(n2983), 
        .QB(n1998) );
  DFZX1 gate512 ( .D(g6923), .TD(n2983), .SEL(test_se), .CK(clk), .Q(n3073) );
  DFZX1 gate513 ( .D(g11261), .TD(n3073), .SEL(test_se), .CK(clk), .Q(n3200), 
        .QB(n1904) );
  DFZX1 gate514 ( .D(g6638), .TD(n3200), .SEL(test_se), .CK(clk), .Q(g8981), 
        .QB(n2043) );
  DFZX1 gate515 ( .D(g6534), .TD(g8981), .SEL(test_se), .CK(clk), .Q(n3199), 
        .QB(n1887) );
  DFZX1 gate516 ( .D(g6895), .TD(n3199), .SEL(test_se), .CK(clk), .Q(n3003) );
  DFZX1 gate517 ( .D(g8771), .TD(n3003), .SEL(test_se), .CK(clk), .Q(n3015) );
  DFZX1 gate518 ( .D(g4506), .TD(n3015), .SEL(test_se), .CK(clk), .Q(n2956), 
        .QB(n2033) );
  DFZX1 gate519 ( .D(g7441), .TD(n2956), .SEL(test_se), .CK(clk), .Q(n2900) );
  DFZX1 gate520 ( .D(g8055), .TD(n2900), .SEL(test_se), .CK(clk), .Q(n2941) );
  DFZX1 gate521 ( .D(g6468), .TD(n2941), .SEL(test_se), .CK(clk), .Q(n3101) );
  DFZX1 gate522 ( .D(g8430), .TD(n3101), .SEL(test_se), .CK(clk), .Q(n2894), 
        .QB(n2027) );
  DFZX1 gate523 ( .D(g11327), .TD(n2894), .SEL(test_se), .CK(clk), .Q(n2987), 
        .QB(n1925) );
  DFZX1 gate524 ( .D(g6508), .TD(n2987), .SEL(test_se), .CK(clk), .Q(n2994), 
        .QB(n1956) );
  DFZX1 gate525 ( .D(g10717), .TD(n2994), .SEL(test_se), .CK(clk), .Q(n3198), 
        .QB(n2024) );
  DFZX1 gate526 ( .D(g4334), .TD(n3198), .SEL(test_se), .CK(clk), .Q(n2955) );
  DFZX1 gate527 ( .D(n1864), .TD(n2955), .SEL(test_se), .CK(clk), .Q(g1360) );
  DFZX1 gate529 ( .D(g6679), .TD(g1360), .SEL(test_se), .CK(clk), .Q(n3191), 
        .QB(n2099) );
  DFZX1 gate530 ( .D(g11336), .TD(n3191), .SEL(test_se), .CK(clk), .Q(n3197), 
        .QB(n1876) );
  DFZX1 gate531 ( .D(g10771), .TD(n3197), .SEL(test_se), .CK(clk), .Q(n3196), 
        .QB(n1935) );
  DFZX1 gate532 ( .D(g5445), .TD(n3196), .SEL(test_se), .CK(clk), .Q(n3091), 
        .QB(n1996) );
  DFZX1 gate533 ( .D(g8559), .TD(n3091), .SEL(test_se), .CK(clk), .Q(n2898), 
        .QB(n2003) );
  DFZX1 gate534 ( .D(g7219), .TD(n2898), .SEL(test_se), .CK(clk), .Q(g8984), 
        .QB(n2035) );
  AN3X1 U1365 ( .I1(n2451), .I2(n1591), .I3(g109), .O(n2455) );
  INVX2 U1366 ( .I(g109), .O(n2295) );
  NR2X2 U1367 ( .I1(n3057), .I2(g1696), .O(n2292) );
  TIE0X1 U1368 ( .O(g11489) );
  TIE1X1 U1369 ( .O(n1591) );
  AOI12X1 U1370 ( .B1(g881), .B2(g109), .A1(n2102), .O(n577) );
  INVCKX1 U1371 ( .I(n2103), .O(n569) );
  ND3X1 U1372 ( .I1(g47), .I2(n2104), .I3(n2105), .O(n1867) );
  OR4B2XLP U1373 ( .I1(n2106), .I2(g47), .B1(n2105), .B2(n2107), .O(n1866) );
  ND3X1 U1374 ( .I1(g46), .I2(n2108), .I3(n2109), .O(n1865) );
  ND3X1 U1375 ( .I1(g47), .I2(n2106), .I3(n2109), .O(n1864) );
  AN3X1 U1376 ( .I1(n2107), .I2(n2110), .I3(n2111), .O(n2109) );
  XOR2X1 U1377 ( .I1(n2947), .I2(n2112), .O(n1861) );
  NR2X1 U1378 ( .I1(n1743), .I2(n2113), .O(n2112) );
  OR3B1XLP U1379 ( .I1(g31), .I2(g30), .B1(n2107), .O(g9961) );
  NR2X1 U1380 ( .I1(n2114), .I2(n2115), .O(g9721) );
  XNR2X1 U1381 ( .I1(n3136), .I2(n2116), .O(n2114) );
  NR2X1 U1382 ( .I1(n2117), .I2(n2118), .O(n2116) );
  AOI112X1 U1383 ( .C1(n2119), .C2(n2120), .A1(n3149), .B1(n2121), .O(n2117)
         );
  MUXB2X1 U1384 ( .EB(n2115), .A(n2122), .B(n2123), .S(n2999), .O(g9555) );
  ND2X1 U1385 ( .I1(n2124), .I2(n2125), .O(n2123) );
  OAI12X1 U1386 ( .B1(n2126), .B2(n1871), .A1(n1953), .O(n2125) );
  NR2X1 U1387 ( .I1(n2127), .I2(n1953), .O(n2122) );
  NR2X1 U1388 ( .I1(n2128), .I2(n2115), .O(g9272) );
  XNR2X1 U1389 ( .I1(n3189), .I2(n2129), .O(n2128) );
  AOI13X1 U1390 ( .B1(n2130), .B2(n2131), .B3(n2132), .A1(n2133), .O(n2129) );
  MXL2XLP U1391 ( .A(n2134), .B(n2135), .S(n1961), .OB(n2132) );
  NR2X1 U1392 ( .I1(n1871), .I2(n1890), .O(n2134) );
  NR2X1 U1393 ( .I1(n2136), .I2(n2115), .O(g9269) );
  XNR2X1 U1394 ( .I1(n2137), .I2(n1890), .O(n2136) );
  OAI13X1 U1395 ( .B1(n2138), .B2(n2139), .B3(n2140), .A1(n2126), .O(n2137) );
  NR2X1 U1396 ( .I1(n2141), .I2(n2115), .O(g9266) );
  XNR2X1 U1397 ( .I1(n2142), .I2(n1871), .O(n2141) );
  OAI13X1 U1398 ( .B1(n2140), .B2(n2135), .B3(n2143), .A1(n2126), .O(n2142) );
  INVCKX1 U1399 ( .I(n2144), .O(n2143) );
  NR2X1 U1400 ( .I1(n2145), .I2(n3155), .O(n2140) );
  NR2X1 U1401 ( .I1(n2115), .I2(n2146), .O(g9150) );
  XOR2X1 U1402 ( .I1(n2948), .I2(n2147), .O(n2146) );
  AOI12X1 U1403 ( .B1(n2148), .B2(n2149), .A1(n2121), .O(n2147) );
  INVCKX1 U1404 ( .I(n2150), .O(n2121) );
  OAI112X1 U1405 ( .C1(n1954), .C2(n2151), .A1(n2152), .B1(n2153), .O(n2149)
         );
  XNR2X1 U1406 ( .I1(n2948), .I2(n1889), .O(n2151) );
  NR2X1 U1407 ( .I1(n2154), .I2(n2115), .O(g9124) );
  XNR2X1 U1408 ( .I1(n3156), .I2(n2155), .O(n2154) );
  OA13X1 U1409 ( .B1(n2156), .B2(n2157), .B3(n2158), .A1(n2159), .O(n2155) );
  NR2X1 U1410 ( .I1(n2160), .I2(n2115), .O(g9110) );
  XNR2X1 U1411 ( .I1(n3165), .I2(n2161), .O(n2160) );
  NR2X1 U1412 ( .I1(n2162), .I2(n2120), .O(n2161) );
  AOI112X1 U1413 ( .C1(n3156), .C2(n1889), .A1(n2119), .B1(n2156), .O(n2162)
         );
  NR2X1 U1414 ( .I1(n2163), .I2(n3156), .O(n2156) );
  OAI12X1 U1415 ( .B1(n2164), .B2(n2148), .A1(n2165), .O(g8973) );
  XNR2X1 U1416 ( .I1(n3170), .I2(n2166), .O(n2164) );
  AOI12X1 U1417 ( .B1(n2167), .B2(n1905), .A1(n2168), .O(n2166) );
  OAI12X1 U1418 ( .B1(n2169), .B2(n2170), .A1(n2171), .O(g8945) );
  XNR2X1 U1419 ( .I1(n3152), .I2(n2172), .O(n2169) );
  MUXB2X1 U1420 ( .EB(n2173), .A(n2174), .B(n3140), .S(n2175), .O(n2172) );
  ND2X1 U1421 ( .I1(n2176), .I2(n2177), .O(n2174) );
  OAI12X1 U1422 ( .B1(n2178), .B2(n2170), .A1(n2171), .O(g8944) );
  XNR2X1 U1423 ( .I1(n2885), .I2(n2179), .O(n2178) );
  MUXB2X1 U1424 ( .EB(n2173), .A(n2180), .B(n3157), .S(n2175), .O(n2179) );
  MXL2XLP U1425 ( .A(n2181), .B(n2182), .S(n2886), .OB(n2180) );
  OR2X1 U1426 ( .I1(n2183), .I2(n2184), .O(n2182) );
  ND2X1 U1427 ( .I1(n2185), .I2(n2186), .O(n2181) );
  OAI12X1 U1428 ( .B1(n2187), .B2(n2170), .A1(n2171), .O(g8943) );
  AOI23X1 U1429 ( .B1(n2188), .B2(n2189), .B3(n2190), .A1(n3119), .A2(n2191), 
        .O(n2187) );
  OR2B1XLP U1430 ( .I1(n2188), .B1(n2189), .O(n2191) );
  OAI12X1 U1431 ( .B1(n2192), .B2(n2193), .A1(n2194), .O(n2190) );
  MXL2XLP U1432 ( .A(n3164), .B(n2195), .S(n2196), .OB(n2194) );
  NR2X1 U1433 ( .I1(n3177), .I2(n2197), .O(n2195) );
  OAI112X1 U1434 ( .C1(n2197), .C2(n2193), .A1(n2198), .B1(n2199), .O(n2188)
         );
  AOI12X1 U1435 ( .B1(n2175), .B2(n1906), .A1(n1878), .O(n2199) );
  INVCKX1 U1436 ( .I(n2200), .O(n2193) );
  OAI12X1 U1437 ( .B1(n2201), .B2(n2170), .A1(n2171), .O(g8941) );
  XOR2X1 U1438 ( .I1(n2202), .I2(n2886), .O(n2201) );
  ND2X1 U1439 ( .I1(n2203), .I2(n2189), .O(n2202) );
  OAI222X1 U1440 ( .A1(n2183), .A2(n2204), .B1(n2205), .B2(n2206), .C1(n2196), 
        .C2(n1989), .O(n2203) );
  INVCKX1 U1441 ( .I(n2185), .O(n2205) );
  OAI12X1 U1442 ( .B1(n2207), .B2(n2170), .A1(n2171), .O(g8940) );
  XNR2X1 U1443 ( .I1(n3154), .I2(n2208), .O(n2207) );
  AOI12X1 U1444 ( .B1(n2209), .B2(n2210), .A1(n2173), .O(n2208) );
  ND2X1 U1445 ( .I1(n2895), .I2(n2175), .O(n2210) );
  MXL2XLP U1446 ( .A(n2211), .B(n2212), .S(n2887), .OB(n2209) );
  NR2X1 U1447 ( .I1(n1972), .I2(n2204), .O(n2212) );
  NR2X1 U1448 ( .I1(n3161), .I2(n2206), .O(n2211) );
  OAI12X1 U1449 ( .B1(n2213), .B2(n2170), .A1(n2171), .O(g8939) );
  XNR2X1 U1450 ( .I1(n2887), .I2(n2214), .O(n2213) );
  AOI12X1 U1451 ( .B1(n2215), .B2(n2216), .A1(n2173), .O(n2214) );
  ND2X1 U1452 ( .I1(n2896), .I2(n2175), .O(n2216) );
  MUX2X1 U1453 ( .A(n2206), .B(n2204), .S(n3161), .O(n2215) );
  OAI12X1 U1454 ( .B1(n2217), .B2(n2170), .A1(n2171), .O(g8938) );
  XNR2X1 U1455 ( .I1(n2218), .I2(n1972), .O(n2217) );
  ND2X1 U1456 ( .I1(n2189), .I2(n2219), .O(n2218) );
  OAI112X1 U1457 ( .C1(n2196), .C2(n1912), .A1(n2206), .B1(n2204), .O(n2219)
         );
  ND2X1 U1458 ( .I1(n2220), .I2(n2196), .O(n2204) );
  ND2X1 U1459 ( .I1(n2186), .I2(n2196), .O(n2206) );
  OAI12X1 U1460 ( .B1(n2221), .B2(n2170), .A1(n2171), .O(g8937) );
  XNR2X1 U1461 ( .I1(n3183), .I2(n2222), .O(n2221) );
  AOI112X1 U1462 ( .C1(n2200), .C2(n1878), .A1(n2223), .B1(n2224), .O(n2222)
         );
  MXL2XLP U1463 ( .A(n2897), .B(n2225), .S(n2196), .OB(n2224) );
  ND2X1 U1464 ( .I1(n2192), .I2(n3119), .O(n2225) );
  ND2X1 U1465 ( .I1(n2189), .I2(n2198), .O(n2223) );
  ND3X1 U1466 ( .I1(n2196), .I2(n1967), .I3(n2197), .O(n2198) );
  INVCKX1 U1467 ( .I(n2175), .O(n2196) );
  INVCKX1 U1468 ( .I(n2173), .O(n2189) );
  NR2X1 U1469 ( .I1(n1967), .I2(n2175), .O(n2200) );
  OAI12X1 U1470 ( .B1(n2226), .B2(n2148), .A1(n2165), .O(g8926) );
  XNR2X1 U1471 ( .I1(n3166), .I2(n2227), .O(n2226) );
  MUXB2X1 U1472 ( .EB(n2168), .A(n2228), .B(n3133), .S(n2167), .O(n2227) );
  ND2X1 U1473 ( .I1(n2229), .I2(n2230), .O(n2228) );
  OAI12X1 U1474 ( .B1(n2231), .B2(n2148), .A1(n2165), .O(g8923) );
  XNR2X1 U1475 ( .I1(n2888), .I2(n2232), .O(n2231) );
  MUXB2X1 U1476 ( .EB(n2168), .A(n2233), .B(n3174), .S(n2167), .O(n2232) );
  MXL2XLP U1477 ( .A(n2234), .B(n2235), .S(n1965), .OB(n2233) );
  ND3X1 U1478 ( .I1(n2236), .I2(n2237), .I3(n2889), .O(n2234) );
  OAI12X1 U1479 ( .B1(n2238), .B2(n2148), .A1(n2165), .O(g8922) );
  AOI23X1 U1480 ( .B1(n2239), .B2(n2240), .B3(n2241), .A1(n3168), .A2(n2242), 
        .O(n2238) );
  OR2B1XLP U1481 ( .I1(n2239), .B1(n2240), .O(n2242) );
  ND2X1 U1482 ( .I1(n3168), .I2(n2241), .O(n2239) );
  MUX2X1 U1483 ( .A(n2243), .B(n3181), .S(n2167), .O(n2241) );
  AO12X1 U1484 ( .B1(n2244), .B2(n3170), .A1(n2245), .O(n2243) );
  OAI12X1 U1485 ( .B1(n2246), .B2(n2170), .A1(n2171), .O(g8921) );
  OR4B2XLP U1486 ( .I1(n2247), .I2(n2138), .B1(n2170), .B2(n2248), .O(n2171)
         );
  NR2X1 U1487 ( .I1(n2139), .I2(n2249), .O(n2248) );
  NR2X1 U1488 ( .I1(n1890), .I2(n3189), .O(n2138) );
  INVCKX1 U1489 ( .I(n2133), .O(n2170) );
  NR2X1 U1490 ( .I1(n2247), .I2(n2126), .O(n2133) );
  AN2X1 U1491 ( .I1(n2250), .I2(n2251), .O(n2126) );
  MXL2XLP U1492 ( .A(n2177), .B(n2176), .S(n3152), .OB(n2250) );
  OR4B2XLP U1493 ( .I1(n2184), .I2(n2183), .B1(n2885), .B2(n2886), .O(n2176)
         );
  ND3X1 U1494 ( .I1(n3154), .I2(n3161), .I3(n2887), .O(n2183) );
  INVCKX1 U1495 ( .I(n2220), .O(n2184) );
  AN4B1XLP U1496 ( .I1(n3183), .I2(n2197), .I3(n3177), .B1(n1878), .O(n2220)
         );
  INVCKX1 U1497 ( .I(n2192), .O(n2197) );
  OR4B2XLP U1498 ( .I1(n2885), .I2(n2886), .B1(n2185), .B2(n2186), .O(n2177)
         );
  AN4B1XLP U1499 ( .I1(n1878), .I2(n1967), .I3(n2192), .B1(n3183), .O(n2186)
         );
  AOI12X1 U1500 ( .B1(n1961), .B2(n2135), .A1(n1890), .O(n2192) );
  NR3X1 U1501 ( .I1(n3154), .I2(n2887), .I3(n3161), .O(n2185) );
  XNR2X1 U1502 ( .I1(n3177), .I2(n2252), .O(n2246) );
  AOI12X1 U1503 ( .B1(n2175), .B2(n2003), .A1(n2173), .O(n2252) );
  NR2X1 U1504 ( .I1(n2251), .I2(n2175), .O(n2173) );
  ND2X1 U1505 ( .I1(n2253), .I2(n2144), .O(n2251) );
  ND2X1 U1506 ( .I1(n2249), .I2(n2124), .O(n2144) );
  NR3X1 U1507 ( .I1(n1871), .I2(n3147), .I3(n1962), .O(n2249) );
  OAI112X1 U1508 ( .C1(n3155), .C2(n3189), .A1(n2124), .B1(n3142), .O(n2253)
         );
  AOI12X1 U1509 ( .B1(n2254), .B2(n1953), .A1(n2127), .O(n2175) );
  OAI12X1 U1510 ( .B1(n2255), .B2(n2148), .A1(n2165), .O(g8920) );
  XOR2X1 U1511 ( .I1(n2256), .I2(n2889), .O(n2255) );
  OAI12X1 U1512 ( .B1(n2257), .B2(n2258), .A1(n2240), .O(n2256) );
  MXL2XLP U1513 ( .A(n2259), .B(n2260), .S(n1965), .OB(n2258) );
  ND2X1 U1514 ( .I1(n2261), .I2(n2262), .O(n2260) );
  ND2X1 U1515 ( .I1(n2263), .I2(n2236), .O(n2259) );
  NR2X1 U1516 ( .I1(n2264), .I2(n1882), .O(n2257) );
  OAI12X1 U1517 ( .B1(n2265), .B2(n2148), .A1(n2165), .O(g8889) );
  XNR2X1 U1518 ( .I1(n2891), .I2(n2266), .O(n2265) );
  NR2X1 U1519 ( .I1(n2267), .I2(n2168), .O(n2266) );
  AOI222X1 U1520 ( .A1(n2893), .A2(n2167), .B1(n2261), .B2(n2262), .C1(n2263), 
        .C2(n2236), .O(n2267) );
  INVCKX1 U1521 ( .I(n2268), .O(n2236) );
  OAI12X1 U1522 ( .B1(n2269), .B2(n2148), .A1(n2165), .O(g8887) );
  XOR2X1 U1523 ( .I1(n2270), .I2(n3122), .O(n2269) );
  OAI12X1 U1524 ( .B1(n2271), .B2(n2272), .A1(n2240), .O(n2270) );
  MXL2XLP U1525 ( .A(n2273), .B(n2274), .S(n2890), .OB(n2272) );
  ND2X1 U1526 ( .I1(n2263), .I2(n3158), .O(n2274) );
  OR2B1XLP U1527 ( .I1(n3158), .B1(n2261), .O(n2273) );
  NR2X1 U1528 ( .I1(n2264), .I2(n1916), .O(n2271) );
  OAI12X1 U1529 ( .B1(n2275), .B2(n2148), .A1(n2165), .O(g8885) );
  XNR2X1 U1530 ( .I1(n3158), .I2(n2276), .O(n2275) );
  AOI12X1 U1531 ( .B1(n2277), .B2(n2278), .A1(n2168), .O(n2276) );
  ND2X1 U1532 ( .I1(n2894), .I2(n2167), .O(n2278) );
  MXL2XLP U1533 ( .A(n2261), .B(n2263), .S(n2890), .OB(n2277) );
  OAI12X1 U1534 ( .B1(n2279), .B2(n2148), .A1(n2165), .O(g8883) );
  OR4B2XLP U1535 ( .I1(n2158), .I2(n2119), .B1(n2148), .B2(n2280), .O(n2165)
         );
  NR2X1 U1536 ( .I1(n2281), .I2(n2157), .O(n2280) );
  NR2X1 U1537 ( .I1(n1954), .I2(n2948), .O(n2158) );
  XNR2X1 U1538 ( .I1(n2890), .I2(n2282), .O(n2279) );
  NR2X1 U1539 ( .I1(n2283), .I2(n2168), .O(n2282) );
  INVCKX1 U1540 ( .I(n2240), .O(n2168) );
  ND2X1 U1541 ( .I1(n2284), .I2(n2264), .O(n2240) );
  AOI112X1 U1542 ( .C1(n3129), .C2(n2167), .A1(n2263), .B1(n2261), .O(n2283)
         );
  AN3B2X1 U1543 ( .I1(n2245), .B1(n2167), .B2(n3168), .O(n2261) );
  AN2X1 U1544 ( .I1(n2237), .I2(n2264), .O(n2263) );
  INVCKX1 U1545 ( .I(n2167), .O(n2264) );
  AOI12X1 U1546 ( .B1(n1968), .B2(n2285), .A1(n2118), .O(n2167) );
  OAI12X1 U1547 ( .B1(n2286), .B2(n1971), .A1(n2150), .O(g8820) );
  ND3X1 U1548 ( .I1(n2159), .I2(n1971), .I3(n2119), .O(n2150) );
  OA12X1 U1549 ( .B1(n2119), .B2(n2281), .A1(n2148), .O(n2286) );
  ND2X1 U1550 ( .I1(n2153), .I2(n2120), .O(n2148) );
  INVCKX1 U1551 ( .I(n2159), .O(n2120) );
  AN2B1XLP U1552 ( .I1(n2287), .B1(n2284), .O(n2159) );
  OAI12X1 U1553 ( .B1(n2119), .B2(n2288), .A1(n2289), .O(n2284) );
  OA12X1 U1554 ( .B1(n3156), .B2(n2948), .A1(n3132), .O(n2288) );
  MXL2XLP U1555 ( .A(n2230), .B(n2229), .S(n3166), .OB(n2287) );
  OR4B2XLP U1556 ( .I1(n1965), .I2(n2268), .B1(n2237), .B2(n2290), .O(n2229)
         );
  AN2X1 U1557 ( .I1(n2889), .I2(n2888), .O(n2290) );
  AN3X1 U1558 ( .I1(n3170), .I2(n2244), .I3(n3168), .O(n2237) );
  ND3X1 U1559 ( .I1(n3122), .I2(n3158), .I3(n2890), .O(n2268) );
  OR3X1 U1560 ( .I1(n2888), .I2(n2891), .I3(n2235), .O(n2230) );
  OR4B2XLP U1561 ( .I1(n3168), .I2(n2889), .B1(n2262), .B2(n2245), .O(n2235)
         );
  NR2X1 U1562 ( .I1(n2244), .I2(n3170), .O(n2245) );
  OAI12X1 U1563 ( .B1(n2948), .B2(n3165), .A1(n3156), .O(n2244) );
  NR3X1 U1564 ( .I1(n3122), .I2(n2890), .I3(n3158), .O(n2262) );
  NR3X1 U1565 ( .I1(n1889), .I2(n3149), .I3(n1963), .O(n2119) );
  MUX2X1 U1566 ( .A(n3011), .B(n2291), .S(n2292), .O(g8779) );
  MUX2X1 U1567 ( .A(n3051), .B(n2293), .S(n2292), .O(g8777) );
  MUX2X1 U1568 ( .A(n3053), .B(n2294), .S(n2292), .O(g8776) );
  NR2X1 U1569 ( .I1(n2295), .I2(n2296), .O(g8775) );
  XNR2X1 U1570 ( .I1(n2919), .I2(n2297), .O(n2296) );
  MUX2X1 U1571 ( .A(n3048), .B(n2297), .S(n2292), .O(g8774) );
  OAI12X1 U1572 ( .B1(g18), .B2(n2298), .A1(n2299), .O(n2297) );
  XOR2X1 U1573 ( .I1(n2300), .I2(n3184), .O(n2298) );
  ND2X1 U1574 ( .I1(n2301), .I2(n1891), .O(n2300) );
  MUX2X1 U1575 ( .A(n3013), .B(n2302), .S(n2292), .O(g8773) );
  NR2X1 U1576 ( .I1(n2295), .I2(n2303), .O(g8772) );
  XNR2X1 U1577 ( .I1(n2918), .I2(n2294), .O(n2303) );
  OAI12X1 U1578 ( .B1(g18), .B2(n2304), .A1(n2305), .O(n2294) );
  XNR2X1 U1579 ( .I1(n2306), .I2(n1908), .O(n2304) );
  ND2X1 U1580 ( .I1(n2301), .I2(n3141), .O(n2306) );
  AN2X1 U1581 ( .I1(n2307), .I2(n2953), .O(n2301) );
  MUX2X1 U1582 ( .A(n3015), .B(n2308), .S(n2292), .O(g8771) );
  MUX2X1 U1583 ( .A(n3017), .B(n2309), .S(n2292), .O(g8770) );
  NR2X1 U1584 ( .I1(n2295), .I2(n2310), .O(g8769) );
  XNR2X1 U1585 ( .I1(n2915), .I2(n2309), .O(n2310) );
  OAI12X1 U1586 ( .B1(g18), .B2(n2311), .A1(n2312), .O(n2309) );
  XNR2X1 U1587 ( .I1(n2313), .I2(n1982), .O(n2311) );
  ND2X1 U1588 ( .I1(n2314), .I2(n3141), .O(n2313) );
  NR2X1 U1589 ( .I1(n2295), .I2(n2315), .O(g8768) );
  XNR2X1 U1590 ( .I1(n2917), .I2(n2293), .O(n2315) );
  OAI12X1 U1591 ( .B1(g18), .B2(n2316), .A1(n2317), .O(n2293) );
  XNR2X1 U1592 ( .I1(n2957), .I2(n2318), .O(n2316) );
  NR2X1 U1593 ( .I1(n3126), .I2(n2319), .O(n2318) );
  NR2X1 U1594 ( .I1(n2295), .I2(n2320), .O(g8767) );
  XNR2X1 U1595 ( .I1(n2921), .I2(n2308), .O(n2320) );
  OAI12X1 U1596 ( .B1(g18), .B2(n2321), .A1(n2322), .O(n2308) );
  XNR2X1 U1597 ( .I1(n2959), .I2(n2323), .O(n2321) );
  NR2X1 U1598 ( .I1(n3141), .I2(n2324), .O(n2323) );
  NR2X1 U1599 ( .I1(n2295), .I2(n2325), .O(g8766) );
  XNR2X1 U1600 ( .I1(n2961), .I2(n2291), .O(n2325) );
  OAI12X1 U1601 ( .B1(g18), .B2(n2326), .A1(n2327), .O(n2291) );
  XNR2X1 U1602 ( .I1(n2958), .I2(n2328), .O(n2326) );
  AN2X1 U1603 ( .I1(n2329), .I2(n2952), .O(n2328) );
  NR2X1 U1604 ( .I1(n2295), .I2(n2330), .O(g8765) );
  XNR2X1 U1605 ( .I1(n2920), .I2(n2302), .O(n2330) );
  OAI12X1 U1606 ( .B1(g18), .B2(n2331), .A1(n2332), .O(n2302) );
  XNR2X1 U1607 ( .I1(n2960), .I2(n2333), .O(n2331) );
  NR2X1 U1608 ( .I1(n1891), .I2(n2324), .O(n2333) );
  ND3X1 U1609 ( .I1(n1893), .I2(n1964), .I3(n2953), .O(n2324) );
  OAI112X1 U1610 ( .C1(n2334), .C2(n1905), .A1(n2335), .B1(n2153), .O(g8649)
         );
  MXL2XLP U1611 ( .A(n2336), .B(n2337), .S(n2153), .OB(g8631) );
  AOI12X1 U1612 ( .B1(n2157), .B2(n1971), .A1(n2338), .O(n2337) );
  AOI13X1 U1613 ( .B1(n2339), .B2(n2340), .B3(g4892), .A1(n2892), .O(n2338) );
  OR4B2XLP U1614 ( .I1(n3136), .I2(n3156), .B1(n2163), .B2(n2285), .O(n2340)
         );
  XOR2X1 U1615 ( .I1(n2341), .I2(n2342), .O(n2339) );
  MXL2XLP U1616 ( .A(n2343), .B(n1889), .S(n3132), .OB(n2342) );
  ND2X1 U1617 ( .I1(n1963), .I2(n2163), .O(n2343) );
  ND2X1 U1618 ( .I1(n3127), .I2(g255), .O(n2341) );
  INVCKX1 U1619 ( .I(n2152), .O(n2157) );
  AOI112X1 U1620 ( .C1(n2344), .C2(n2345), .A1(n1674), .B1(n2346), .O(n2336)
         );
  OA22X1 U1621 ( .A1(n1614), .A2(n1738), .B1(n1672), .B2(n1676), .O(n2346) );
  OR2B1XLP U1622 ( .I1(n1707), .B1(g802), .O(n2345) );
  ND2X1 U1623 ( .I1(n2347), .I2(n2130), .O(g8559) );
  MXL2XLP U1624 ( .A(n3140), .B(n2898), .S(n2348), .OB(n2347) );
  NR2X1 U1625 ( .I1(n2115), .I2(n2349), .O(g8505) );
  XNR2X1 U1626 ( .I1(n3149), .I2(n2350), .O(n2349) );
  OAI12X1 U1627 ( .B1(n2118), .B2(n2285), .A1(n2335), .O(n2350) );
  ND2X1 U1628 ( .I1(n3133), .I2(n2334), .O(n2335) );
  ND3X1 U1629 ( .I1(n3165), .I2(n1968), .I3(n2351), .O(n2285) );
  OAI22X1 U1630 ( .A1(n2352), .A2(n1922), .B1(n2077), .B2(n2353), .O(g8435) );
  OAI22X1 U1631 ( .A1(n1882), .A2(n2352), .B1(n2353), .B2(n1922), .O(g8434) );
  OAI22X1 U1632 ( .A1(n2029), .A2(n2352), .B1(n1882), .B2(n2353), .O(g8433) );
  OAI22X1 U1633 ( .A1(n1916), .A2(n2352), .B1(n2029), .B2(n2353), .O(g8432) );
  OAI22X1 U1634 ( .A1(n2027), .A2(n2352), .B1(n1916), .B2(n2353), .O(g8431) );
  OAI22X1 U1635 ( .A1(n1927), .A2(n2352), .B1(n2027), .B2(n2353), .O(g8430) );
  OAI22X1 U1636 ( .A1(n2030), .A2(n2352), .B1(n1927), .B2(n2353), .O(g8429) );
  OAI22X1 U1637 ( .A1(n2352), .A2(n1905), .B1(n2030), .B2(n2353), .O(g8428) );
  ND2X1 U1638 ( .I1(n2153), .I2(n2352), .O(n2353) );
  INVCKX1 U1639 ( .I(n2334), .O(n2352) );
  NR3X1 U1640 ( .I1(n2118), .I2(n3136), .I3(n1968), .O(n2334) );
  NR2X1 U1641 ( .I1(n2115), .I2(n2354), .O(g8384) );
  XNR2X1 U1642 ( .I1(n1953), .I2(n2355), .O(n2354) );
  OA22X1 U1643 ( .A1(n2006), .A2(n2348), .B1(n2254), .B2(n2127), .O(n2355) );
  OAI22X1 U1644 ( .A1(n2348), .A2(n1923), .B1(n2006), .B2(n2356), .O(g8288) );
  OAI22X1 U1645 ( .A1(n1989), .A2(n2348), .B1(n2356), .B2(n1923), .O(g8287) );
  OAI22X1 U1646 ( .A1(n1928), .A2(n2348), .B1(n1989), .B2(n2356), .O(g8286) );
  OAI22X1 U1647 ( .A1(n2028), .A2(n2348), .B1(n1928), .B2(n2356), .O(g8285) );
  OAI22X1 U1648 ( .A1(n1912), .A2(n2348), .B1(n2028), .B2(n2356), .O(g8284) );
  OAI22X1 U1649 ( .A1(n2348), .A2(n2005), .B1(n1912), .B2(n2356), .O(g8283) );
  OAI22X1 U1650 ( .A1(n1906), .A2(n2348), .B1(n2356), .B2(n2005), .O(g8282) );
  OAI22X1 U1651 ( .A1(n2348), .A2(n2003), .B1(n1906), .B2(n2356), .O(g8281) );
  ND2X1 U1652 ( .I1(n2130), .I2(n2348), .O(n2356) );
  ND3X1 U1653 ( .I1(n2124), .I2(n1962), .I3(n3147), .O(n2348) );
  AN2B1XLP U1654 ( .I1(n3124), .B1(n2357), .O(g8260) );
  AN2B1XLP U1655 ( .I1(n3162), .B1(n2357), .O(g8254) );
  AN2B1XLP U1656 ( .I1(n3092), .B1(n2357), .O(g8250) );
  NR2X1 U1657 ( .I1(n2358), .I2(n2359), .O(g8245) );
  XOR2X1 U1658 ( .I1(n1674), .I2(n2360), .O(n2359) );
  NR2X1 U1659 ( .I1(n1614), .I2(n2361), .O(n2360) );
  NR2X1 U1660 ( .I1(n2362), .I2(n2363), .O(g8244) );
  XNR2X1 U1661 ( .I1(n1743), .I2(n2113), .O(n2363) );
  OR2B1XLP U1662 ( .I1(n1661), .B1(n2364), .O(n2113) );
  ND2X1 U1663 ( .I1(n2047), .I2(n2365), .O(g8349) );
  ND2X1 U1664 ( .I1(n2035), .I2(n2365), .O(g8340) );
  ND2X1 U1665 ( .I1(n2042), .I2(n2365), .O(g8335) );
  ND2X1 U1666 ( .I1(n2036), .I2(n2365), .O(g8331) );
  ND2X1 U1667 ( .I1(n2043), .I2(n2365), .O(g8328) );
  ND2X1 U1668 ( .I1(n2037), .I2(n2365), .O(g8323) );
  ND2X1 U1669 ( .I1(n2044), .I2(n2365), .O(g8318) );
  ND2X1 U1670 ( .I1(n2038), .I2(n2365), .O(g8316) );
  ND2X1 U1671 ( .I1(n2045), .I2(n2365), .O(g8313) );
  ND2X1 U1672 ( .I1(n2039), .I2(n2365), .O(g8347) );
  MXL2XLP U1673 ( .A(n2041), .B(n2366), .S(n2292), .OB(g8194) );
  XNR2X1 U1674 ( .I1(n2956), .I2(n2367), .O(n2366) );
  NR2X1 U1675 ( .I1(n2319), .I2(n1893), .O(n2367) );
  ND3X1 U1676 ( .I1(n1891), .I2(n1966), .I3(n2952), .O(n2319) );
  MXL2XLP U1677 ( .A(n2021), .B(n2368), .S(n2292), .OB(g8193) );
  XNR2X1 U1678 ( .I1(n2369), .I2(n1913), .O(n2368) );
  ND2X1 U1679 ( .I1(n2314), .I2(n1891), .O(n2369) );
  AN2X1 U1680 ( .I1(n2307), .I2(n1966), .O(n2314) );
  NR2X1 U1681 ( .I1(n1893), .I2(n2952), .O(n2307) );
  ND2X1 U1682 ( .I1(n2046), .I2(n2365), .O(g8352) );
  INVCKX1 U1683 ( .I(g82), .O(n2365) );
  NR2X1 U1684 ( .I1(n2370), .I2(g1713), .O(g8173) );
  XNR2X1 U1685 ( .I1(n2997), .I2(n2371), .O(n2370) );
  AN2B1XLP U1686 ( .I1(n2995), .B1(n2372), .O(n2371) );
  NR2X1 U1687 ( .I1(n1979), .I2(n2357), .O(g8147) );
  OAI13X1 U1688 ( .B1(g114), .B2(g881), .B3(n2102), .A1(g109), .O(n2357) );
  INVCKX1 U1689 ( .I(n2373), .O(n2102) );
  NR2X1 U1690 ( .I1(n2295), .I2(n2374), .O(g8060) );
  XNR2X1 U1691 ( .I1(n2904), .I2(g6002), .O(n2374) );
  NR2X1 U1692 ( .I1(n2375), .I2(n2295), .O(g8059) );
  XNR2X1 U1693 ( .I1(g6042), .I2(n2907), .O(n2375) );
  NR2X1 U1694 ( .I1(n2295), .I2(n2376), .O(g8055) );
  XNR2X1 U1695 ( .I1(n2914), .I2(n2377), .O(n2376) );
  NR2X1 U1696 ( .I1(n2295), .I2(n2378), .O(g8054) );
  XNR2X1 U1697 ( .I1(n2902), .I2(g6015), .O(n2378) );
  NR2X1 U1698 ( .I1(n2379), .I2(n2295), .O(g8053) );
  XNR2X1 U1699 ( .I1(g6045), .I2(n2905), .O(n2379) );
  NR2X1 U1700 ( .I1(n2295), .I2(n2380), .O(g8052) );
  XNR2X1 U1701 ( .I1(n1910), .I2(n2381), .O(n2380) );
  NR2X1 U1702 ( .I1(n2295), .I2(n2382), .O(g8051) );
  XNR2X1 U1703 ( .I1(n1985), .I2(n2383), .O(n2382) );
  NR2X1 U1704 ( .I1(n2295), .I2(n2384), .O(g8050) );
  XNR2X1 U1705 ( .I1(n2901), .I2(g6026), .O(n2384) );
  NR2X1 U1706 ( .I1(n2385), .I2(n2295), .O(g8049) );
  XNR2X1 U1707 ( .I1(g6049), .I2(n2903), .O(n2385) );
  NR2X1 U1708 ( .I1(n2295), .I2(n2386), .O(g8048) );
  XNR2X1 U1709 ( .I1(n2924), .I2(g5996), .O(n2386) );
  NR2X1 U1710 ( .I1(n2295), .I2(n2387), .O(g8047) );
  XNR2X1 U1711 ( .I1(n2909), .I2(g6035), .O(n2387) );
  NR2X1 U1712 ( .I1(n2295), .I2(n2388), .O(g8046) );
  XOR2X1 U1713 ( .I1(n2912), .I2(n2389), .O(n2388) );
  NR2X1 U1714 ( .I1(n2295), .I2(n2390), .O(g8045) );
  XNR2X1 U1715 ( .I1(n1986), .I2(n2391), .O(n2390) );
  NR2X1 U1716 ( .I1(n2295), .I2(n2392), .O(g8044) );
  XNR2X1 U1717 ( .I1(n2908), .I2(g6038), .O(n2392) );
  NR2X1 U1718 ( .I1(n2295), .I2(n2393), .O(g8043) );
  XOR2X1 U1719 ( .I1(n2911), .I2(n2394), .O(n2393) );
  NR2X1 U1720 ( .I1(n2295), .I2(n2395), .O(g8042) );
  XNR2X1 U1721 ( .I1(n2913), .I2(n2396), .O(n2395) );
  NR2X1 U1722 ( .I1(n2295), .I2(n2397), .O(g8041) );
  XNR2X1 U1723 ( .I1(n2941), .I2(n2398), .O(n2397) );
  NR2X1 U1724 ( .I1(n2295), .I2(n2399), .O(g8040) );
  XOR2X1 U1725 ( .I1(n2916), .I2(n2400), .O(n2399) );
  NR2X1 U1726 ( .I1(n2295), .I2(n2401), .O(g8039) );
  XNR2X1 U1727 ( .I1(n1909), .I2(n2402), .O(n2401) );
  NR2X1 U1728 ( .I1(n2358), .I2(n2403), .O(g8024) );
  XNR2X1 U1729 ( .I1(n1614), .I2(n2361), .O(n2403) );
  OR2B1XLP U1730 ( .I1(n1738), .B1(n2404), .O(n2361) );
  NR2X1 U1731 ( .I1(n2362), .I2(n2405), .O(g8019) );
  XOR2X1 U1732 ( .I1(n1661), .I2(n2364), .O(n2405) );
  NR2X1 U1733 ( .I1(n2406), .I2(n1688), .O(n2364) );
  NR2X1 U1734 ( .I1(n2407), .I2(g1713), .O(g7930) );
  XOR2X1 U1735 ( .I1(n2372), .I2(n2995), .O(n2407) );
  ND2X1 U1736 ( .I1(n3186), .I2(n2408), .O(n2372) );
  NR2X1 U1737 ( .I1(n2295), .I2(n2409), .O(g7843) );
  XNR2X1 U1738 ( .I1(n2906), .I2(g6000), .O(n2409) );
  NR2X1 U1739 ( .I1(n2358), .I2(n2410), .O(g7709) );
  XOR2X1 U1740 ( .I1(n1738), .I2(n2404), .O(n2410) );
  NR2X1 U1741 ( .I1(n2411), .I2(n1676), .O(n2404) );
  NR2X1 U1742 ( .I1(n2362), .I2(n2412), .O(g7705) );
  XNR2X1 U1743 ( .I1(n1688), .I2(n2406), .O(n2412) );
  OR2B1XLP U1744 ( .I1(n1620), .B1(n2413), .O(n2406) );
  OAI12X1 U1745 ( .B1(n2414), .B2(n2001), .A1(n2415), .O(g7660) );
  MUXB2X1 U1746 ( .EB(n2951), .A(n2416), .B(n2417), .S(n2978), .O(g7632) );
  OAI12X1 U1747 ( .B1(n2295), .B2(n2418), .A1(n2419), .O(n2417) );
  NR2X1 U1748 ( .I1(n2295), .I2(n2420), .O(n2416) );
  ND2X1 U1749 ( .I1(n2421), .I2(n2153), .O(g7626) );
  MXL2XLP U1750 ( .A(n2422), .B(n2118), .S(n3132), .OB(n2421) );
  AOI13X1 U1751 ( .B1(n2152), .B2(n1954), .B3(n2163), .A1(n2118), .O(n2422) );
  ND2X1 U1752 ( .I1(n2948), .I2(n3165), .O(n2163) );
  ND3X1 U1753 ( .I1(n1889), .I2(n1954), .I3(n2948), .O(n2152) );
  NR2X1 U1754 ( .I1(n2423), .I2(n2424), .O(g7590) );
  AOI13X1 U1755 ( .B1(n2975), .B2(n2976), .B3(n2425), .A1(n2977), .O(n2423) );
  NR2X1 U1756 ( .I1(n2426), .I2(n2424), .O(g7586) );
  XNR2X1 U1757 ( .I1(n2976), .I2(n2427), .O(n2426) );
  NR2X1 U1758 ( .I1(n1994), .I2(n2428), .O(n2427) );
  NR2X1 U1759 ( .I1(n2429), .I2(n2424), .O(g7581) );
  OR2B1XLP U1760 ( .I1(n2951), .B1(g109), .O(n2424) );
  XNR2X1 U1761 ( .I1(n2975), .I2(n2425), .O(n2429) );
  INVCKX1 U1762 ( .I(n2428), .O(n2425) );
  ND3X1 U1763 ( .I1(n2978), .I2(n2418), .I3(n2430), .O(n2428) );
  INVCKX1 U1764 ( .I(n2431), .O(n2418) );
  NR2X1 U1765 ( .I1(n2432), .I2(g1713), .O(g7541) );
  XNR2X1 U1766 ( .I1(n3186), .I2(n2408), .O(n2432) );
  NR2X1 U1767 ( .I1(n2433), .I2(n2434), .O(n2408) );
  INVCKX1 U1768 ( .I(n2435), .O(n2434) );
  ND2X1 U1769 ( .I1(n2436), .I2(n2415), .O(g7441) );
  XNR2X1 U1770 ( .I1(n2900), .I2(n3143), .O(n2436) );
  OAI22X1 U1771 ( .A1(n1879), .A2(n2420), .B1(n1978), .B2(n2419), .O(g7303) );
  OAI22X1 U1772 ( .A1(n1903), .A2(n2420), .B1(n1879), .B2(n2419), .O(g7302) );
  OAI22X1 U1773 ( .A1(n1980), .A2(n2420), .B1(n1903), .B2(n2419), .O(g7301) );
  OAI22X1 U1774 ( .A1(n1869), .A2(n2420), .B1(n1980), .B2(n2419), .O(g7300) );
  OAI22X1 U1775 ( .A1(n1977), .A2(n2420), .B1(n1869), .B2(n2419), .O(g7299) );
  OAI22X1 U1776 ( .A1(n1877), .A2(n2420), .B1(n1977), .B2(n2419), .O(g7298) );
  OAI22X1 U1777 ( .A1(n1998), .A2(n2420), .B1(n1877), .B2(n2419), .O(g7297) );
  OAI22X1 U1778 ( .A1(n1896), .A2(n2420), .B1(n1998), .B2(n2419), .O(g7296) );
  OAI22X1 U1779 ( .A1(n1900), .A2(n2420), .B1(n2093), .B2(n2419), .O(g7295) );
  OAI22X1 U1780 ( .A1(n2420), .A2(n1988), .B1(n1900), .B2(n2419), .O(g7294) );
  OAI22X1 U1781 ( .A1(n2420), .A2(n1921), .B1(n2419), .B2(n1988), .O(g7293) );
  OAI22X1 U1782 ( .A1(n2420), .A2(n2007), .B1(n2419), .B2(n1921), .O(g7292) );
  OAI22X1 U1783 ( .A1(n2420), .A2(n1914), .B1(n2419), .B2(n2007), .O(g7291) );
  OAI22X1 U1784 ( .A1(n1978), .A2(n2420), .B1(n2419), .B2(n1914), .O(g7290) );
  MXL2XLP U1785 ( .A(n2063), .B(n1936), .S(n2292), .OB(g7257) );
  MUX2X1 U1786 ( .A(n3001), .B(n2938), .S(n2292), .O(g7244) );
  ND2X1 U1787 ( .I1(n2035), .I2(n2437), .O(g7219) );
  ND2X1 U1788 ( .I1(n2036), .I2(n2437), .O(g7204) );
  NR2X1 U1789 ( .I1(n2358), .I2(n2438), .O(g7202) );
  XNR2X1 U1790 ( .I1(n1676), .I2(n2411), .O(n2438) );
  OR2B1XLP U1791 ( .I1(n1672), .B1(n2439), .O(n2411) );
  NR2X1 U1792 ( .I1(n2362), .I2(n2440), .O(g7191) );
  XOR2X1 U1793 ( .I1(n1620), .I2(n2413), .O(n2440) );
  NR2X1 U1794 ( .I1(n2441), .I2(n1719), .O(n2413) );
  ND2X1 U1795 ( .I1(n2037), .I2(n2437), .O(g7189) );
  ND2X1 U1796 ( .I1(n2038), .I2(n2437), .O(g7183) );
  ND2X1 U1797 ( .I1(n2039), .I2(n2437), .O(g7143) );
  NR2X1 U1798 ( .I1(n2442), .I2(n2443), .O(g7137) );
  AOI12X1 U1799 ( .B1(n2899), .B2(n2444), .A1(n2414), .O(n2442) );
  AOI12X1 U1800 ( .B1(n2444), .B2(n2445), .A1(n2443), .O(g7134) );
  INVCKX1 U1801 ( .I(n2415), .O(n2443) );
  NR2X1 U1802 ( .I1(n2289), .I2(n2281), .O(n2415) );
  INVCKX1 U1803 ( .I(n2153), .O(n2281) );
  INVCKX1 U1804 ( .I(n2118), .O(n2289) );
  ND2X1 U1805 ( .I1(n2414), .I2(n2001), .O(n2118) );
  NR2X1 U1806 ( .I1(n2444), .I2(n2899), .O(n2414) );
  OAI12X1 U1807 ( .B1(n2900), .B2(n2004), .A1(n3130), .O(n2445) );
  OR3X1 U1808 ( .I1(n3130), .I2(n2900), .I3(n2004), .O(n2444) );
  ND2X1 U1809 ( .I1(n2446), .I2(n1823), .O(g7133) );
  XNR2X1 U1810 ( .I1(n2447), .I2(n2993), .O(n2446) );
  OAI23X1 U1811 ( .B1(n2448), .B2(n2449), .B3(n2450), .A1(n2295), .A2(n2100), 
        .O(g7032) );
  OR4B2XLP U1812 ( .I1(n2908), .I2(n2909), .B1(n1883), .B2(n1981), .O(n2450)
         );
  OR4B2XLP U1813 ( .I1(n2904), .I2(n2907), .B1(n1934), .B2(n2008), .O(n2449)
         );
  OR4B2XLP U1814 ( .I1(n2451), .I2(n2073), .B1(g6786), .B2(n2452), .O(n2448)
         );
  AN4B1XLP U1815 ( .I1(n2903), .I2(n2901), .I3(n1911), .B1(n2009), .O(n2452)
         );
  NR2X1 U1816 ( .I1(n2453), .I2(g1713), .O(g6983) );
  XNR2X1 U1817 ( .I1(n2996), .I2(n2454), .O(n2453) );
  NR2X1 U1818 ( .I1(n1874), .I2(n2433), .O(n2454) );
  MUX2X1 U1819 ( .A(n2901), .B(n3109), .S(n2455), .O(g6934) );
  MUX2X1 U1820 ( .A(n3006), .B(n2929), .S(n2292), .O(g6930) );
  MUX2X1 U1821 ( .A(n2925), .B(n3071), .S(n2455), .O(g6929) );
  MXL2XLP U1822 ( .A(n2009), .B(n1933), .S(n2455), .OB(g6928) );
  MUX2X1 U1823 ( .A(n3005), .B(n2930), .S(n2292), .O(g6924) );
  MUX2X1 U1824 ( .A(n2903), .B(n3073), .S(n2455), .O(g6923) );
  MUX2X1 U1825 ( .A(n2904), .B(n3070), .S(n2455), .O(g6922) );
  MUX2X1 U1826 ( .A(n3008), .B(n2931), .S(n2292), .O(g6918) );
  MXL2XLP U1827 ( .A(n1934), .B(n2058), .S(n2455), .OB(g6916) );
  MXL2XLP U1828 ( .A(n2008), .B(n1945), .S(n2455), .OB(g6915) );
  MUX2X1 U1829 ( .A(n3007), .B(n2932), .S(n2292), .O(g6912) );
  MUX2X1 U1830 ( .A(n2907), .B(n3087), .S(n2455), .O(g6911) );
  MXL2XLP U1831 ( .A(n1883), .B(n1931), .S(n2455), .OB(g6910) );
  OAI12X1 U1832 ( .B1(n2456), .B2(n2002), .A1(n2457), .O(g6909) );
  MUX2X1 U1833 ( .A(n3004), .B(n2933), .S(n2292), .O(g6908) );
  MUX2X1 U1834 ( .A(n2908), .B(n3096), .S(n2455), .O(g6907) );
  MXL2XLP U1835 ( .A(n1981), .B(n1932), .S(n2455), .OB(g6906) );
  MUX2X1 U1836 ( .A(n3009), .B(n2934), .S(n2292), .O(g6902) );
  MUX2X1 U1837 ( .A(n2909), .B(n3100), .S(n2455), .O(g6901) );
  MUX2X1 U1838 ( .A(n2910), .B(n3097), .S(n2455), .O(g6900) );
  MUX2X1 U1839 ( .A(n3010), .B(n2935), .S(n2292), .O(g6898) );
  MUX2X1 U1840 ( .A(n2923), .B(n3099), .S(n2455), .O(g6897) );
  ND2X1 U1841 ( .I1(n2458), .I2(n1997), .O(n2451) );
  MUX2X1 U1842 ( .A(n3003), .B(n2936), .S(n2292), .O(g6895) );
  MUX2X1 U1843 ( .A(n3002), .B(n2937), .S(n2292), .O(g6894) );
  NR2X1 U1844 ( .I1(n2295), .I2(n2067), .O(g6841) );
  NR2X1 U1845 ( .I1(n2295), .I2(n1907), .O(g6840) );
  AN2X1 U1846 ( .I1(n2945), .I2(g109), .O(g6839) );
  NR2X1 U1847 ( .I1(n2295), .I2(n1880), .O(g6838) );
  NR2X1 U1848 ( .I1(n2295), .I2(n1888), .O(g6834) );
  AN2X1 U1849 ( .I1(n3019), .I2(g109), .O(g6833) );
  NR2X1 U1850 ( .I1(n2295), .I2(n2074), .O(g6832) );
  NR2X1 U1851 ( .I1(n2295), .I2(n2061), .O(g6831) );
  AN2X1 U1852 ( .I1(n2944), .I2(g109), .O(g6830) );
  NR2X1 U1853 ( .I1(n2295), .I2(n2078), .O(g6829) );
  AN2X1 U1854 ( .I1(n2943), .I2(g109), .O(g6828) );
  NR2X1 U1855 ( .I1(n2295), .I2(n2070), .O(g6827) );
  NR2X1 U1856 ( .I1(n2295), .I2(n1943), .O(g6826) );
  NR2X1 U1857 ( .I1(n2295), .I2(n1944), .O(g6824) );
  NR2X1 U1858 ( .I1(n2295), .I2(n1951), .O(g6823) );
  AN2X1 U1859 ( .I1(n3049), .I2(g109), .O(g6822) );
  AN2X1 U1860 ( .I1(n3054), .I2(g109), .O(g6821) );
  NR2X1 U1861 ( .I1(n2295), .I2(n2064), .O(g6820) );
  AN2X1 U1862 ( .I1(n3052), .I2(g109), .O(g6819) );
  NR2X1 U1863 ( .I1(n2459), .I2(n2460), .O(g6795) );
  AOI12X1 U1864 ( .B1(n2992), .B2(n2461), .A1(n2456), .O(n2459) );
  AN2B1XLP U1865 ( .I1(n2910), .B1(n2295), .O(g6786) );
  NR2X1 U1866 ( .I1(n2295), .I2(n1981), .O(g6759) );
  NR2X1 U1867 ( .I1(n2295), .I2(n1911), .O(g6757) );
  ND2X1 U1868 ( .I1(n2462), .I2(n1970), .O(g6755) );
  AOI112X1 U1869 ( .C1(n1584), .C2(n2031), .A1(n2295), .B1(n3179), .O(g6747)
         );
  NR2X1 U1870 ( .I1(n2358), .I2(n2463), .O(g6733) );
  XOR2X1 U1871 ( .I1(n1672), .I2(n2439), .O(n2463) );
  NR2X1 U1872 ( .I1(n2464), .I2(n1707), .O(n2439) );
  NR2X1 U1873 ( .I1(n2362), .I2(n2465), .O(g6728) );
  XNR2X1 U1874 ( .I1(n1719), .I2(n2441), .O(n2465) );
  OR3B1XLP U1875 ( .I1(n1724), .I2(n1731), .B1(n2466), .O(n2441) );
  OAI23X1 U1876 ( .B1(n2467), .B2(n2468), .B3(n2469), .A1(n2295), .A2(n2099), 
        .O(g6679) );
  OR4B2XLP U1877 ( .I1(n1885), .I2(n2034), .B1(n2918), .B2(n2915), .O(n2469)
         );
  OR4B2XLP U1878 ( .I1(n2921), .I2(n2964), .B1(n1919), .B2(n2032), .O(n2468)
         );
  OR4B2XLP U1879 ( .I1(n1917), .I2(n2065), .B1(n2962), .B2(n2470), .O(n2467)
         );
  AN4B1XLP U1880 ( .I1(n2920), .I2(n2961), .I3(g6234), .B1(n2471), .O(n2470)
         );
  OR2X1 U1881 ( .I1(g4117), .I2(n3143), .O(g6672) );
  OAI23X1 U1882 ( .B1(n2472), .B2(n2473), .B3(n2474), .A1(n2295), .A2(n2101), 
        .O(g6656) );
  OR4B2XLP U1883 ( .I1(n2939), .I2(n1986), .B1(n2911), .B2(n2914), .O(n2474)
         );
  OR4B2XLP U1884 ( .I1(n2912), .I2(n2913), .B1(n1985), .B2(n1910), .O(n2473)
         );
  OR4B2XLP U1885 ( .I1(n2475), .I2(n1987), .B1(n3145), .B2(g6215), .O(n2472)
         );
  OR4B2XLP U1886 ( .I1(n1909), .I2(n2471), .B1(n2941), .B2(n2916), .O(n2475)
         );
  NR2X1 U1887 ( .I1(n2476), .I2(n2042), .O(g6653) );
  NR2X1 U1888 ( .I1(n2476), .I2(n2043), .O(g6638) );
  NR2X1 U1889 ( .I1(n2476), .I2(n2044), .O(g6627) );
  NR2X1 U1890 ( .I1(n2476), .I2(n2045), .O(g6621) );
  MUX2X1 U1891 ( .A(n2911), .B(n3112), .S(n2479), .O(g6551) );
  MUX2X1 U1892 ( .A(n2940), .B(n3065), .S(n2479), .O(g6546) );
  MUX2X1 U1893 ( .A(n2912), .B(n3115), .S(n2479), .O(g6545) );
  MUX2X1 U1894 ( .A(n2913), .B(n3074), .S(n2479), .O(g6542) );
  MXL2XLP U1895 ( .A(n1910), .B(n2056), .S(n2479), .OB(g6541) );
  MXL2XLP U1896 ( .A(n1986), .B(n1886), .S(n2479), .OB(g6538) );
  MUX2X1 U1897 ( .A(n2914), .B(n3072), .S(n2479), .O(g6537) );
  MXL2XLP U1898 ( .A(n1985), .B(n1887), .S(n2479), .OB(g6534) );
  MUX2X1 U1899 ( .A(n2941), .B(n3079), .S(n2479), .O(g6533) );
  NR2X1 U1900 ( .I1(n2476), .I2(n2046), .O(g6531) );
  MXL2XLP U1901 ( .A(n1909), .B(n2059), .S(n2479), .OB(g6529) );
  MUX2X1 U1902 ( .A(n2939), .B(n3085), .S(n2479), .O(g6528) );
  NR2X1 U1903 ( .I1(n2476), .I2(n2047), .O(g6526) );
  INVCKX1 U1904 ( .I(n2437), .O(n2476) );
  NR2X1 U1905 ( .I1(n2477), .I2(g1713), .O(g6525) );
  XNR2X1 U1906 ( .I1(n2433), .I2(n1874), .O(n2477) );
  ND2X1 U1907 ( .I1(n3160), .I2(n2478), .O(n2433) );
  MUX2X1 U1908 ( .A(n2915), .B(n3111), .S(n2479), .O(g6524) );
  MUX2X1 U1909 ( .A(n2916), .B(n3102), .S(n2479), .O(g6523) );
  MUX2X1 U1910 ( .A(n2928), .B(n3182), .S(n2479), .O(g6522) );
  NR2X1 U1911 ( .I1(n2480), .I2(g1713), .O(g6516) );
  XNR2X1 U1912 ( .I1(n3160), .I2(n2478), .O(n2480) );
  NR2X1 U1913 ( .I1(n1956), .I2(n2481), .O(n2478) );
  MUX2X1 U1914 ( .A(n2961), .B(n3067), .S(n2479), .O(g6515) );
  MUX2X1 U1915 ( .A(n2927), .B(n3114), .S(n2479), .O(g6514) );
  MUX2X1 U1916 ( .A(n3145), .B(n3098), .S(n2479), .O(g6513) );
  NR2X1 U1917 ( .I1(n2482), .I2(g1713), .O(g6508) );
  XNR2X1 U1918 ( .I1(n2481), .I2(n1956), .O(n2482) );
  ND2X1 U1919 ( .I1(n3151), .I2(n2483), .O(n2481) );
  MXL2XLP U1920 ( .A(n2034), .B(n1930), .S(n2479), .OB(g6507) );
  MXL2XLP U1921 ( .A(n2010), .B(n1929), .S(n2479), .OB(g6506) );
  NR2X1 U1922 ( .I1(n2484), .I2(g1713), .O(g6502) );
  XNR2X1 U1923 ( .I1(n3151), .I2(n2483), .O(n2484) );
  NR2X1 U1924 ( .I1(n1901), .I2(n2485), .O(n2483) );
  MUX2X1 U1925 ( .A(n2918), .B(n3078), .S(n2479), .O(g6501) );
  MXL2XLP U1926 ( .A(n1919), .B(n2057), .S(n2479), .OB(g6500) );
  MXL2XLP U1927 ( .A(n1885), .B(n1946), .S(n2479), .OB(g6481) );
  MUX2X1 U1928 ( .A(n2962), .B(n3080), .S(n2479), .O(g6480) );
  MUX2X1 U1929 ( .A(n2920), .B(n3089), .S(n2479), .O(g6479) );
  MUX2X1 U1930 ( .A(n2963), .B(n3086), .S(n2479), .O(g6478) );
  NR2X1 U1931 ( .I1(n2486), .I2(n2460), .O(g6471) );
  INVCKX1 U1932 ( .I(n2457), .O(n2460) );
  AOI12X1 U1933 ( .B1(n3137), .B2(n1970), .A1(n2487), .O(n2486) );
  MUX2X1 U1934 ( .A(n2921), .B(n3104), .S(n2479), .O(g6470) );
  MUX2X1 U1935 ( .A(n2926), .B(n3095), .S(n2479), .O(g6469) );
  MUX2X1 U1936 ( .A(n2964), .B(n3101), .S(n2479), .O(g6468) );
  AN2X1 U1937 ( .I1(n2471), .I2(g109), .O(n2479) );
  ND2X1 U1938 ( .I1(n2458), .I2(n1996), .O(n2471) );
  NR2X1 U1939 ( .I1(n2488), .I2(n2295), .O(g6439) );
  XOR4XLP U1940 ( .I1(n1883), .I2(n1911), .I3(n2073), .I4(n2922), .O(n2488) );
  NR2X1 U1941 ( .I1(n2295), .I2(n2025), .O(g6334) );
  NR2X1 U1942 ( .I1(n2295), .I2(n1984), .O(g6333) );
  AN2X1 U1943 ( .I1(n2946), .I2(g109), .O(g6332) );
  NR2X1 U1944 ( .I1(n2295), .I2(n1919), .O(g6244) );
  ND2X1 U1945 ( .I1(n2489), .I2(n2490), .O(g6243) );
  XNR2X1 U1946 ( .I1(n1812), .I2(n1651), .O(n2489) );
  NR2X1 U1947 ( .I1(n2010), .I2(n2295), .O(g6234) );
  NR2X1 U1948 ( .I1(n2295), .I2(n2065), .O(g6224) );
  NR2X1 U1949 ( .I1(n2295), .I2(n2032), .O(g6216) );
  AN2B1XLP U1950 ( .I1(n2928), .B1(n2295), .O(g6215) );
  NR2X1 U1951 ( .I1(n2295), .I2(n1917), .O(g6205) );
  AN2X1 U1952 ( .I1(n2939), .I2(g109), .O(g6198) );
  AN2X1 U1953 ( .I1(n2962), .I2(g109), .O(g6193) );
  NR2X1 U1954 ( .I1(n2295), .I2(n1987), .O(g6180) );
  NR2X1 U1955 ( .I1(n2491), .I2(n2031), .O(g6179) );
  INVCKX1 U1956 ( .I(n2491), .O(g6163) );
  ND3X1 U1957 ( .I1(n2492), .I2(n2025), .I3(g6331), .O(n2491) );
  NR2X1 U1958 ( .I1(n1999), .I2(n2295), .O(g6331) );
  MXL2XLP U1959 ( .A(n2493), .B(n2494), .S(n1870), .OB(g6155) );
  ND2X1 U1960 ( .I1(n2949), .I2(g1700), .O(n2494) );
  INVCKX1 U1961 ( .I(g4076), .O(n2493) );
  MXL2XLP U1962 ( .A(n2495), .B(n2496), .S(n1707), .OB(g6126) );
  ND3X1 U1963 ( .I1(g798), .I2(g802), .I3(n2103), .O(n2496) );
  ND2X1 U1964 ( .I1(n2490), .I2(n2464), .O(n2495) );
  OR2X1 U1965 ( .I1(n2344), .I2(n1727), .O(n2464) );
  MXL2XLP U1966 ( .A(n2497), .B(n2498), .S(n1731), .OB(g6123) );
  OR3B2X1 U1967 ( .I1(n1724), .B1(n2466), .B2(n2499), .O(n2498) );
  AOI12X1 U1968 ( .B1(n1724), .B2(n2499), .A1(n2500), .O(n2497) );
  MUX2X1 U1969 ( .A(n2965), .B(n2929), .S(n2501), .O(g6099) );
  MUX2X1 U1970 ( .A(n2966), .B(n2930), .S(n2501), .O(g6096) );
  MUX2X1 U1971 ( .A(n2967), .B(n2931), .S(n2501), .O(g6093) );
  MUX2X1 U1972 ( .A(n2968), .B(n2932), .S(n2501), .O(g6088) );
  MUX2X1 U1973 ( .A(n2969), .B(n2933), .S(n2501), .O(g6080) );
  MUX2X1 U1974 ( .A(n2970), .B(n2934), .S(n2501), .O(g6071) );
  MUX2X1 U1975 ( .A(n2971), .B(n2935), .S(n2501), .O(g6068) );
  MUX2X1 U1976 ( .A(n2972), .B(n2936), .S(n2501), .O(g6059) );
  MUX2X1 U1977 ( .A(n2950), .B(n2937), .S(n2501), .O(g6054) );
  MXL2XLP U1978 ( .A(n2053), .B(n1880), .S(g18), .OB(g6049) );
  MXL2XLP U1979 ( .A(n2054), .B(n1907), .S(g18), .OB(g6045) );
  MUX2X1 U1980 ( .A(n3050), .B(n3052), .S(g18), .O(g6042) );
  OAI12X1 U1981 ( .B1(g18), .B2(n2024), .A1(n2327), .O(g6038) );
  OAI12X1 U1982 ( .B1(g18), .B2(n2016), .A1(n2317), .O(g6035) );
  OAI12X1 U1983 ( .B1(g18), .B2(n2017), .A1(n2305), .O(g6026) );
  OAI12X1 U1984 ( .B1(g18), .B2(n2018), .A1(n2299), .O(g6015) );
  OAI12X1 U1985 ( .B1(g18), .B2(n2019), .A1(n2332), .O(g6002) );
  OAI12X1 U1986 ( .B1(g18), .B2(n2020), .A1(n2322), .O(g6000) );
  OAI12X1 U1987 ( .B1(g18), .B2(n2022), .A1(n2312), .O(g5996) );
  OAI12X1 U1988 ( .B1(n2295), .B2(n1997), .A1(n2502), .O(g5918) );
  MXL2XLP U1989 ( .A(n2040), .B(n1936), .S(n2501), .OB(g5914) );
  MUX2X1 U1990 ( .A(n2973), .B(n2938), .S(n2501), .O(g5910) );
  NR2X1 U1991 ( .I1(n2503), .I2(n2295), .O(g5770) );
  XOR4XLP U1992 ( .I1(n2939), .I2(n1987), .I3(n3145), .I4(n2941), .O(n2503) );
  NR2X1 U1993 ( .I1(n2295), .I2(n2504), .O(g5755) );
  XOR4XLP U1994 ( .I1(n2942), .I2(n1984), .I3(n3171), .I4(n2505), .O(n2504) );
  AO12X1 U1995 ( .B1(n1999), .B2(n2492), .A1(n3131), .O(n2505) );
  AN4B2X1 U1996 ( .I1(n2506), .I2(n2507), .B1(n2508), .B2(n2509), .O(n2492) );
  OR4B2XLP U1997 ( .I1(n2945), .I2(n2946), .B1(n2510), .B2(n2067), .O(n2509)
         );
  NR2X1 U1998 ( .I1(n2943), .I2(n2944), .O(n2510) );
  OR4B2XLP U1999 ( .I1(n3054), .I2(n3052), .B1(n2061), .B2(n2511), .O(n2508)
         );
  NR2X1 U2000 ( .I1(n3019), .I2(n3049), .O(n2511) );
  AN4B2X1 U2001 ( .I1(n2074), .I2(n1951), .B1(n2942), .B2(n2512), .O(n2507) );
  ND3X1 U2002 ( .I1(n2064), .I2(n1944), .I3(n1888), .O(n2512) );
  AN4B2X1 U2003 ( .I1(n2070), .I2(n1943), .B1(n3018), .B2(n2513), .O(n2506) );
  ND3X1 U2004 ( .I1(n1880), .I2(n1984), .I3(n1907), .O(n2513) );
  AN4B1XLP U2005 ( .I1(n2994), .I2(n2514), .I3(n2435), .B1(n2515), .O(g5556)
         );
  ND3X1 U2006 ( .I1(n2993), .I2(n1992), .I3(n3151), .O(n2515) );
  AN4B2X1 U2007 ( .I1(n2949), .I2(n3153), .B1(n1993), .B2(n2516), .O(n2514) );
  ND2X1 U2008 ( .I1(n2995), .I2(n3186), .O(n2516) );
  MXL2XLP U2009 ( .A(n2517), .B(n2518), .S(g802), .OB(g5543) );
  ND2X1 U2010 ( .I1(n2490), .I2(n2344), .O(n2518) );
  OR2X1 U2011 ( .I1(n1812), .I2(n1651), .O(n2344) );
  INVCKX1 U2012 ( .I(n2358), .O(n2490) );
  ND2X1 U2013 ( .I1(n2103), .I2(g798), .O(n2517) );
  NR2X1 U2014 ( .I1(n2358), .I2(n1812), .O(n2103) );
  OR3B2X1 U2015 ( .I1(n1794), .B1(g745), .B2(g109), .O(n2358) );
  MXL2XLP U2016 ( .A(n2519), .B(n2520), .S(n1724), .OB(g5536) );
  ND2X1 U2017 ( .I1(n2499), .I2(n2466), .O(n2520) );
  INVCKX1 U2018 ( .I(n2500), .O(n2519) );
  NR2X1 U2019 ( .I1(n2362), .I2(n2466), .O(n2500) );
  NR2X1 U2020 ( .I1(n1742), .I2(n1836), .O(n2466) );
  MXL2XLP U2021 ( .A(n2521), .B(n2522), .S(n1742), .OB(g5529) );
  OR2X1 U2022 ( .I1(n1836), .I2(n2362), .O(n2522) );
  INVCKX1 U2023 ( .I(n2499), .O(n2362) );
  OAI12X1 U2024 ( .B1(n2295), .B2(n1996), .A1(n2502), .O(g5445) );
  OAI12B2X1 U2025 ( .B1(g109), .B2(n3084), .A1(n2502), .O(g5421) );
  ND2X1 U2026 ( .I1(n2458), .I2(g109), .O(n2502) );
  AN2X1 U2027 ( .I1(n3179), .I2(g18), .O(n2458) );
  MXL2XLP U2028 ( .A(n1958), .B(n1823), .S(n2292), .OB(g5404) );
  MXL2XLP U2029 ( .A(n1823), .B(n1426), .S(n2292), .OB(g5396) );
  INVCKX1 U2030 ( .I(n2523), .O(g5392) );
  NR2X1 U2031 ( .I1(n1891), .I2(n2524), .O(g5390) );
  NR2X1 U2032 ( .I1(g1696), .I2(g4089), .O(g6842) );
  AN2X1 U2033 ( .I1(n3159), .I2(n2485), .O(g5194) );
  NR2X1 U2034 ( .I1(n1964), .I2(n2524), .O(g5173) );
  NR2X1 U2035 ( .I1(n1966), .I2(n2524), .O(g5148) );
  NR2X1 U2036 ( .I1(n1893), .I2(n2524), .O(g5126) );
  ND2X1 U2037 ( .I1(g109), .I2(n1606), .O(n2524) );
  AOI12X1 U2038 ( .B1(n2501), .B2(n2485), .A1(g4089), .O(g5083) );
  INVCKX1 U2039 ( .I(n2521), .O(g4940) );
  ND2X1 U2040 ( .I1(n1836), .I2(n2499), .O(n2521) );
  NR2X1 U2041 ( .I1(n2295), .I2(n2947), .O(n2499) );
  NR2X1 U2042 ( .I1(g3524), .I2(n1576), .O(g4905) );
  NR2X1 U2043 ( .I1(g3524), .I2(n1405), .O(g4903) );
  NR2X1 U2044 ( .I1(g3524), .I2(n1549), .O(g4902) );
  NR2X1 U2045 ( .I1(g4117), .I2(n1525), .O(g4893) );
  AN2B1XLP U2046 ( .I1(g632), .B1(g4117), .O(g4892) );
  NR2X1 U2047 ( .I1(g4117), .I2(n1508), .O(g4891) );
  NR2X1 U2048 ( .I1(g4117), .I2(n1434), .O(g4890) );
  OR2X1 U2049 ( .I1(n2974), .I2(n2951), .O(g4556) );
  NR2X1 U2050 ( .I1(n2295), .I2(n2033), .O(g4506) );
  AN2B1XLP U2051 ( .I1(n3055), .B1(n2292), .O(g4500) );
  NR2X1 U2052 ( .I1(n2295), .I2(n1924), .O(g4498) );
  NR2X1 U2053 ( .I1(n2295), .I2(n2076), .O(g4490) );
  NR2X1 U2054 ( .I1(n2295), .I2(n1908), .O(g4484) );
  AN2B1XLP U2055 ( .I1(n3184), .B1(n2295), .O(g4480) );
  NR2X1 U2056 ( .I1(n2295), .I2(n1884), .O(g4477) );
  NR2X1 U2057 ( .I1(n2295), .I2(n2013), .O(g4473) );
  NR2X1 U2058 ( .I1(n2295), .I2(n1982), .O(g4471) );
  NR2X1 U2059 ( .I1(n2295), .I2(n1913), .O(g4465) );
  AN2X1 U2060 ( .I1(n3169), .I2(g109), .O(g4342) );
  AN2X1 U2061 ( .I1(n3121), .I2(g109), .O(g4340) );
  NR2X1 U2062 ( .I1(n2295), .I2(n2072), .O(g4338) );
  AN2X1 U2063 ( .I1(n2955), .I2(g109), .O(g4334) );
  NR2X1 U2064 ( .I1(n2295), .I2(n1949), .O(g4330) );
  AN2X1 U2065 ( .I1(n2954), .I2(g109), .O(g4325) );
  MUX2X1 U2066 ( .A(n3116), .B(n2997), .S(n2525), .O(g4309) );
  MUX2X1 U2067 ( .A(n3066), .B(n2995), .S(n2525), .O(g4293) );
  MUX2X1 U2068 ( .A(n3077), .B(n3186), .S(n2525), .O(g4283) );
  MXL2XLP U2069 ( .A(n2014), .B(n1920), .S(n2525), .OB(g4274) );
  MXL2XLP U2070 ( .A(n2015), .B(n1874), .S(n2525), .OB(g4264) );
  MXL2XLP U2071 ( .A(n1947), .B(n1992), .S(n2525), .OB(g4255) );
  MUX2X1 U2072 ( .A(n3103), .B(n2994), .S(n2525), .O(g4239) );
  MUX2X1 U2073 ( .A(n3110), .B(n3151), .S(n2525), .O(g4238) );
  MXL2XLP U2074 ( .A(n2060), .B(n1901), .S(n2525), .OB(g4231) );
  OAI12X1 U2075 ( .B1(n3165), .B2(n1963), .A1(n2153), .O(g4117) );
  ND2X1 U2076 ( .I1(n2351), .I2(n1889), .O(n2153) );
  NR3X1 U2077 ( .I1(n3136), .I2(n2948), .I3(n3156), .O(n2351) );
  AN4B1XLP U2078 ( .I1(n3178), .I2(n3192), .I3(n3190), .B1(n2000), .O(g4114)
         );
  ND2X1 U2079 ( .I1(g1700), .I2(n1595), .O(g4089) );
  NR2X1 U2080 ( .I1(n681), .I2(n2949), .O(g4076) );
  INVCKX1 U2081 ( .I(g1700), .O(n681) );
  INVCKX1 U2082 ( .I(n2462), .O(g3524) );
  AN4B1XLP U2083 ( .I1(n3125), .I2(n3082), .I3(n3107), .B1(n1969), .O(g3506)
         );
  OAI22X1 U2084 ( .A1(n1768), .A2(n2526), .B1(n1794), .B2(n2437), .O(g3462) );
  INVCKX1 U2085 ( .I(g4171), .O(n2526) );
  MXL2XLP U2086 ( .A(n2055), .B(n1937), .S(n1870), .OB(g8566) );
  MXL2XLP U2087 ( .A(n2048), .B(n1938), .S(n1870), .OB(g6949) );
  MXL2XLP U2088 ( .A(n2049), .B(n1939), .S(n1870), .OB(g8564) );
  MXL2XLP U2089 ( .A(n2050), .B(n1940), .S(n1870), .OB(g8563) );
  AN3X1 U2090 ( .I1(g743), .I2(g109), .I3(g744), .O(g5659) );
  MXL2XLP U2091 ( .A(n2051), .B(n1941), .S(n1870), .OB(g6926) );
  AN3X1 U2092 ( .I1(g741), .I2(g109), .I3(g742), .O(g5658) );
  MXL2XLP U2093 ( .A(n2052), .B(n1942), .S(n1870), .OB(g6920) );
  AN4B1XLP U2094 ( .I1(n3092), .I2(n3124), .I3(n3162), .B1(n1979), .O(g3381)
         );
  INVCKX1 U2095 ( .I(g23), .O(g3327) );
  NR2X1 U2096 ( .I1(g750), .I2(n1794), .O(g4171) );
  NR2X1 U2097 ( .I1(n3159), .I2(g1737), .O(g2478) );
  MXL2XLP U2098 ( .A(n2527), .B(n2082), .S(n2437), .OB(g11647) );
  MXL2XLP U2099 ( .A(n2528), .B(n2529), .S(n2530), .OB(n2527) );
  NR2X1 U2100 ( .I1(n2531), .I2(n2532), .O(g11641) );
  XNR2X1 U2101 ( .I1(n3190), .I2(n2533), .O(n2531) );
  AN2B1XLP U2102 ( .I1(n3192), .B1(n2534), .O(n2533) );
  NR2X1 U2103 ( .I1(n2535), .I2(n2532), .O(g11640) );
  XOR2X1 U2104 ( .I1(n2534), .I2(n3192), .O(n2535) );
  ND2X1 U2105 ( .I1(n2536), .I2(n3178), .O(n2534) );
  NR2X1 U2106 ( .I1(n2537), .I2(n2532), .O(g11639) );
  XNR2X1 U2107 ( .I1(n3178), .I2(n2536), .O(n2537) );
  NR2X1 U2108 ( .I1(n2538), .I2(n2000), .O(n2536) );
  NR2X1 U2109 ( .I1(n2539), .I2(n2532), .O(g11636) );
  AO12X1 U2110 ( .B1(n592), .B2(n2951), .A1(n2295), .O(n2532) );
  ND2X1 U2111 ( .I1(g109), .I2(n2540), .O(n592) );
  OAI12X1 U2112 ( .B1(n3060), .B2(n3061), .A1(n3058), .O(n2540) );
  XNR2X1 U2113 ( .I1(n3163), .I2(n519), .O(n2539) );
  MXL2XLP U2114 ( .A(n2541), .B(n2040), .S(n2437), .OB(g11625) );
  XNR2X1 U2115 ( .I1(n2529), .I2(n2528), .O(n2541) );
  XNR3X1 U2116 ( .I1(n2542), .I2(n2543), .I3(n2544), .O(n2528) );
  XOR4XLP U2117 ( .I1(n2545), .I2(n2546), .I3(n2547), .I4(n2548), .O(n2543) );
  XOR4XLP U2118 ( .I1(n2549), .I2(n2550), .I3(n2551), .I4(n2552), .O(n2542) );
  MUX2X1 U2119 ( .A(n2553), .B(n1983), .S(n2554), .O(n2529) );
  XOR2X1 U2120 ( .I1(n2555), .I2(n2556), .O(n2553) );
  NR2X1 U2121 ( .I1(n3148), .I2(n2557), .O(n2555) );
  MUX2X1 U2122 ( .A(n3138), .B(n2997), .S(n2558), .O(g11610) );
  MUX2X1 U2123 ( .A(n3175), .B(n2995), .S(n2558), .O(g11609) );
  MUX2X1 U2124 ( .A(n3144), .B(n3186), .S(n2558), .O(g11608) );
  MUX2X1 U2125 ( .A(n3081), .B(n2996), .S(n2558), .O(g11607) );
  MUX2X1 U2126 ( .A(n3088), .B(n3187), .S(n2558), .O(g11606) );
  MUX2X1 U2127 ( .A(n3193), .B(n3160), .S(n2558), .O(g11605) );
  MXL2XLP U2128 ( .A(n1948), .B(n1956), .S(n2558), .OB(g11604) );
  MUX2X1 U2129 ( .A(n3180), .B(n3151), .S(n2558), .O(g11603) );
  MUX2X1 U2130 ( .A(n3135), .B(n2993), .S(n2558), .O(g11602) );
  AN2X1 U2131 ( .I1(g1317), .I2(n519), .O(n2558) );
  INVCKX1 U2132 ( .I(n2538), .O(n519) );
  OAI112X1 U2133 ( .C1(n2559), .C2(n2560), .A1(n2431), .B1(n2430), .O(n2538)
         );
  INVCKX1 U2134 ( .I(n2420), .O(n2430) );
  OR4B2XLP U2135 ( .I1(n2561), .I2(n2562), .B1(n2563), .B2(n2564), .O(n2560)
         );
  XNR2X1 U2136 ( .I1(n3010), .I2(n2983), .O(n2564) );
  NR2X1 U2137 ( .I1(n2565), .I2(n2566), .O(n2563) );
  XNR2X1 U2138 ( .I1(n1978), .I2(n3001), .O(n2566) );
  XNR2X1 U2139 ( .I1(n1877), .I2(n3009), .O(n2565) );
  XNR2X1 U2140 ( .I1(n1896), .I2(n3003), .O(n2562) );
  XNR2X1 U2141 ( .I1(n1977), .I2(n3004), .O(n2561) );
  OR4B2XLP U2142 ( .I1(n2567), .I2(n2568), .B1(n2569), .B2(n2570), .O(n2559)
         );
  NR2X1 U2143 ( .I1(n2571), .I2(n2572), .O(n2570) );
  XNR2X1 U2144 ( .I1(n1903), .I2(n3005), .O(n2572) );
  XNR2X1 U2145 ( .I1(n1879), .I2(n3006), .O(n2571) );
  XOR2X1 U2146 ( .I1(n2573), .I2(n2574), .O(n2569) );
  XNR2X1 U2147 ( .I1(n1980), .I2(n3008), .O(n2568) );
  XNR2X1 U2148 ( .I1(n1869), .I2(n3007), .O(n2567) );
  MXL2XLP U2149 ( .A(n2023), .B(n2575), .S(n2292), .OB(g11579) );
  XOR4XLP U2150 ( .I1(n2576), .I2(n3159), .I3(n2577), .I4(n2578), .O(n2575) );
  ND2X1 U2151 ( .I1(n2329), .I2(n1964), .O(n2577) );
  NR3X1 U2152 ( .I1(n3126), .I2(n2953), .I3(n1891), .O(n2329) );
  MXL2XLP U2153 ( .A(n2579), .B(n3169), .S(n3121), .OB(n2576) );
  AOI12X1 U2154 ( .B1(n2580), .B2(n2581), .A1(n3169), .O(n2579) );
  AN4B2X1 U2155 ( .I1(n1913), .I2(n2033), .B1(n2957), .B2(n2582), .O(n2581) );
  OR4B2XLP U2156 ( .I1(n2954), .I2(n2955), .B1(n2072), .B2(n1949), .O(n2582)
         );
  AN4B2X1 U2157 ( .I1(n1982), .I2(n1908), .B1(n3184), .B2(n2583), .O(n2580) );
  ND3X1 U2158 ( .I1(n2013), .I2(n1924), .I3(n1884), .O(n2583) );
  NR2X1 U2159 ( .I1(n2295), .I2(n2584), .O(g11514) );
  XOR4XLP U2160 ( .I1(n1917), .I2(n2585), .I3(n2964), .I4(n2578), .O(n2584) );
  MUX3X1 U2161 ( .A(n2586), .B(n2062), .C(n3171), .S0(n2587), .S1(g18), .O(
        n2578) );
  AN4B2X1 U2162 ( .I1(n2075), .I2(n1952), .B1(n3046), .B2(n3047), .O(n2587) );
  ND2X1 U2163 ( .I1(n2588), .I2(n2589), .O(n2586) );
  XOR2X1 U2164 ( .I1(n2961), .I2(n2962), .O(n2585) );
  MXL2XLP U2165 ( .A(n2548), .B(n2083), .S(n2437), .OB(g11488) );
  MXL2XLP U2166 ( .A(n3038), .B(n2590), .S(n2591), .OB(n2548) );
  XNR2X1 U2167 ( .I1(n1894), .I2(n2592), .O(n2590) );
  AN4B1XLP U2168 ( .I1(n3139), .I2(n3150), .I3(n1873), .B1(n3148), .O(n2592)
         );
  MXL2XLP U2169 ( .A(n2547), .B(n2084), .S(n2437), .OB(g11487) );
  MXL2XLP U2170 ( .A(n3042), .B(n2593), .S(n2591), .OB(n2547) );
  XNR2X1 U2171 ( .I1(n1876), .I2(n2594), .O(n2593) );
  NR2X1 U2172 ( .I1(n3123), .I2(n2595), .O(n2594) );
  MXL2XLP U2173 ( .A(n2546), .B(n2085), .S(n2437), .OB(g11486) );
  MXL2XLP U2174 ( .A(n2596), .B(n3045), .S(n2554), .OB(n2546) );
  XNR2X1 U2175 ( .I1(n1960), .I2(n2597), .O(n2596) );
  MXL2XLP U2176 ( .A(n2545), .B(n2086), .S(n2437), .OB(g11485) );
  MXL2XLP U2177 ( .A(n2598), .B(n3043), .S(n2554), .OB(n2545) );
  XNR2X1 U2178 ( .I1(n1868), .I2(n2599), .O(n2598) );
  NR2X1 U2179 ( .I1(n1873), .I2(n2600), .O(n2599) );
  MXL2XLP U2180 ( .A(n2552), .B(n2087), .S(n2437), .OB(g11484) );
  MXL2XLP U2181 ( .A(n3034), .B(n2601), .S(n2591), .OB(n2552) );
  XNR2X1 U2182 ( .I1(n1974), .I2(n2602), .O(n2601) );
  NR2X1 U2183 ( .I1(n2557), .I2(n1892), .O(n2602) );
  ND3X1 U2184 ( .I1(n1955), .I2(n1873), .I3(n3150), .O(n2557) );
  MXL2XLP U2185 ( .A(n2551), .B(n2088), .S(n2437), .OB(g11483) );
  MXL2XLP U2186 ( .A(n3035), .B(n2603), .S(n2591), .OB(n2551) );
  XNR2X1 U2187 ( .I1(n1898), .I2(n2604), .O(n2603) );
  NR2X1 U2188 ( .I1(n3123), .I2(n2600), .O(n2604) );
  ND3X1 U2189 ( .I1(n1872), .I2(n1955), .I3(n3148), .O(n2600) );
  MXL2XLP U2190 ( .A(n2550), .B(n2089), .S(n2437), .OB(g11482) );
  MXL2XLP U2191 ( .A(n2605), .B(n3033), .S(n2554), .OB(n2550) );
  XNR2X1 U2192 ( .I1(n1959), .I2(n2606), .O(n2605) );
  NR2X1 U2193 ( .I1(n1872), .I2(n2607), .O(n2606) );
  MXL2XLP U2194 ( .A(n2549), .B(n2090), .S(n2437), .OB(g11481) );
  MXL2XLP U2195 ( .A(n3029), .B(n2608), .S(n2591), .OB(n2549) );
  XNR2X1 U2196 ( .I1(n1897), .I2(n2609), .O(n2608) );
  NR2X1 U2197 ( .I1(n3150), .I2(n2607), .O(n2609) );
  ND3X1 U2198 ( .I1(n1892), .I2(n1955), .I3(n3123), .O(n2607) );
  MXL2XLP U2199 ( .A(n2544), .B(n2091), .S(n2437), .OB(g11478) );
  ND2X1 U2200 ( .I1(n1768), .I2(g750), .O(n2437) );
  MXL2XLP U2201 ( .A(n2610), .B(n3040), .S(n2554), .OB(n2544) );
  XNR2X1 U2202 ( .I1(n1975), .I2(n2611), .O(n2610) );
  NR2X1 U2203 ( .I1(n2595), .I2(n1873), .O(n2611) );
  ND3X1 U2204 ( .I1(n1872), .I2(n1892), .I3(n3139), .O(n2595) );
  OAI22X1 U2205 ( .A1(n2573), .A2(n2420), .B1(n1896), .B2(n2419), .O(g11443)
         );
  ND2X1 U2206 ( .I1(g109), .I2(n2420), .O(n2419) );
  ND3X1 U2207 ( .I1(n1823), .I2(n2292), .I3(n2974), .O(n2420) );
  MXL2XLP U2208 ( .A(n2574), .B(n2612), .S(n2431), .OB(n2573) );
  AN4B1XLP U2209 ( .I1(n2978), .I2(n2977), .I3(n2976), .B1(n1994), .O(n2431)
         );
  MUX2X1 U2210 ( .A(n2613), .B(n1900), .S(n2979), .O(n2612) );
  OAI13X1 U2211 ( .B1(n2614), .B2(n2615), .B3(n2616), .A1(n1900), .O(n2613) );
  ND3X1 U2212 ( .I1(n1896), .I2(n1877), .I3(n1869), .O(n2616) );
  OR4B2XLP U2213 ( .I1(n2980), .I2(n2981), .B1(n1988), .B2(n1914), .O(n2615)
         );
  OR4B2XLP U2214 ( .I1(n2985), .I2(n2986), .B1(n1879), .B2(n2617), .O(n2614)
         );
  NR3X1 U2215 ( .I1(n2984), .I2(n2982), .I3(n2983), .O(n2617) );
  XOR2X1 U2216 ( .I1(n3002), .I2(n2618), .O(n2574) );
  NR2X1 U2217 ( .I1(n2530), .I2(n2063), .O(n2618) );
  NR2X1 U2218 ( .I1(n2619), .I2(n2620), .O(g11393) );
  XNR2X1 U2219 ( .I1(n3082), .I2(n2621), .O(n2619) );
  NR2X1 U2220 ( .I1(n1969), .I2(n2622), .O(n2621) );
  NR2X1 U2221 ( .I1(n2623), .I2(n2620), .O(g11392) );
  XNR2X1 U2222 ( .I1(n2622), .I2(n1969), .O(n2623) );
  ND2X1 U2223 ( .I1(n2624), .I2(n3125), .O(n2622) );
  NR2X1 U2224 ( .I1(n2625), .I2(n2620), .O(g11391) );
  XNR2X1 U2225 ( .I1(n3125), .I2(n2624), .O(n2625) );
  AN2X1 U2226 ( .I1(n3107), .I2(n523), .O(n2624) );
  AOI12X1 U2227 ( .B1(n1955), .B2(n2626), .A1(n2627), .O(g11380) );
  OR2B1XLP U2228 ( .I1(n2628), .B1(n2597), .O(n2626) );
  AN4B1XLP U2229 ( .I1(n3148), .I2(n1955), .I3(n3123), .B1(n1872), .O(n2597)
         );
  NR2X1 U2230 ( .I1(n2629), .I2(n2627), .O(g11376) );
  XNR2X1 U2231 ( .I1(n2630), .I2(n1892), .O(n2629) );
  ND2X1 U2232 ( .I1(n2631), .I2(n3123), .O(n2630) );
  NR2X1 U2233 ( .I1(n2632), .I2(n2627), .O(g11372) );
  XNR2X1 U2234 ( .I1(n3123), .I2(n2631), .O(n2632) );
  NR2X1 U2235 ( .I1(n2628), .I2(n1872), .O(n2631) );
  NR2X1 U2236 ( .I1(n2633), .I2(n2620), .O(g11349) );
  AO12X1 U2237 ( .B1(n2634), .B2(n3000), .A1(n2295), .O(n2620) );
  XNR2X1 U2238 ( .I1(n523), .I2(n3107), .O(n2633) );
  NR2X1 U2239 ( .I1(n2635), .I2(n2627), .O(g11340) );
  ND2X1 U2240 ( .I1(g109), .I2(n1594), .O(n2627) );
  XNR2X1 U2241 ( .I1(n2628), .I2(n1872), .O(n2635) );
  ND2X1 U2242 ( .I1(n2636), .I2(n2591), .O(n2628) );
  OR4B2XLP U2243 ( .I1(n1892), .I2(n1873), .B1(n3139), .B2(n3150), .O(n2636)
         );
  MXL2XLP U2244 ( .A(n1975), .B(n1894), .S(n2591), .OB(g11338) );
  MXL2XLP U2245 ( .A(n1894), .B(n1876), .S(n2591), .OB(g11337) );
  MXL2XLP U2246 ( .A(n1876), .B(n1960), .S(n2591), .OB(g11336) );
  MXL2XLP U2247 ( .A(n1960), .B(n1868), .S(n2591), .OB(g11335) );
  MXL2XLP U2248 ( .A(n1868), .B(n1974), .S(n2591), .OB(g11334) );
  MXL2XLP U2249 ( .A(n1974), .B(n1898), .S(n2591), .OB(g11333) );
  MXL2XLP U2250 ( .A(n1898), .B(n1959), .S(n2591), .OB(g11332) );
  MXL2XLP U2251 ( .A(n1959), .B(n1897), .S(n2591), .OB(g11331) );
  MUX2X1 U2252 ( .A(n3185), .B(n3176), .S(n2554), .O(g11330) );
  MUX2X1 U2253 ( .A(n2988), .B(n3185), .S(n2554), .O(g11329) );
  MXL2XLP U2254 ( .A(n2026), .B(n1925), .S(n2591), .OB(g11328) );
  MXL2XLP U2255 ( .A(n1925), .B(n2011), .S(n2591), .OB(g11327) );
  MXL2XLP U2256 ( .A(n2011), .B(n1918), .S(n2591), .OB(g11326) );
  MXL2XLP U2257 ( .A(n1918), .B(n1975), .S(n2591), .OB(g11325) );
  MXL2XLP U2258 ( .A(n1897), .B(n2556), .S(n2591), .OB(g11324) );
  MUX2X1 U2259 ( .A(n2637), .B(n3185), .S(n3176), .O(n2556) );
  AOI12X1 U2260 ( .B1(n2638), .B2(n2639), .A1(n3185), .O(n2637) );
  AN4B2X1 U2261 ( .I1(n1959), .I2(n1897), .B1(n2990), .B2(n2640), .O(n2639) );
  OR4B2XLP U2262 ( .I1(n2987), .I2(n2989), .B1(n1918), .B2(n2026), .O(n2640)
         );
  AN4B2X1 U2263 ( .I1(n1960), .I2(n1898), .B1(n2991), .B2(n2641), .O(n2638) );
  ND3X1 U2264 ( .I1(n1894), .I2(n1876), .I3(n1868), .O(n2641) );
  NR2X1 U2265 ( .I1(n2642), .I2(n2643), .O(g11320) );
  XNR2X1 U2266 ( .I1(n2644), .I2(n3030), .O(n2642) );
  MUX2X1 U2267 ( .A(n3117), .B(n3020), .S(n2645), .O(g11314) );
  MUX2X1 U2268 ( .A(n3069), .B(n3024), .S(n2645), .O(g11312) );
  MUX2X1 U2269 ( .A(n3075), .B(n3028), .S(n2645), .O(g11310) );
  MUX2X1 U2270 ( .A(n3083), .B(n3026), .S(n2645), .O(g11308) );
  MUX2X1 U2271 ( .A(n3172), .B(n3021), .S(n2645), .O(g11306) );
  MUX2X1 U2272 ( .A(n3093), .B(n3022), .S(n2645), .O(g11305) );
  MUX2X1 U2273 ( .A(n3106), .B(n3023), .S(n2645), .O(g11303) );
  MUX2X1 U2274 ( .A(n3108), .B(n3025), .S(n2645), .O(g11300) );
  MUX2X1 U2275 ( .A(n3118), .B(n3027), .S(n2645), .O(g11298) );
  AN2X1 U2276 ( .I1(n2634), .I2(n523), .O(n2645) );
  OA112X1 U2277 ( .C1(n2646), .C2(n2647), .A1(n2591), .B1(n2648), .O(n523) );
  OR4B2XLP U2278 ( .I1(n2649), .I2(n2650), .B1(n2651), .B2(n2652), .O(n2647)
         );
  XNR2X1 U2279 ( .I1(n3035), .I2(n3036), .O(n2652) );
  NR2X1 U2280 ( .I1(n2653), .I2(n2654), .O(n2651) );
  XNR2X1 U2281 ( .I1(n1973), .I2(n3038), .O(n2654) );
  XNR2X1 U2282 ( .I1(n1875), .I2(n3034), .O(n2653) );
  XNR2X1 U2283 ( .I1(n3029), .I2(n1957), .O(n2650) );
  XNR2X1 U2284 ( .I1(n1895), .I2(n3033), .O(n2649) );
  OR4B2XLP U2285 ( .I1(n2655), .I2(n2656), .B1(n2657), .B2(n2658), .O(n2646)
         );
  NR2X1 U2286 ( .I1(n2659), .I2(n2660), .O(n2658) );
  XNR2X1 U2287 ( .I1(n1881), .I2(n3040), .O(n2660) );
  XNR2X1 U2288 ( .I1(n1902), .I2(n3042), .O(n2659) );
  XNR2X1 U2289 ( .I1(n1983), .I2(n2661), .O(n2657) );
  XNR2X1 U2290 ( .I1(n1976), .I2(n3045), .O(n2656) );
  XNR2X1 U2291 ( .I1(n1899), .I2(n3043), .O(n2655) );
  ND2X1 U2292 ( .I1(g109), .I2(n2662), .O(n2634) );
  OAI12X1 U2293 ( .B1(n3063), .B2(n3064), .A1(n3062), .O(n2662) );
  OAI12X1 U2294 ( .B1(n2663), .B2(n2130), .A1(n2664), .O(g11294) );
  MXL2XLP U2295 ( .A(n2665), .B(n2457), .S(n3142), .OB(n2664) );
  NR2X1 U2296 ( .I1(n2247), .I2(n2124), .O(n2457) );
  INVCKX1 U2297 ( .I(n2127), .O(n2124) );
  AOI13X1 U2298 ( .B1(n2131), .B2(n1890), .B3(n2145), .A1(n2127), .O(n2665) );
  ND2X1 U2299 ( .I1(n2456), .I2(n2002), .O(n2127) );
  NR2X1 U2300 ( .I1(n2461), .I2(n2992), .O(n2456) );
  INVCKX1 U2301 ( .I(n2487), .O(n2461) );
  NR2X1 U2302 ( .I1(n1970), .I2(n3137), .O(n2487) );
  INVCKX1 U2303 ( .I(n2139), .O(n2131) );
  MUXB2X1 U2304 ( .EB(n2666), .A(n2667), .B(n2668), .S(n3153), .O(n2663) );
  OAI22X1 U2305 ( .A1(n2669), .A2(n2670), .B1(n2671), .B2(n2588), .O(n2668) );
  NR2X1 U2306 ( .I1(n2672), .I2(n2673), .O(n2667) );
  AOI22X1 U2307 ( .A1(n3160), .A2(n2674), .B1(n3151), .B2(n2675), .O(n2673) );
  AOI12X1 U2308 ( .B1(n2995), .B2(n3186), .A1(n2435), .O(n2672) );
  NR2X1 U2309 ( .I1(n1920), .I2(n1874), .O(n2435) );
  AOI122X1 U2310 ( .B1(n2674), .B2(n533), .C1(n2675), .C2(n540), .A1(n1870), 
        .O(n2666) );
  MXL2XLP U2311 ( .A(n1901), .B(n2676), .S(n3153), .OB(n2675) );
  MXL2XLP U2312 ( .A(n1956), .B(n2677), .S(n3153), .OB(n2674) );
  MXL2XLP U2313 ( .A(n2678), .B(n2679), .S(n2130), .OB(g11293) );
  NR2X1 U2314 ( .I1(n2680), .I2(n2139), .O(n2679) );
  NR3X1 U2315 ( .I1(n3188), .I2(n3155), .I3(n1961), .O(n2139) );
  AOI13X1 U2316 ( .B1(n2681), .B2(n2682), .B3(g4904), .A1(n2998), .O(n2680) );
  AN2X1 U2317 ( .I1(g1850), .I2(n2462), .O(g4904) );
  AOI12X1 U2318 ( .B1(n1871), .B2(n2999), .A1(n2247), .O(n2462) );
  INVCKX1 U2319 ( .I(n2130), .O(n2247) );
  ND2X1 U2320 ( .I1(n2683), .I2(n1871), .O(n2130) );
  OR4B2XLP U2321 ( .I1(n2999), .I2(n3155), .B1(n2145), .B2(n2254), .O(n2682)
         );
  ND3X1 U2322 ( .I1(n3188), .I2(n1953), .I3(n2683), .O(n2254) );
  NR3X1 U2323 ( .I1(n3155), .I2(n2999), .I3(n3189), .O(n2683) );
  XOR2X1 U2324 ( .I1(n2684), .I2(n2685), .O(n2681) );
  MXL2XLP U2325 ( .A(n2686), .B(n2135), .S(n3142), .OB(n2685) );
  NR2X1 U2326 ( .I1(n1890), .I2(n3188), .O(n2135) );
  ND2X1 U2327 ( .I1(n2145), .I2(n1962), .O(n2686) );
  ND2X1 U2328 ( .I1(n3189), .I2(n3188), .O(n2145) );
  MXL2XLP U2329 ( .A(n2676), .B(n1993), .S(n1870), .OB(n2678) );
  AOI12X1 U2330 ( .B1(n2066), .B2(n2687), .A1(n2643), .O(g11292) );
  OR2B1XLP U2331 ( .I1(n2688), .B1(n3173), .O(n2687) );
  NR2X1 U2332 ( .I1(n2689), .I2(n2643), .O(g11291) );
  XOR2X1 U2333 ( .I1(n2688), .I2(n3173), .O(n2689) );
  ND2X1 U2334 ( .I1(n2690), .I2(n3146), .O(n2688) );
  NR2X1 U2335 ( .I1(n2691), .I2(n2643), .O(g11290) );
  OR2B1XLP U2336 ( .I1(n3000), .B1(g109), .O(n2643) );
  XNR2X1 U2337 ( .I1(n3146), .I2(n2690), .O(n2691) );
  AN2X1 U2338 ( .I1(n2644), .I2(n3030), .O(n2690) );
  NR2X1 U2339 ( .I1(n2554), .I2(n2648), .O(n2644) );
  INVCKX1 U2340 ( .I(n2591), .O(n2554) );
  MXL2XLP U2341 ( .A(n1881), .B(n1973), .S(n2591), .OB(g11270) );
  MXL2XLP U2342 ( .A(n1973), .B(n1902), .S(n2591), .OB(g11269) );
  MXL2XLP U2343 ( .A(n1902), .B(n1976), .S(n2591), .OB(g11268) );
  MXL2XLP U2344 ( .A(n1976), .B(n1899), .S(n2591), .OB(g11267) );
  MXL2XLP U2345 ( .A(n1899), .B(n1875), .S(n2591), .OB(g11266) );
  MXL2XLP U2346 ( .A(n1875), .B(n1995), .S(n2591), .OB(g11265) );
  MXL2XLP U2347 ( .A(n1995), .B(n1895), .S(n2591), .OB(g11264) );
  MXL2XLP U2348 ( .A(n1895), .B(n1957), .S(n2591), .OB(g11263) );
  MXL2XLP U2349 ( .A(n1990), .B(n1904), .S(n2591), .OB(g11262) );
  MXL2XLP U2350 ( .A(n1904), .B(n1991), .S(n2591), .OB(g11261) );
  MXL2XLP U2351 ( .A(n1991), .B(n1926), .S(n2591), .OB(g11260) );
  MXL2XLP U2352 ( .A(n1926), .B(n2012), .S(n2591), .OB(g11259) );
  MXL2XLP U2353 ( .A(n2012), .B(n1915), .S(n2591), .OB(g11258) );
  MXL2XLP U2354 ( .A(n1915), .B(n1881), .S(n2591), .OB(g11257) );
  MXL2XLP U2355 ( .A(n1957), .B(n2661), .S(n2591), .OB(g11256) );
  ND2X1 U2356 ( .I1(n2692), .I2(n2693), .O(n2591) );
  NR4XLP U2357 ( .I1(n3024), .I2(n3023), .I3(n3025), .I4(n2694), .O(n2693) );
  OR3X1 U2358 ( .I1(n3021), .I2(n3020), .I3(n3022), .O(n2694) );
  AOI112X1 U2359 ( .C1(n2695), .C2(n2696), .A1(n2697), .B1(n2295), .O(n2692)
         );
  OR3X1 U2360 ( .I1(n3027), .I2(n3026), .I3(n3028), .O(n2697) );
  AN4B1XLP U2361 ( .I1(n2588), .I2(n2670), .I3(n2669), .B1(n546), .O(n2696) );
  AN4B1XLP U2362 ( .I1(n2698), .I2(n2677), .I3(n2676), .B1(n533), .O(n2695) );
  MUX2X1 U2363 ( .A(n1983), .B(n2699), .S(n2648), .O(n2661) );
  AN4B1XLP U2364 ( .I1(n3173), .I2(n3030), .I3(n3146), .B1(n2066), .O(n2648)
         );
  MXL2XLP U2365 ( .A(n1990), .B(n2700), .S(n1904), .OB(n2699) );
  OAI13X1 U2366 ( .B1(n2701), .B2(n2702), .B3(n2703), .A1(n1990), .O(n2700) );
  ND3X1 U2367 ( .I1(n1895), .I2(n1957), .I3(n1875), .O(n2703) );
  OR4B2XLP U2368 ( .I1(n3031), .I2(n3032), .B1(n1991), .B2(n1915), .O(n2702)
         );
  OR4B2XLP U2369 ( .I1(n3041), .I2(n3044), .B1(n1899), .B2(n2704), .O(n2701)
         );
  NR3X1 U2370 ( .I1(n3039), .I2(n3036), .I3(n3037), .O(n2704) );
  MXL2XLP U2371 ( .A(n2705), .B(n2062), .S(n2485), .OB(g10936) );
  AN4B1XLP U2372 ( .I1(n2698), .I2(n2677), .I3(n2676), .B1(n2706), .O(n2705)
         );
  ND3X1 U2373 ( .I1(n2589), .I2(n533), .I3(n2684), .O(n2706) );
  MXL2XLP U2374 ( .A(n2092), .B(n2707), .S(n2292), .OB(g10898) );
  NR2X1 U2375 ( .I1(n2530), .I2(n2708), .O(n2707) );
  XOR4XLP U2376 ( .I1(n2709), .I2(n2710), .I3(n3001), .I4(n3002), .O(n2708) );
  XOR4XLP U2377 ( .I1(n3009), .I2(n3010), .I3(n3007), .I4(n3008), .O(n2710) );
  XOR4XLP U2378 ( .I1(n3005), .I2(n3006), .I3(n3003), .I4(n3004), .O(n2709) );
  AN2X1 U2379 ( .I1(n2589), .I2(n2669), .O(n2530) );
  ND3X1 U2380 ( .I1(n2104), .I2(n2108), .I3(n2105), .O(n2589) );
  AN2X1 U2381 ( .I1(n2111), .I2(g42), .O(n2105) );
  AN4B1XLP U2382 ( .I1(n2711), .I2(n2712), .I3(n2713), .B1(g48), .O(n2111) );
  MXL2XLP U2383 ( .A(n2048), .B(n2714), .S(n2292), .OB(g10866) );
  MXL2XLP U2384 ( .A(n2715), .B(n1937), .S(n2501), .OB(g10865) );
  OAI12X1 U2385 ( .B1(n533), .B2(n2295), .A1(n2716), .O(n2715) );
  MXL2XLP U2386 ( .A(n2049), .B(n2717), .S(n2292), .OB(g10864) );
  MXL2XLP U2387 ( .A(n2718), .B(n1938), .S(n2501), .OB(g10863) );
  ND2X1 U2388 ( .I1(n2719), .I2(n2720), .O(n2718) );
  OAI12X1 U2389 ( .B1(n2677), .B2(n2295), .A1(n1958), .O(n2719) );
  MXL2XLP U2390 ( .A(n2050), .B(n2721), .S(n2292), .OB(g10862) );
  MXL2XLP U2391 ( .A(n2722), .B(n1939), .S(n2501), .OB(g10861) );
  MXL2XLP U2392 ( .A(n2051), .B(n2723), .S(n2292), .OB(g10860) );
  MXL2XLP U2393 ( .A(n2724), .B(n1940), .S(n2501), .OB(g10859) );
  MXL2XLP U2394 ( .A(n2052), .B(n2725), .S(n2292), .OB(g10858) );
  MXL2XLP U2395 ( .A(n2053), .B(n2722), .S(n2292), .OB(g10855) );
  OAI122X1 U2396 ( .B1(n2396), .B2(n2720), .C1(n540), .C2(n2726), .A1(n2727), 
        .O(n2722) );
  MXL2XLP U2397 ( .A(n1880), .B(n2041), .S(n2115), .OB(n2396) );
  MXL2XLP U2398 ( .A(n2054), .B(n2724), .S(n2292), .OB(g10800) );
  MOAI1X1 U2399 ( .A1(n527), .A2(n2728), .B1(n2391), .B2(n2729), .O(n2724) );
  MXL2XLP U2400 ( .A(n3012), .B(n3011), .S(n2115), .OB(n2391) );
  MXL2XLP U2401 ( .A(n2016), .B(n2730), .S(n2292), .OB(g10799) );
  MXL2XLP U2402 ( .A(n2017), .B(n2714), .S(n2292), .OB(g10798) );
  OA22X1 U2403 ( .A1(n2684), .A2(n2726), .B1(n2394), .B2(n2720), .O(n2714) );
  AOI12X1 U2404 ( .B1(n2115), .B2(n3013), .A1(n2731), .O(n2394) );
  INVCKX1 U2405 ( .I(n2305), .O(n2731) );
  ND2X1 U2406 ( .I1(n3014), .I2(g18), .O(n2305) );
  MXL2XLP U2407 ( .A(n2018), .B(n2717), .S(n2292), .OB(g10797) );
  OA22X1 U2408 ( .A1(n2389), .A2(n2720), .B1(n2732), .B2(n2728), .O(n2717) );
  AOI12X1 U2409 ( .B1(n2115), .B2(n3015), .A1(n2733), .O(n2389) );
  INVCKX1 U2410 ( .I(n2299), .O(n2733) );
  ND2X1 U2411 ( .I1(n3016), .I2(g18), .O(n2299) );
  MXL2XLP U2412 ( .A(n2019), .B(n2721), .S(n2292), .OB(g10795) );
  OA22X1 U2413 ( .A1(n2381), .A2(n2720), .B1(n2677), .B2(n2728), .O(n2721) );
  AOI12X1 U2414 ( .B1(n2115), .B2(n3017), .A1(n2734), .O(n2381) );
  INVCKX1 U2415 ( .I(n2332), .O(n2734) );
  ND2X1 U2416 ( .I1(n3018), .I2(g18), .O(n2332) );
  MXL2XLP U2417 ( .A(n2020), .B(n2723), .S(n2292), .OB(g10793) );
  OAI22X1 U2418 ( .A1(n2377), .A2(n2720), .B1(n540), .B2(n2728), .O(n2723) );
  ND3X1 U2419 ( .I1(n2720), .I2(n1958), .I3(g109), .O(n2728) );
  OAI12X1 U2420 ( .B1(g18), .B2(n2021), .A1(n2322), .O(n2377) );
  ND2X1 U2421 ( .I1(n3120), .I2(g18), .O(n2322) );
  MXL2XLP U2422 ( .A(n2022), .B(n2725), .S(n2292), .OB(g10791) );
  AOI23X1 U2423 ( .B1(n2716), .B2(n527), .B3(g109), .A1(n2398), .A2(n2729), 
        .O(n2725) );
  OAI12X1 U2424 ( .B1(g18), .B2(n2023), .A1(n2312), .O(n2398) );
  ND2X1 U2425 ( .I1(n3019), .I2(g18), .O(n2312) );
  AN2B1XLP U2426 ( .I1(n3046), .B1(n2447), .O(g10785) );
  AN2X1 U2427 ( .I1(n3047), .I2(n2485), .O(g10784) );
  INVCKX1 U2428 ( .I(n2447), .O(n2485) );
  NR2X1 U2429 ( .I1(n2447), .I2(n1952), .O(g10782) );
  NR2X1 U2430 ( .I1(n2447), .I2(n2075), .O(g10780) );
  NR2X1 U2431 ( .I1(n2735), .I2(n3057), .O(n2447) );
  XNR2X1 U2432 ( .I1(n2736), .I2(n526), .O(g11163) );
  INVCKX1 U2433 ( .I(n2737), .O(n526) );
  MXL2XLP U2434 ( .A(n2055), .B(n2730), .S(n2292), .OB(g10776) );
  INVCKX1 U2435 ( .I(n2738), .O(n2730) );
  OAI122X1 U2436 ( .B1(n2400), .B2(n2720), .C1(n2588), .C2(n2726), .A1(n2727), 
        .O(n2738) );
  AOI12X1 U2437 ( .B1(n2115), .B2(n3048), .A1(n2739), .O(n2400) );
  INVCKX1 U2438 ( .I(n2317), .O(n2739) );
  ND2X1 U2439 ( .I1(n3049), .I2(g18), .O(n2317) );
  OAI22X1 U2440 ( .A1(n2740), .A2(n2068), .B1(n2677), .B2(n2741), .O(g10773)
         );
  OAI22X1 U2441 ( .A1(n2740), .A2(n1935), .B1(n2698), .B2(n2741), .O(g10771)
         );
  OAI22X1 U2442 ( .A1(n2740), .A2(n2069), .B1(n2676), .B2(n2741), .O(g10770)
         );
  MXL2XLP U2443 ( .A(n2742), .B(n1941), .S(n2501), .OB(g10767) );
  MXL2XLP U2444 ( .A(n2743), .B(n1942), .S(n2501), .OB(g10765) );
  ND2X1 U2445 ( .I1(n3057), .I2(n2735), .O(n2501) );
  INVCKX1 U2446 ( .I(g1696), .O(n2735) );
  MXL2XLP U2447 ( .A(n2094), .B(n2742), .S(n2292), .OB(g10718) );
  OAI122X1 U2448 ( .B1(n2744), .B2(n2720), .C1(n578), .C2(n2726), .A1(n2727), 
        .O(n2742) );
  INVCKX1 U2449 ( .I(n2383), .O(n2744) );
  MXL2XLP U2450 ( .A(n3052), .B(n3051), .S(n2115), .OB(n2383) );
  MXL2XLP U2451 ( .A(n2024), .B(n2743), .S(n2292), .OB(g10717) );
  INVCKX1 U2452 ( .I(n2745), .O(n2743) );
  OAI122X1 U2453 ( .B1(n2402), .B2(n2720), .C1(n2669), .C2(n2726), .A1(n2727), 
        .O(n2745) );
  ND2X1 U2454 ( .I1(n2716), .I2(n2295), .O(n2727) );
  INVCKX1 U2455 ( .I(n2726), .O(n2716) );
  ND2X1 U2456 ( .I1(n2720), .I2(n1958), .O(n2726) );
  INVCKX1 U2457 ( .I(n2729), .O(n2720) );
  NR2X1 U2458 ( .I1(n3055), .I2(n3134), .O(n2729) );
  AOI12X1 U2459 ( .B1(n2115), .B2(n3053), .A1(n2746), .O(n2402) );
  INVCKX1 U2460 ( .I(n2327), .O(n2746) );
  ND2X1 U2461 ( .I1(n3054), .I2(g18), .O(n2327) );
  INVCKX1 U2462 ( .I(g18), .O(n2115) );
  ND2X1 U2463 ( .I1(n2747), .I2(n2737), .O(g10801) );
  XOR4XLP U2464 ( .I1(n541), .I2(n2732), .I3(n2671), .I4(n2748), .O(n2737) );
  XOR4XLP U2465 ( .I1(n547), .I2(n578), .I3(n527), .I4(n2749), .O(n2748) );
  XNR3X1 U2466 ( .I1(n552), .I2(n540), .I3(n2750), .O(n2749) );
  ND2X1 U2467 ( .I1(n3056), .I2(n2751), .O(n2750) );
  INVCKX1 U2468 ( .I(n2588), .O(n552) );
  INVCKX1 U2469 ( .I(n2669), .O(n547) );
  INVCKX1 U2470 ( .I(n2677), .O(n541) );
  MXL2XLP U2471 ( .A(n2071), .B(n2684), .S(n2740), .OB(g10711) );
  NR2X1 U2472 ( .I1(n2295), .I2(n546), .O(n2684) );
  INVCKX1 U2473 ( .I(n2671), .O(n546) );
  OAI22X1 U2474 ( .A1(n2740), .A2(n1950), .B1(n2732), .B2(n2741), .O(g10707)
         );
  ND2X1 U2475 ( .I1(n2740), .I2(g109), .O(n2741) );
  AN2X1 U2476 ( .I1(n3057), .I2(g1696), .O(n2740) );
  INVCKX1 U2477 ( .I(n2752), .O(g10628) );
  NR2X1 U2478 ( .I1(n2736), .I2(n2752), .O(g11206) );
  OAI22X1 U2479 ( .A1(n2677), .A2(n2373), .B1(n2753), .B2(n2295), .O(n2752) );
  AOI122X1 U2480 ( .B1(g881), .B2(n540), .C1(g877), .C2(n527), .A1(n2754), .O(
        n2753) );
  OAI23X1 U2481 ( .B1(n2671), .B2(n3063), .B3(n3064), .A1(n3062), .A2(n2732), 
        .O(n2754) );
  INVCKX1 U2482 ( .I(n2676), .O(n527) );
  INVCKX1 U2483 ( .I(n2698), .O(n540) );
  ND3X1 U2484 ( .I1(g2986), .I2(n1834), .I3(g109), .O(n2373) );
  OAI22X1 U2485 ( .A1(n2669), .A2(n2523), .B1(n2755), .B2(n2295), .O(n2736) );
  AOI122X1 U2486 ( .B1(n533), .B2(n2080), .C1(n578), .C2(g2648), .A1(n2756), 
        .O(n2755) );
  OAI23X1 U2487 ( .B1(n2671), .B2(n3060), .B3(n3061), .A1(n3059), .A2(n2588), 
        .O(n2756) );
  INVCKX1 U2488 ( .I(n2670), .O(n578) );
  INVCKX1 U2489 ( .I(n2732), .O(n533) );
  ND2X1 U2490 ( .I1(n2525), .I2(g109), .O(n2523) );
  AN2X1 U2491 ( .I1(n3159), .I2(g1765), .O(n2525) );
  ND2X1 U2492 ( .I1(n2747), .I2(n2588), .O(g10465) );
  AN4B2X1 U2493 ( .I1(n2757), .I2(n2758), .B1(n2759), .B2(n2760), .O(n2588) );
  OAI122X1 U2494 ( .B1(n2761), .B2(n1929), .C1(n2762), .C2(n2056), .A1(n2763), 
        .O(n2760) );
  AOI23X1 U2495 ( .B1(n2764), .B2(n2765), .B3(n2766), .A1(n3069), .A2(n2767), 
        .O(n2763) );
  AO222X1 U2496 ( .A1(n2768), .A2(n3070), .B1(n2769), .B2(n3066), .C1(n2770), 
        .C2(n3071), .O(n2759) );
  AOI222X1 U2497 ( .A1(n3067), .A2(n2771), .B1(n3068), .B2(n2751), .C1(n3065), 
        .C2(n2772), .O(n2758) );
  AOI222X1 U2498 ( .A1(g1185), .A2(n2773), .B1(g913), .B2(n2774), .C1(n3175), 
        .C2(n2775), .O(n2757) );
  ND2X1 U2499 ( .I1(n2747), .I2(n2671), .O(g10463) );
  AN4B2X1 U2500 ( .I1(n2776), .I2(n2777), .B1(n2778), .B2(n2779), .O(n2671) );
  OAI122X1 U2501 ( .B1(n2780), .B2(n1930), .C1(n2761), .C2(n2057), .A1(n2781), 
        .O(n2779) );
  AOI22X1 U2502 ( .A1(n3074), .A2(n2772), .B1(n3073), .B2(n2770), .O(n2781) );
  OAI122X1 U2503 ( .B1(n2782), .B2(n2081), .C1(n2783), .C2(n1945), .A1(n2784), 
        .O(n2778) );
  MAOI1X1 U2504 ( .A1(n3077), .A2(n2769), .B1(n2071), .B2(n2785), .O(n2784) );
  AOI122X1 U2505 ( .B1(n3072), .B2(n2786), .C1(g910), .C2(n2774), .A1(n2787), 
        .O(n2777) );
  MOAI1X1 U2506 ( .A1(n2788), .A2(n1448), .B1(n2775), .B2(n3144), .O(n2787) );
  AOI122X1 U2507 ( .B1(g1182), .B2(n2773), .C1(n2789), .C2(g16), .A1(n2790), 
        .O(n2776) );
  MXL2XLP U2508 ( .A(n2791), .B(n3076), .S(n2792), .OB(n2790) );
  OR4B2XLP U2509 ( .I1(n2789), .I2(n2793), .B1(n2766), .B2(n2764), .O(n2791)
         );
  ND2X1 U2510 ( .I1(n2747), .I2(n2732), .O(g10461) );
  AN4B2X1 U2511 ( .I1(n2794), .I2(n2795), .B1(n2796), .B2(n2797), .O(n2732) );
  OR4B2XLP U2512 ( .I1(n2798), .I2(n2799), .B1(n2800), .B2(n2801), .O(n2797)
         );
  AOI222X1 U2513 ( .A1(g907), .A2(n2774), .B1(n3082), .B2(n2802), .C1(n3083), 
        .C2(n2767), .O(n2801) );
  AOI22X1 U2514 ( .A1(n3124), .A2(n2803), .B1(g895), .B2(n2804), .O(n2800) );
  OAI22X1 U2515 ( .A1(n2788), .A2(n1417), .B1(n2805), .B2(n2014), .O(n2799) );
  OAI222X1 U2516 ( .A1(n2780), .A2(n2097), .B1(n2806), .B2(n1886), .C1(n2785), 
        .C2(n1950), .O(n2798) );
  OAI122X1 U2517 ( .B1(n2783), .B2(n1931), .C1(n2807), .C2(n2058), .A1(n2808), 
        .O(n2796) );
  AOI222X1 U2518 ( .A1(n3079), .A2(n2786), .B1(n2789), .B2(g17), .C1(n3080), 
        .C2(n2809), .O(n2808) );
  AOI122X1 U2519 ( .B1(g1203), .B2(n2810), .C1(n2792), .C2(g8), .A1(n2811), 
        .O(n2795) );
  AOI222X1 U2520 ( .A1(g1179), .A2(n2773), .B1(n3081), .B2(n2775), .C1(n3190), 
        .C2(n2812), .O(n2794) );
  ND2X1 U2521 ( .I1(n2747), .I2(n2677), .O(g10459) );
  AN4B2X1 U2522 ( .I1(n2813), .I2(n2814), .B1(n2815), .B2(n2816), .O(n2677) );
  OR4B2XLP U2523 ( .I1(n2817), .I2(n2818), .B1(n2819), .B2(n2820), .O(n2816)
         );
  AOI222X1 U2524 ( .A1(g904), .A2(n2774), .B1(n3128), .B2(n2802), .C1(n3172), 
        .C2(n2767), .O(n2820) );
  AOI22X1 U2525 ( .A1(n3162), .A2(n2803), .B1(g892), .B2(n2804), .O(n2819) );
  OAI22X1 U2526 ( .A1(n2788), .A2(n1500), .B1(n2805), .B2(n2015), .O(n2818) );
  OAI222X1 U2527 ( .A1(n2780), .A2(n1946), .B1(n2806), .B2(n1887), .C1(n2785), 
        .C2(n2068), .O(n2817) );
  OAI122X1 U2528 ( .B1(n2783), .B2(n1932), .C1(n2807), .C2(n2096), .A1(n2821), 
        .O(n2815) );
  AOI222X1 U2529 ( .A1(n3085), .A2(n2786), .B1(n3084), .B2(n2789), .C1(n3086), 
        .C2(n2809), .O(n2821) );
  AOI122X1 U2530 ( .B1(g1200), .B2(n2810), .C1(n3191), .C2(n2792), .A1(n2811), 
        .O(n2814) );
  AOI222X1 U2531 ( .A1(g1176), .A2(n2773), .B1(n3088), .B2(n2775), .C1(n3192), 
        .C2(n2812), .O(n2813) );
  ND2X1 U2532 ( .I1(n2747), .I2(n2698), .O(g10457) );
  AN4B2X1 U2533 ( .I1(n2822), .I2(n2823), .B1(n2824), .B2(n2825), .O(n2698) );
  OAI122X1 U2534 ( .B1(n2785), .B2(n1935), .C1(n2806), .C2(n2059), .A1(n2826), 
        .O(n2825) );
  AOI222X1 U2535 ( .A1(n3091), .A2(n2789), .B1(n3093), .B2(n2767), .C1(n3090), 
        .C2(n2792), .O(n2826) );
  AO222X1 U2536 ( .A1(n2803), .A2(n3092), .B1(n2770), .B2(n3096), .C1(n2802), 
        .C2(n3125), .O(n2824) );
  AN4B1XLP U2537 ( .I1(n2827), .I2(n2828), .I3(n2829), .B1(n2830), .O(n2823)
         );
  OAI222X1 U2538 ( .A1(n2805), .A2(n1947), .B1(n2780), .B2(n2079), .C1(n2788), 
        .C2(n3094), .O(n2830) );
  AOI222X1 U2539 ( .A1(n3178), .A2(n2812), .B1(n3182), .B2(n2786), .C1(g1173), 
        .C2(n2773), .O(n2829) );
  AOI222X1 U2540 ( .A1(g925), .A2(n2831), .B1(g901), .B2(n2774), .C1(g1197), 
        .C2(n2810), .O(n2828) );
  AOI22X1 U2541 ( .A1(g889), .A2(n2804), .B1(n3193), .B2(n2775), .O(n2827) );
  AOI122X1 U2542 ( .B1(n3097), .B2(n2768), .C1(n3095), .C2(n2809), .A1(n2811), 
        .O(n2822) );
  ND2X1 U2543 ( .I1(n2747), .I2(n2676), .O(g10455) );
  AN4B2X1 U2544 ( .I1(n2832), .I2(n2833), .B1(n2834), .B2(n2835), .O(n2676) );
  OR4B2XLP U2545 ( .I1(n2836), .I2(n2837), .B1(n2838), .B2(n2839), .O(n2835)
         );
  AOI112X1 U2546 ( .C1(n3102), .C2(n2772), .A1(n2793), .B1(n2811), .O(n2839)
         );
  AN4B2X1 U2547 ( .I1(n2840), .I2(n2841), .B1(n2792), .B2(n2842), .O(n2811) );
  ND2X1 U2548 ( .I1(n2843), .I2(n2765), .O(n2842) );
  AOI222X1 U2549 ( .A1(n3101), .A2(n2809), .B1(n3104), .B2(n2771), .C1(n3103), 
        .C2(n2769), .O(n2838) );
  OAI222X1 U2550 ( .A1(n2844), .A2(n1948), .B1(n2788), .B2(n1431), .C1(n2785), 
        .C2(n2069), .O(n2837) );
  AO222X1 U2551 ( .A1(n2768), .A2(n3099), .B1(n2786), .B2(n3098), .C1(n2770), 
        .C2(n3100), .O(n2836) );
  INVCKX1 U2552 ( .I(n2807), .O(n2770) );
  OAI112X1 U2553 ( .C1(n2845), .C2(n1979), .A1(n2846), .B1(n2847), .O(n2834)
         );
  AOI222X1 U2554 ( .A1(g898), .A2(n2774), .B1(g1170), .B2(n2773), .C1(n3163), 
        .C2(n2812), .O(n2847) );
  AOI22X1 U2555 ( .A1(g1194), .A2(n2810), .B1(n3106), .B2(n2767), .O(n2846) );
  INVCKX1 U2556 ( .I(n2843), .O(n2810) );
  ND2X1 U2557 ( .I1(n2848), .I2(n2849), .O(n2843) );
  AOI222X1 U2558 ( .A1(g922), .A2(n2831), .B1(n3107), .B2(n2802), .C1(n3167), 
        .C2(n2789), .O(n2833) );
  INVCKX1 U2559 ( .I(n2840), .O(n2789) );
  ND2X1 U2560 ( .I1(n2850), .I2(n2110), .O(n2840) );
  INVCKX1 U2561 ( .I(n2851), .O(n2831) );
  AOI22X1 U2562 ( .A1(g886), .A2(n2804), .B1(n3105), .B2(n2792), .O(n2832) );
  AN2X1 U2563 ( .I1(n2850), .I2(g42), .O(n2792) );
  AN3B2X1 U2564 ( .I1(n2852), .B1(n2853), .B2(g44), .O(n2850) );
  ND2X1 U2565 ( .I1(n2747), .I2(n2670), .O(g10379) );
  AN4B2X1 U2566 ( .I1(n2854), .I2(n2855), .B1(n2856), .B2(n2857), .O(n2670) );
  AO22X1 U2567 ( .A1(n2786), .A2(n3112), .B1(n2809), .B2(n3111), .O(n2857) );
  AO222X1 U2568 ( .A1(n2768), .A2(n3109), .B1(n2751), .B2(n2098), .C1(n2802), 
        .C2(n3108), .O(n2856) );
  INVCKX1 U2569 ( .I(n2783), .O(n2768) );
  AOI22X1 U2570 ( .A1(g919), .A2(n2774), .B1(n3180), .B2(n2812), .O(n2855) );
  AOI12X1 U2571 ( .B1(g1191), .B2(n2773), .A1(n2858), .O(n2854) );
  MXL2XLP U2572 ( .A(n2095), .B(n2859), .S(n2785), .OB(n2858) );
  OR4B2XLP U2573 ( .I1(n2812), .I2(n2773), .B1(n2765), .B2(n2860), .O(n2859)
         );
  INVCKX1 U2574 ( .I(n2793), .O(n2765) );
  AN4B2X1 U2575 ( .I1(n2107), .I2(n2861), .B1(n2862), .B2(n2106), .O(n2793) );
  NR2X1 U2576 ( .I1(n2863), .I2(n2108), .O(n2861) );
  ND2X1 U2577 ( .I1(n2747), .I2(n2669), .O(g10377) );
  AN4B2X1 U2578 ( .I1(n2864), .I2(n2865), .B1(n2866), .B2(n2867), .O(n2669) );
  AO222X1 U2579 ( .A1(n2809), .A2(n3114), .B1(n2769), .B2(n3116), .C1(n2786), 
        .C2(n3115), .O(n2867) );
  INVCKX1 U2580 ( .I(n2762), .O(n2786) );
  ND2X1 U2581 ( .I1(n2806), .I2(n2868), .O(n2762) );
  INVCKX1 U2582 ( .I(n2805), .O(n2769) );
  INVCKX1 U2583 ( .I(n2761), .O(n2809) );
  ND2X1 U2584 ( .I1(n2780), .I2(n2869), .O(n2761) );
  OAI122X1 U2585 ( .B1(n2783), .B2(n1933), .C1(n2785), .C2(n2060), .A1(n2870), 
        .O(n2866) );
  AOI22X1 U2586 ( .A1(n3118), .A2(n2802), .B1(n3117), .B2(n2767), .O(n2870) );
  ND2X1 U2587 ( .I1(n2871), .I2(n2807), .O(n2783) );
  ND2X1 U2588 ( .I1(n2871), .I2(n2110), .O(n2807) );
  AOI222X1 U2589 ( .A1(g1188), .A2(n2773), .B1(n3113), .B2(n2751), .C1(n3138), 
        .C2(n2775), .O(n2865) );
  AOI122X1 U2590 ( .B1(g916), .B2(n2774), .C1(n3135), .C2(n2812), .A1(n2841), 
        .O(n2864) );
  AN3X1 U2591 ( .I1(n2764), .I2(n2872), .I3(n2766), .O(n2841) );
  NR2X1 U2592 ( .I1(n2775), .I2(n2773), .O(n2766) );
  AN2B1XLP U2593 ( .I1(n2848), .B1(n2873), .O(n2773) );
  INVCKX1 U2594 ( .I(n2844), .O(n2775) );
  ND2X1 U2595 ( .I1(n2848), .I2(n2874), .O(n2844) );
  AN3X1 U2596 ( .I1(n2805), .I2(n2785), .I3(n2860), .O(n2764) );
  AN4B2X1 U2597 ( .I1(n2875), .I2(n2876), .B1(n2868), .B2(n2869), .O(n2860) );
  OAI12X1 U2598 ( .B1(n2853), .B2(n2877), .A1(n2780), .O(n2869) );
  INVCKX1 U2599 ( .I(n2771), .O(n2780) );
  AN2B1XLP U2600 ( .I1(n2874), .B1(n2853), .O(n2771) );
  OAI12X1 U2601 ( .B1(n2853), .B2(n2873), .A1(n2806), .O(n2868) );
  INVCKX1 U2602 ( .I(n2772), .O(n2806) );
  NR2X1 U2603 ( .I1(n2863), .I2(n2853), .O(n2772) );
  AN4B2X1 U2604 ( .I1(n2851), .I2(n2878), .B1(n2804), .B2(n2871), .O(n2876) );
  AN4B1XLP U2605 ( .I1(n2713), .I2(n2712), .I3(g44), .B1(n2853), .O(n2871) );
  ND3X1 U2606 ( .I1(n2879), .I2(n2108), .I3(n2104), .O(n2853) );
  INVCKX1 U2607 ( .I(g47), .O(n2108) );
  AN4B1XLP U2608 ( .I1(n2880), .I2(n2881), .I3(g45), .B1(n2712), .O(n2804) );
  NR2X1 U2609 ( .I1(g44), .I2(n2110), .O(n2881) );
  NR2X1 U2610 ( .I1(n2774), .I2(n2767), .O(n2878) );
  INVCKX1 U2611 ( .I(n2782), .O(n2767) );
  ND2X1 U2612 ( .I1(n2874), .I2(n2880), .O(n2782) );
  AN4B1XLP U2613 ( .I1(n2110), .I2(n2711), .I3(g45), .B1(g43), .O(n2874) );
  ND2X1 U2614 ( .I1(n2849), .I2(n2880), .O(n2851) );
  INVCKX1 U2615 ( .I(n2863), .O(n2849) );
  ND3X1 U2616 ( .I1(g44), .I2(n2110), .I3(n2852), .O(n2863) );
  NR3X1 U2617 ( .I1(n2751), .I2(n2802), .I3(n2803), .O(n2875) );
  INVCKX1 U2618 ( .I(n2845), .O(n2803) );
  ND3X1 U2619 ( .I1(n2882), .I2(g44), .I3(n2880), .O(n2845) );
  AN2B1XLP U2620 ( .I1(n2880), .B1(n2877), .O(n2802) );
  ND2X1 U2621 ( .I1(n2883), .I2(g42), .O(n2785) );
  ND2X1 U2622 ( .I1(n2883), .I2(n2110), .O(n2805) );
  AN4B1XLP U2623 ( .I1(g44), .I2(g45), .I3(n2848), .B1(n2712), .O(n2883) );
  INVCKX1 U2624 ( .I(n2872), .O(n2812) );
  OR2B1XLP U2625 ( .I1(n2877), .B1(n2848), .O(n2872) );
  AN3X1 U2626 ( .I1(n2104), .I2(n2879), .I3(g47), .O(n2848) );
  AN2X1 U2627 ( .I1(n2107), .I2(n2106), .O(n2104) );
  INVCKX1 U2628 ( .I(g46), .O(n2106) );
  ND2X1 U2629 ( .I1(n2882), .I2(n2711), .O(n2877) );
  INVCKX1 U2630 ( .I(g44), .O(n2711) );
  NR3X1 U2631 ( .I1(n2110), .I2(g43), .I3(n2713), .O(n2882) );
  INVCKX1 U2632 ( .I(g45), .O(n2713) );
  INVCKX1 U2633 ( .I(g42), .O(n2110) );
  AN2B1XLP U2634 ( .I1(n2880), .B1(n2873), .O(n2774) );
  ND3X1 U2635 ( .I1(g42), .I2(g44), .I3(n2852), .O(n2873) );
  NR2X1 U2636 ( .I1(n2712), .I2(g45), .O(n2852) );
  INVCKX1 U2637 ( .I(g43), .O(n2712) );
  AN4B1XLP U2638 ( .I1(n2879), .I2(g46), .I3(n2107), .B1(g47), .O(n2880) );
  OAI23X1 U2639 ( .B1(g30), .B2(g48), .B3(g41), .A1(n2751), .A2(n2862), .O(
        n2107) );
  INVCKX1 U2640 ( .I(n2879), .O(n2862) );
  NR2X1 U2641 ( .I1(n2884), .I2(g41), .O(n2879) );
  NR2X1 U2642 ( .I1(n2751), .I2(g30), .O(n2747) );
  INVCKX1 U2643 ( .I(n2788), .O(n2751) );
  NR2X1 U2644 ( .I1(n2884), .I2(g31), .O(n2788) );
  INVCKX1 U2645 ( .I(g48), .O(n2884) );
endmodule

