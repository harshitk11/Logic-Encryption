module s15850(clk, g18, g27, g109, g741, g742, g743, g744, g872, g873, g877, g881, g1712, g1960, g1961, g1696, g750, g85, g42, g1700, g102, g104, g101, g29, g28, g103, g83, g23, g87, g922, g892, g84, g919, g1182, g925, g48, g895, g889, g1185, g41, g43, g99, g1173, g1203, g1188, g1197, g46, g31, g45, g92, g89, g898, g91, g93, g913, g82, g88, g1194, g47, g96, g910, g95, g904, g1176, g901, g44, g916, g100, g886, g30, g86, g1170, g1200, g1191, g907, g90, g94, g1179, g2355, g2601, g2602, g2603, g2604, g2605, g2606, g2607, g2608, g2609, g2610, g2611, g2612, g2648, g2986, g3007, g3069, g4172, g4173, g4174, g4175, g4176, g4177, g4178, g4179, g4180, g4181, g4887, g4888, g5101, g5105, g5658, g5659, g5816, g6920, g6926, g6932, g6942, g6949, g6955, g7744, g8061, g8062, g8271, g8313, g8316, g8318, g8323, g8328, g8331, g8335, g8340, g8347, g8349, g8352, g8561, g8562, g8563, g8564, g8565, g8566, g8976, g8977, g8978, g8979, g8980, g8981, g8982, g8983, g8984, g8985, g8986, g9451, g9961, g10377, g10379, g10455, g10457, g10459, g10461, g10463, g10465, g10628, g10801, g11163, g11206, g11489, g6842, g4171, g6267, g6257, g1957, g6282, g6284, g6281, g6253, g6285, g6283, g6265, g3327, g6269, g4204, g4193, g6266, g4203, g4212, g4196, g6263, g4194, g4192, g4213, g6256, g6258, g6279, g4209, g4208, g4214, g4206, g6261, g6255, g6260, g6274, g6271, g4195, g6273, g6275, g4201, g6264, g6270, g4216, g6262, g6278, g4200, g6277, g4198, g4210, g4197, g6259, g4202, g6280, g4191, g6254, g6268, g4205, g4207, g4215, g4199, g6272, g6276, g4211);
input clk, g18, g27, g109, g741, g742, g743, g744, g872, g873, g877, g881, g1712, g1960, g1961, g1696, g750, g85, g42, g1700, g102, g104, g101, g29, g28, g103, g83, g23, g87, g922, g892, g84, g919, g1182, g925, g48, g895, g889, g1185, g41, g43, g99, g1173, g1203, g1188, g1197, g46, g31, g45, g92, g89, g898, g91, g93, g913, g82, g88, g1194, g47, g96, g910, g95, g904, g1176, g901, g44, g916, g100, g886, g30, g86, g1170, g1200, g1191, g907, g90, g94, g1179;
output g2355, g2601, g2602, g2603, g2604, g2605, g2606, g2607, g2608, g2609, g2610, g2611, g2612, g2648, g2986, g3007, g3069, g4172, g4173, g4174, g4175, g4176, g4177, g4178, g4179, g4180, g4181, g4887, g4888, g5101, g5105, g5658, g5659, g5816, g6920, g6926, g6932, g6942, g6949, g6955, g7744, g8061, g8062, g8271, g8313, g8316, g8318, g8323, g8328, g8331, g8335, g8340, g8347, g8349, g8352, g8561, g8562, g8563, g8564, g8565, g8566, g8976, g8977, g8978, g8979, g8980, g8981, g8982, g8983, g8984, g8985, g8986, g9451, g9961, g10377, g10379, g10455, g10457, g10459, g10461, g10463, g10465, g10628, g10801, g11163, g11206, g11489, g6842, g4171, g6267, g6257, g1957, g6282, g6284, g6281, g6253, g6285, g6283, g6265, g3327, g6269, g4204, g4193, g6266, g4203, g4212, g4196, g6263, g4194, g4192, g4213, g6256, g6258, g6279, g4209, g4208, g4214, g4206, g6261, g6255, g6260, g6274, g6271, g4195, g6273, g6275, g4201, g6264, g6270, g4216, g6262, g6278, g4200, g6277, g4198, g4210, g4197, g6259, g4202, g6280, g4191, g6254, g6268, g4205, g4207, g4215, g4199, g6272, g6276, g4211;
wire clk, g18, g27, g109, g741, g742, g743, g744, g872, g873, g877, g881, g1712, g1960, g1961, g1696, g750, g85, g42, g1700, g102, g104, g101, g29, g28, g103, g83, g23, g87, g922, g892, g84, g919, g1182, g925, g48, g895, g889, g1185, g41, g43, g99, g1173, g1203, g1188, g1197, g46, g31, g45, g92, g89, g898, g91, g93, g913, g82, g88, g1194, g47, g96, g910, g95, g904, g1176, g901, g44, g916, g100, g886, g30, g86, g1170, g1200, g1191, g907, g90, g94, g1179;
wire g1289, g1882, g312, g452, g123, g207, g713, g1153, g1209, g1744, g1558;
wire g695, g461, g940, g976, g709, g1092, g1574, g1864, g369, g1580, g1736;
wire g39, g1651, g1424, g1737, g1672, g1077, g1231, g4, g774, g1104, g1304;
wire g243, g1499, g1044, g1444, g757, g786, g1543, g552, g315, g1534, g622;
wire g1927, g1660, g278, g1436, g718, g76, g554, g496, g981, g878, g590;
wire g829, g1095, g704, g1265, g1786, g682, g1296, g587, g52, g646, g327;
wire g1389, g1371, g1956, g1675, g354, g113, g639, g1684, g1639, g1791, g248;
wire g1707, g1759, g351, g1957, g1604, g1098, g932, g126, g1896, g736, g1019;
wire g1362, g745, g1419, g58, g32, g876, g1086, g1486, g1730, g1504, g1470;
wire g822, g583, g1678, g174, g1766, g1801, g186, g959, g1169, g1007, g1407;
wire g1059, g1868, g758, g1718, g396, g1015, g38, g632, g1415, g1227, g1721;
wire g882, g16, g284, g426, g219, g1216, g806, g1428, g579, g1564, g1741;
wire g225, g281, g1308, g611, g631, g1217, g1589, g1466, g1571, g1861, g1365;
wire g1448, g1711, g1133, g1333, g153, g962, g766, g588, g486, g471, g1397;
wire g580, g1950, g756, g635, g1101, g549, g1041, g105, g1669, g1368, g1531;
wire g1458, g572, g1011, g33, g1411, g1074, g444, g1474, g1080, g1713, g333;
wire g269, g401, g1857, g9, g664, g965, g1400, g309, g814, g231, g557;
wire g586, g869, g1383, g158, g627, g1023, g259, g1361, g1327, g654, g293;
wire g1346, g1633, g1753, g1508, g1240, g538, g416, g542, g1681, g374, g563;
wire g1914, g530, g575, g1936, g55, g1117, g1317, g357, g386, g1601, g553;
wire g166, g501, g262, g1840, g70, g318, g1356, g794, g36, g302, g342;
wire g1250, g1163, g1810, g1032, g1432, g1053, g1453, g363, g330, g1157, g1357;
wire g35, g928, g261, g516, g254, g778, g861, g1627, g1292, g290, g1850;
wire g770, g1583, g466, g1561, g1527, g1546, g287, g560, g617, g17, g336;
wire g456, g305, g345, g8, g1771, g865, g255, g1945, g1738, g1478, g1035;
wire g1959, g1690, g1482, g1110, g296, g1663, g700, g1762, g360, g192, g1657;
wire g722, g61, g566, g1394, g1089, g883, g1071, g986, g971, g1955, g143;
wire g1814, g1038, g1212, g1918, g782, g1822, g237, g746, g1062, g1462, g178;
wire g366, g837, g599, g1854, g944, g1941, g170, g1520, g686, g953, g1958;
wire g40, g1765, g1733, g1270, g1610, g1796, g1324, g1540, g1377, g1206, g491;
wire g1849, g213, g1781, g1900, g1245, g108, g630, g148, g833, g1923, g936;
wire g1215, g1314, g849, g1336, g272, g1806, g826, g1065, g1887, g37, g968;
wire g1845, g1137, g1891, g1255, g257, g874, g591, g731, g636, g1218, g605;
wire g79, g182, g950, g1129, g857, g448, g1828, g1727, g1592, g1703, g1932;
wire g1624, g26, g1068, g578, g440, g476, g119, g668, g139, g1149, g34;
wire g1848, g263, g818, g1747, g802, g275, g1524, g1577, g810, g391, g658;
wire g1386, g253, g875, g1125, g201, g1280, g1083, g650, g1636, g853, g421;
wire g762, g956, g378, g1756, g589, g841, g1027, g1003, g1403, g1145, g1107;
wire g1223, g406, g1811, g1642, g1047, g1654, g197, g1595, g1537, g727, g999;
wire g798, g481, g754, g1330, g845, g790, g1512, g114, g1490, g1166, g1056;
wire g348, g868, g1260, g260, g131, g7, g258, g521, g1318, g1872, g677;
wire g582, g1393, g1549, g947, g1834, g1598, g1121, g1321, g506, g546, g1909;
wire g755, g1552, g584, g1687, g1586, g324, g1141, g1570, g1341, g1710, g1645;
wire g115, g135, g525, g581, g1607, g321, g67, g1275, g1311, g1615, g382;
wire g1374, g266, g1284, g1380, g673, g1853, g162, g411, g431, g1905, g1515;
wire g1630, g49, g991, g1300, g339, g256, g1750, g585, g1440, g1666, g1528;
wire g1351, g1648, g127, g1618, g1235, g299, g435, g64, g1555, g995, g1621;
wire g1113, g643, g1494, g1567, g691, g534, g1776, g569, g1160, g1360, g1050;
wire g1, g511, g1724, g12, g1878, g73, I8854, g5652, I12913, g11354, g6837;
wire I10941, I6979, g5843, g2771, g3537, g6062, I9984, I14382, g7706, I13618, I15181;
wire g6620, I12436, g5193, g6462, g8925, I14519, g10289, I14176, I14185, g11181, I14675;
wire g2299, I12607, g3272, g2547, g9291, I6001, I7048, g10309, g7029, g4440, I9544;
wire g10288, I12274, I9483, g7787, I6676, I8520, g10571, I17692, I17761, I13469, g9344;
wire g7956, g3417, g4323, I11286, I8031, g7675, g8320, I12565, I16644, I11306, g1981;
wire I7333, I13039, g3982, g6249, g9259, I15190, g11426, g9819, g8277, I5050, I5641;
wire g5121, g1997, g3629, g3328, I12641, g5670, g6842, g8617, I15520, I7396, I7803;
wire g3330, g2991, I9461, g2244, g6192, g6298, g6085, I12153, g4351, I11677, g10687;
wire g4530, g8516, g5232, I13975, g2078, I8911, g2340, g7684, I12409, g7745, g8987;
wire g11546, I10729, g5253, g7338, I7509, I9427, g3800, I15088, g2907, g7791, I11143;
wire g6854, g11088, g7309, g8299, I9046, g6941, g2435, I14439, g4010, g2082, I6932;
wire I7662, I9446, g5519, g5740, I5289, I9514, g7808, g2482, I5658, I15497, I6624;
wire g8892, I11169, g3213, I6068, g11497, I13791, I16867, I10349, g10260, g7759, I8473;
wire I14349, g6708, g10668, I5271, I9191, I9391, g6219, I15250, I17100, I14906, g9825;
wire g7201, I14083, g10195, I8324, g6031, g2915, I13666, I9695, I11363, I11217, g6431;
wire g6252, g4172, g6812, g8991, g4372, g7049, I6576, g10525, g10488, I10566, I13478;
wire g5586, g8709, g2214, I9536, g6176, g4618, I15296, g4143, I7381, I9159, g11339;
wire g8140, I16979, I16496, g8078, I7847, I9359, g8340, g2110, I15338, g6405, g8478;
wire I16111, g4282, g11644, g7604, g9768, g4566, g7098, g10893, I4961, g4988, g6286;
wire g8959, I13580, I9016, I6398, g8517, g3348, I15060, I15968, I5332, g8482, g2002;
wire I10138, g11060, I17407, I12303, g5645, I15855, g2824, g11197, g4555, g5691, I9642;
wire g7539, g7896, g8656, g9887, I8199, g6974, g6270, I14415, g3260, g11411, I10852;
wire g10042, g10255, g6073, g10189, I4903, g2877, I11531, g10679, g6796, I8900, I16735;
wire g1968, g5879, I10963, g10270, g3463, g7268, g7362, I11740, g10188, I12174, I12796;
wire g5659, g7419, I15503, I17441, g6980, I17206, g4113, g6069, g11503, g7052, g8110;
wire g2556, g4313, I16196, I7817, g8310, g10460, g2222, I11953, I13373, I6818, g4202;
wire I6867, I9880, g10093, I10484, g9845, g3720, g10267, g10294, I11800, g4908, g5111;
wire g11450, I13800, g5275, I11417, I17758, g3318, g11315, g4094, I17435, g10065, I5092;
wire g8002, g5615, g4567, I8259, g11202, g7728, g6287, I14312, I9612, g10875, I9243;
wire g11055, g3393, g9807, g11111, g4776, I9935, g4593, I11964, I7441, I15986, g3971;
wire g7070, g2237, g6399, g5284, I11423, g7470, I15741, g7897, g7025, I6370, g7425;
wire I11587, g2844, I12553, I12862, I8215, I10813, g11384, I14799, I6821, g2194, g10160;
wire g6797, g11067, g9342, I12326, g8928, g3121, I16280, g4160, g3321, g2089, g4933;
wire I14973, g2731, I16688, I11543, g5420, I15801, I12948, g10455, g8064, g4521, I14805;
wire g6291, g2557, g4050, I13117, I12904, I4873, g8785, g4450, g5794, g9097, g2071;
wire g7678, g6144, I11569, g3253, I7743, g6344, g3938, g7331, I15196, g9354, g10201;
wire g7406, g10277, g2242, I9213, g3909, I6106, g7635, I4869, I13568, I13747, I15526;
wire g8563, g10075, g4724, g6259, g4179, g7766, I5722, g7682, I13242, I17500, g6694;
wire g4379, g3519, g7801, g7305, I7411, g8295, g2955, I8136, g5628, I6061, I12183;
wire g6852, I11814, g5515, I6461, g5630, I12397, I4917, g2254, g2814, g11402, g4289;
wire g7748, g4777, I11807, g11457, I9090, g4835, I14400, g2350, g7755, g9267, g9312;
wire I13639, g2038, I8943, I16763, I12933, g7226, g8089, g10352, g2438, I11293, I13230;
wire g2773, g4271, I6904, I12508, I11638, I12634, g10155, I17613, g10822, I4786, I6046;
wire I9056, g6951, g10266, I8228, I14005, g10170, I8465, I16660, g7045, I10538, I8934;
wire I5424, I5795, g7445, g6114, I5737, I6403, I5809, g6314, I7713, g9761, I11841;
wire I11992, I11391, I9851, g2212, I13391, g6870, g4674, g8948, g3141, I6391, I5672;
wire I15688, g5040, I5077, g1983, g6825, g3710, g7369, g7602, g10167, g10194, g10589;
wire I16550, g4541, g7007, I17371, I17234, g7920, I11578, I12574, g10524, g2229, I15157;
wire I16307, g4332, I12205, g7767, I6159, g11157, g4680, g6136, g8150, g4209, g4353;
wire g5666, g6336, g8350, I13586, g10119, I8337, g8438, g6594, g11066, g4802, I13442;
wire g8009, I5304, g10118, I6016, I6757, g7793, I9279, g5648, g6806, g5875, g6943;
wire I16269, I9720, I12592, g10616, g4558, g5655, I13615, g7415, g7227, I9872, g10313;
wire I5926, I13720, I9652, I5754, I10991, I15763, I11275, g10276, g11511, g4901, I7760;
wire I16670, I11746, I13430, g10305, g10254, g4511, g10900, g9576, g2837, g10466, g5884;
wire I5044, g6433, g5839, g8229, I6654, g8993, g2620, I12846, g2462, g9349, I8815;
wire g10101, g10177, I16667, I13806, I7220, I5862, I9598, I7779, I17724, g6845, g7502;
wire I8154, I10584, I17359, g3545, I15314, g11550, I15287, g6195, I7423, g6137, g5667;
wire g6395, g3380, g5143, g6337, I16487, g6913, g10064, g11287, I15085, g2249, I9625;
wire g4580, I10759, g11307, g11076, I9232, g7188, g7689, I17121, g11596, g7388, I10114;
wire I9253, I9938, g10874, g11054, g6807, I9813, I6417, g5693, g11243, I17344, g3507;
wire g4262, g2298, g2085, I7665, g10630, g11431, g6859, g7028, I6982, g6266, I15269;
wire g10166, g7030, I12583, I9519, g8062, g7430, I15341, I5414, I16286, I7999, g2854;
wire I17173, I5946, I10849, g11341, I7633, g4889, g2941, g6248, g11655, g9258, g3905;
wire g10892, g9818, g9352, I7303, I8293, I10398, I13475, g11180, g7826, g3628, g6255;
wire g4175, g6081, g6815, I10141, g4375, I10804, I5513, g3630, g8788, I11222, I12282;
wire I15335, I16601, g5113, g6692, I16187, g6097, I7732, g7910, I12357, g2219, g9893;
wire g2640, g6154, g4285, g6354, g2031, g10907, g5202, g6960, I15694, I5378, g2431;
wire I15965, g2252, g2812, I7240, g7609, I10135, g7308, g8192, g2958, g8085, g10074;
wire g5094, I13347, g2176, g9026, g8485, g4184, g5494, g3750, g2005, g7883, I7043;
wire g4384, I9141, I9860, g5567, g4339, I9341, g10238, I16169, I9525, I14361, g2829;
wire g11619, g2765, g9821, g11502, g7758, I5916, I13236, g7066, g7589, g4424, g3040;
wire g4737, I11351, I13952, g5593, g6112, I13351, g6218, g6267, g3440, g6312, g11618;
wire g9984, I11821, g10176, g10185, g10675, I16479, g10092, I10048, I16363, I16217, g3323;
wire I15278, g7571, g7365, g2733, g4077, g6001, g7048, g10154, g2270, I5798, I17240;
wire g7711, g4523, I10221, I11790, g8520, g6293, g11469, g8219, g2225, g8640, g10935;
wire g2610, g2073, g2796, g11468, g11039, I6851, g4205, I7697, I10613, I11873, g10883;
wire I17755, g7333, g9106, I7210, g7774, g5521, g3528, g8958, I16580, I17770, g11038;
wire g5050, g2124, g3351, g5641, I17563, g2980, g6727, g8376, I5632, I5095, I6260;
wire g2069, I9111, g7196, g4551, I15601, I9311, I15187, g7803, I12248, I13209, g4499;
wire I8848, g2540, g7538, I13834, I5579, g7780, g5724, g9027, g2206, I12779, g10729;
wire g6703, I9174, I5719, g10577, I17767, g7509, g9427, I10033, I7820, I10234, g4754;
wire I16531, g10439, I11021, I12081, g5878, g6932, g7662, g4273, I16178, I12786, I17633;
wire g5658, g5777, I10795, I13726, g7467, g1990, I6118, g8225, I17191, I17719, I11614;
wire g8610, I6367, I9180, I12647, I16676, I16685, I11436, I9380, g10349, g9345, I16953;
wire I13436, I9591, I16373, g4444, g8473, g2199, g11410, g2399, g9763, g7093, I12999;
wire g3372, I10514, I12380, g10906, I15479, I13320, g10083, I9020, g8124, g10284, g7256;
wire g8980, g7816, g8324, g11479, I6193, I11593, g3143, g11363, g3343, I11122, g2797;
wire I13122, I6549, g4543, I10421, I11464, g3566, I6971, g6716, I14421, g2245, g6149;
wire g3988, I6686, g6349, g7847, g3693, I11034, I10012, g3334, I5725, g7685, g7197;
wire I11641, I11797, g5997, I15580, I13797, I6598, g7021, g4729, g4961, g7421, g10139;
wire g2344, I8211, I9905, g6398, I10541, I6121, g1963, I17324, g7263, I14473, g2207;
wire g10138, I17701, I10789, I12448, I13409, I17534, g3792, g5353, g8849, g2259, g6241;
wire g2819, I11408, I12505, I11635, I10724, g11084, g4885, g4414, I10325, g11110, g3621;
wire I6938, I7668, g2852, I7840, I16543, g10852, g8781, I8614, I10920, I10535, I12026;
wire I10434, g11179, g2701, g3113, g7562, I14358, I7390, I10828, I10946, g8797, g6644;
wire g4513, g7631, I5171, g7723, g6119, I9973, g7817, g5901, I4920, g8291, g11373;
wire g3094, g6258, g4178, g4436, g6818, g4679, g11654, g4378, g7605, g5511, I11575;
wire g3518, I10682, g10576, I9040, g8144, g8344, g6717, I9440, g11417, I13711, I16814;
wire I12433, g4335, I9123, I11109, g7751, g4182, I9323, I13109, g4288, I11537, g4382;
wire I16772, g3776, g6893, g5574, g5864, g10200, g8694, g2825, g2650, g10608, g10115;
wire g6386, g7585, I17447, I5684, I8061, g4805, I7163, I5963, I7810, g7041, I7363;
wire I16638, g2008, I13606, I12971, I11303, g6274, I7432, g6426, g11423, g2336, I16416;
wire I12369, I9875, I7453, g6170, I14506, g7673, I9655, g6125, I5707, g8886, g3521;
wire g8951, I16510, g5262, g3050, I11091, g10973, g5736, g6984, g6280, g6939, g7669;
wire I17246, g11543, g3996, g10184, I12412, I8403, g10674, g8314, g5623, g7772, I7157;
wire g7058, I12133, I5957, I7357, g2122, g2228, g7531, g4095, g9554, g8870, g2322;
wire I10927, g7458, g5889, I12229, I6962, g4495, I9839, g2230, g4437, g4102, I17591;
wire g4208, g7890, g8650, I13840, I16586, g3379, I15568, g10934, g6106, g5175, g6306;
wire g7505, g3878, g11242, I5098, g8008, I10240, g7011, g4719, g10692, g5651, I6587;
wire I10648, I15814, g8336, I14903, I5833, g6387, g5285, g6461, I15807, I15974, I8858;
wire g2550, g7074, I16720, g3271, g10400, g2845, I9282, I15639, I10563, I5584, g10214;
wire g9490, g9823, g2195, g4265, I15293, I9988, g6427, I12627, g2395, g2891, g5184;
wire g2337, I11483, g2913, g10329, g10207, g4442, I6985, g6904, g6200, g11638, g10539;
wire g4786, g6046, g8065, g3799, I8315, I8811, g6446, g8122, g3981, g8465, g9529;
wire g4164, g10538, g4233, g5424, g9348, I11326, I13949, g6403, I13326, I9804, g6145;
wire g2859, g3997, I15510, g9355, I9792, I6832, g4454, g8033, g11510, g6191, g7569;
wire g5672, g4296, I11904, I10633, I10898, g5231, I17318, g3332, I11252, g10241, g9260;
wire g6695, I10719, I13621, g5643, g3353, I7735, I6507, I14191, g8096, g2248, g11578;
wire g2342, I7782, g6107, I17540, I12857, g11014, g6307, g3744, g6536, I4883, g5205;
wire I15586, I8880, g2255, I5728, g7688, I12793, g2481, I9202, g8195, g7976, g8137;
wire g8891, g8337, g10235, g4012, I11183, I16193, g11442, g2097, I12765, g10683, g5742;
wire g2726, g4412, I11397, I13397, g2154, g6016, I12690, g4189, I5070, g2960, I10861;
wire I10573, I9567, g8807, I14573, g4888, g7126, I13933, I17377, g7326, I10045, g6115;
wire g6251, g4171, g6315, g6811, I15275, g4371, I14045, I17739, g4429, g4787, I8982;
wire g11041, g10882, g5754, I9776, I10099, I16475, g6447, I10388, I8234, g7760, I14388;
wire I8328, I17146, I16863, g3092, I14701, I10251, I14534, g4281, I9965, g5613, g6874;
wire g8142, g2112, g8342, g2218, I15983, g2267, I17698, g11035, g8255, g8081, g8481;
wire g2001, g7608, g7924, I5406, g7220, g5572, g5862, I12245, g7779, I4780, I6040;
wire g6595, g10584, I15517, I13574, g2329, g8354, I14140, g7023, I7952, g4963, g10206;
wire I5801, I7276, g9670, I16781, g4791, g7977, g2828, g6272, I16236, g3262, g2727;
wire g3736, g5534, g5729, g7361, g10114, I16175, g9813, I15193, g6417, I13051, I15362;
wire g6935, g11193, g7051, g10107, I11756, g2221, g3076, I13592, g8783, I15523, g7327;
wire I12232, I6528, I16264, g8979, I16790, I8490, g4201, I6648, g8218, I9658, g8312;
wire I7546, g6128, g6629, g5885, g10345, g7999, g7146, g5660, I5445, g6330, g7346;
wire I10162, g7633, g4049, g3375, g8001, I12261, g4449, g3722, I8456, g7103, g5903;
wire g4575, g10848, g11475, g8293, g8129, I6010, g2068, I11152, g8329, g10141, g7696;
wire g10804, g6800, g4098, g3500, I15437, I16209, I8851, I11731, g8828, g11437, g2677;
wire g10263, g7753, I9981, g8727, g5679, g7508, g3384, g10332, g6213, g8592, g7944;
wire I15347, g7072, I15253, g10135, I12445, g11347, g4896, I7906, g2349, g7043, I12499;
wire I11405, g5288, g9341, g3424, I9132, g10361, g3737, g7443, I9332, g9525, I9153;
wire I9680, I10147, I6343, I10355, g7116, g5805, g5916, g7316, g2198, I6282, g4268;
wire I7771, I16607, g2855, g4362, I11929, I14355, I12989, g11351, g3077, g5422, g7034;
wire I10825, g4419, I9744, I12056, I10370, g6166, g8624, g3523, I14370, g8953, I10858;
wire I13020, I13583, g4452, I8872, I15063, g2241, g7147, g6056, g5947, g7347, g11063;
wire I11046, I10996, I12271, g7681, g6649, I8989, g8677, g110, I10367, I10394, I9901;
wire g7697, I14367, I14394, I16641, g3742, g7914, g8576, g2524, g7210, g4728, I16292;
wire g2644, g6698, g4730, g8716, I17546, g8149, g10947, g4504, I11357, g6964, g8349;
wire g2119, g5095, g6260, g5037, I13357, I12199, g4185, I7244, g9311, g11422, I11743;
wire I13105, g5653, g4385, g7413, g5102, g2258, I14319, g2352, g2818, I7140, g6063;
wire I12529, I5940, g2867, I16635, g10463, g11208, g4470, g8198, g4897, g8747, I7478;
wire g5719, g4425, I12843, I15542, g10972, g10033, I5388, g10234, I7435, g7936, g11542;
wire g11453, g5752, I6094, I13803, g3044, g2211, I14540, g6279, g2186, g7317, g6720;
wire I8253, g6118, g3983, g11614, g7601, I5430, g5265, g11436, g3862, g5042, I15320;
wire g9832, g6652, g4678, g6057, g6843, I15530, g11073, g4331, g3543, g2170, g2614;
wire g7775, g11593, g7922, g2125, g8319, g11346, I15565, g2821, g9507, I15464, I6965;
wire I10120, g4766, I11662, I10739, g4087, g4105, g8152, g10421, I16537, g8352, g4305;
wire g6971, I13027, I12258, g3729, I6264, I16108, g6686, g10163, g8717, g11034, g7460;
wire g7597, g5296, I11249, I5638, I14645, I16283, g2083, I6360, g4748, I16492, I13482;
wire I5308, I11710, g7784, I4992, g4755, g10541, I10698, g6121, I15409, I7002, g8186;
wire g10473, g4226, I11204, g6670, I7402, g11409, I6996, g3946, I13779, I7236, I15635;
wire I16982, g8599, g7995, g2790, g11408, g7079, g11635, I11778, g3903, g5012, g9100;
wire g8274, I10427, g7479, g8426, g1994, g4445, g6253, g2061, g2187, g6938, g4173;
wire g6813, g4373, I11786, I16796, g10535, g4491, g8125, g7190, g8325, I11647, g7390;
wire I12878, g5888, I13945, I12171, g10121, g8984, g3436, g4369, g8280, I7556, g4602;
wire g7501, I17450, g3378, g5787, I9424, I9795, I17315, g10344, I9737, g2904, g2200;
wire g6552, g7356, g2046, I17707, g4920, I5827, g2446, g4459, I17202, g3335, I13233;
wire g8483, g4767, I7064, g11575, g2003, g5281, g3382, I9077, I7899, g4535, I8358;
wire I6611, I8506, g2345, g10173, I17070, g8106, g11109, g8306, g2763, g2191, g2391;
wire g6586, I12919, I6799, I11932, g3749, g8790, I9205, g11108, g2695, g9666, g8061;
wire g5684, I8275, I8311, g4415, g5639, I14127, I17384, g7810, g7363, g10134, I7295;
wire I11961, I16553, g5109, g5791, g3798, I13448, I9099, g2159, g7432, I14490, g6141;
wire g8622, g6570, g6860, g7053, I11505, g9351, I5662, g9875, g8427, I5067, g9530;
wire g6710, g5808, I5418, g2858, I12598, I7194, I14376, I14385, g4203, I8985, I13717;
wire g11381, g4721, g2016, I13212, g2757, g8446, g7568, g5759, I9754, I10888, g8514;
wire I6802, g3632, g3095, g3037, g8003, I14888, I16252, g3437, I12817, I9273, I10671;
wire I17695, g3102, I4924, g3208, I12322, g7912, g8145, g8345, g2251, g2642, I12159;
wire g7357, g2047, I12532, I12901, g8191, g10927, g9884, g6158, g3719, I12783, g11390;
wire I13723, g5865, g8695, I5847, I6901, I11149, g2874, g7929, g3752, I16673, I11433;
wire I16847, I11387, g5604, I13433, g5098, g2654, I11620, g4188, g5498, I9712, g6587;
wire g4388, g10491, g10903, I11097, I5421, g8359, g6111, g6275, g6311, g4216, g10604;
wire g9343, g8858, g4671, g2880, g4428, g2537, I10546, g5896, g4430, I14546, I7438;
wire g3164, g3364, I7009, I10024, I8204, I12631, g8115, g4564, g8251, g8315, g2612;
wire I15326, g2017, g6284, g2243, g8447, I6580, g3770, g6239, g10794, I15536, g10395;
wire g5419, g9804, g10262, g7683, g11040, g10899, g6591, I11412, g5052, I13412, I5101;
wire g8874, g3532, g7778, g2234, g6853, I10126, I10659, I16574, g2629, g4638, g2328;
wire I12289, I6968, g6420, g11621, g2130, g10191, g2542, I8973, g2330, g7735, I16311;
wire g4308, I11228, I17231, g7782, g6559, I12571, g3012, I11011, I5751, g8595, g6931;
wire g5728, g5486, I10296, I11716, g5730, g5504, g7949, g4217, g11183, I8123, g3990;
wire g2554, g4758, g4066, g8272, I16592, g4589, g5185, g11397, g5881, g7627, g9094;
wire I5041, I9135, g4466, g1992, g6905, g8978, I5441, g3371, g11062, I10060, g2213;
wire g11509, g7998, g10247, g4165, g4365, I13627, g5425, g10389, g10926, I10855, I13959;
wire I13379, g11508, g4711, g6100, I11112, g8982, g11634, g10612, g6300, g7603, g4055;
wire g7039, I9749, g10388, I8351, g8234, g2902, g7439, g8128, g8328, g7850, g10534;
wire g10098, I17456, g4333, I7837, g8330, g10251, g10272, g2090, g4774, I7462, I9798;
wire I13096, g2166, g6750, g9264, I6424, g7702, g4196, g5678, I10503, I16413, g10462;
wire g4396, g3138, g8800, I14503, I8410, g2056, I16691, g9360, g3109, g3791, g2456;
wire g7919, g10032, g2529, g2649, g10140, g4780, I8839, g6040, g2348, I6077, g11574;
wire g11452, g11047, g5682, g5766, g5105, g4509, g6440, g1976, g11205, I6477, I9632;
wire g7952, I15311, g9450, g5305, g5801, I5734, I6523, g2155, I4820, I17243, g2355;
wire g2851, I7249, I12559, I14315, I6643, g8213, I10819, g11311, I10910, I12424, I9102;
wire I9208, g3707, I9302, I14910, g7616, g7561, g4067, g3759, I8278, I14257, g5748;
wire I10979, g2964, g4418, I9869, g4467, I15072, I14979, g4290, I10111, I14055, g10871;
wire g11051, I5992, g7004, I16583, g11072, I17773, I15592, I15756, g7527, I17268, I6742;
wire I12544, g4093, I8282, g6151, g7764, g4256, g6648, g9777, g7546, I5080, I15350;
wire I10384, g10162, g3715, I9265, I16787, g11350, I5713, I15820, g5091, g8056, I13317;
wire I12610, g4181, I6754, g8529, I14094, g4381, g7925, I9786, g2118, g8348, I12255;
wire I6273, g2872, I16105, g10629, I10150, g5169, g4197, I10801, g8155, g11396, I13002;
wire g8355, g10220, g5007, I13057, g2652, g2057, g10628, I12678, I13128, g2843, g10911;
wire g7320, g2989, g3539, g4263, I13245, I11626, I16769, g5718, I12460, I12939, g5767;
wire I15691, I9296, I10018, I11299, I13323, I7176, I5976, g2549, I6572, I10526, g8063;
wire g2834, g2971, g6172, g6278, g7617, I7405, g7906, g7789, g11405, g5261, g10591;
wire I6543, g3362, g3419, I7829, g6667, g7516, g4562, g6343, g10754, g9353, g3052;
wire g10355, g5415, g6282, g7771, g6566, I11737, g8279, g2121, g4631, I12875, g10825;
wire I10917, I15583, g9802, g1999, I11232, g4257, g6134, g5664, g8318, g8872, I9706;
wire g2232, g10172, g11046, g3086, g5203, g2253, g3728, g2813, I9029, g8989, I14077;
wire I9171, g6555, I10706, I9371, g6804, I15787, I6414, g3730, g2909, I9956, I10689;
wire g3385, I5383, I15302, g11357, g7991, I6513, g2606, g10319, g4441, g6113, g6313;
wire g7078, g7340, I10102, I16778, I13831, g10318, I8050, I13445, I5588, g8121, g10227;
wire g7907, I6436, I6679, g8321, g4673, g6202, g8670, g5689, I8996, I9684, g7035;
wire I15768, I9138, I9639, g7959, I10066, I9338, I10231, g8625, g7082, g2586, g5216;
wire g10540, I17410, g6094, I11498, I12595, I16647, g10058, I16356, g4669, I8724, g6567;
wire g5671, g4368, I11989, I17666, I10885, I8379, g3331, g10203, I14876, I11611, g7656;
wire g4772, g3406, I11722, I7399, g10044, g3635, I6022, g4458, g2570, g2860, g2341;
wire g9262, g3682, g6593, I9759, g8519, g3105, g7915, g3305, g10281, g98, g2645;
wire I8835, g5826, I12418, I12822, g10902, g10377, g8606, g7214, I6947, g10120, g4011;
wire g9076, g5741, g3748, g4411, g4734, I11342, g9889, g7110, g6264, g7310, I6560;
wire I7291, I8611, I10456, I15482, g5638, g3226, g6933, g7663, I11650, g10699, g2607;
wire I12853, I16897, I5240, g2962, g6521, I17084, g4474, g10290, g2158, g6050, g6641;
wire I11198, I9498, I12589, g10698, g2506, g6450, I6037, I17321, g5883, I10314, g7402;
wire I6495, I9833, I17179, I11528, I6102, I16717, I17531, I7694, I11330, I6302, g3373;
wire I15778, g7762, g3491, g4080, I5116, g11081, I7852, I7923, g5758, g8141, g8570;
wire g5066, g5589, g6724, g8341, I10054, g2275, I9539, I9896, g4713, I10243, I11132;
wire I11869, g7877, I7701, g3369, I5565, g3007, g9339, I15356, g7657, g6878, I15826;
wire I6917, I15380, I4894, g2174, g3459, g6289, g9024, g2374, I12616, I9162, g7556;
wire I9268, I16723, g3767, g10547, g9424, g10895, I7886, I9362, g6835, g2985, g9809;
wire g5827, g6882, g7928, I10156, I10655, I15672, g3582, I16387, I17334, g6271, I11225;
wire g10226, I9452, g11182, g11651, g7064, I5210, g2239, I10180, g9672, I13708, g5774;
wire g7899, g3793, g7464, I12053, g8358, I12809, g7785, I16811, g10551, I6233, g2832;
wire I12466, g3415, g3227, I7825, g6799, g2853, I11043, I6454, I13043, I17216, g2420;
wire g6674, I9486, g11513, I12177, g10127, g3664, g8275, g2507, g8311, g3246, I15448;
wire g5509, g4326, I14694, I7408, g7237, g10490, I9185, I7336, g3721, g11505, I11602;
wire I11810, g11404, g6132, g5662, I6553, I4850, g7844, I17543, I11068, I13068, g6680;
wire g6209, g8985, I11879, g5994, g10889, I16850, I11970, g7394, I10557, g10354, g2905;
wire g7089, g7731, g10888, g6802, g8239, g4183, g9273, g4608, g5816, I5922, I7465;
wire g7966, g2100, I10278, g3940, g6558, I12009, I6888, I8262, I11967, g8020, I10286;
wire g8420, I5060, g10931, g3388, I10039, I14306, I11459, g11433, g9572, g5685, g5197;
wire g5700, g8794, g5397, g2750, I8889, g11620, g10190, I8476, g4361, I9766, I15811;
wire g3428, I7096, I12454, I9087, I9105, I9305, I9801, g3430, g7814, I12712, g11646;
wire g4051, I10601, I13010, g11343, I13918, I16379, g4127, g4451, I15971, g4327, I17265;
wire g7350, g2040, g6574, I12907, I5995, I11079, g10546, g7038, I11444, I17416, g10211;
wire g9534, g9961, g6714, g7438, g7773, I11599, g7009, g11369, g2123, I6639, g4346;
wire g8515, g10088, I8285, I10937, I12239, I5840, I15368, I17510, I16742, g8100, I16944;
wire g3910, I13086, g7769, I15412, g3638, I8139, g7212, g5723, I14884, g11412, I11817;
wire I10168, g5101, g5817, I11322, g7918, g5301, g7967, g6262, I15229, g2351, I11159;
wire g10700, g2648, I9491, g10126, I8024, I11901, I16802, g2530, g6736, I13125, g8750;
wire I10666, g4508, g10250, g2655, g4944, g4240, I11783, I16793, I7342, I9602, g4472;
wire I10015, I5704, g7993, I7255, g6076, I4906, I11656, I6049, g5751, g3758, g3066;
wire I8231, g4443, g10296, g8440, I11680, g8969, I17116, g2410, g9679, I7726, g6175;
wire g4116, I7154, g8323, g6871, g2884, I7354, g2839, g3365, g3861, I6498, I17746;
wire g3055, I5053, I15959, g6285, g11627, g7921, g10197, g5673, g4347, I8551, I10084;
wire g2172, g3333, I9415, g11112, I17237, g4681, g10870, g11050, I8499, I12577, g8151;
wire g10527, g3774, g8351, I17340, g4533, I13017, I13364, I15386, g6184, g2235, g2343;
wire I12439, g5669, I10531, I17684, g6339, I14179, g4210, I14531, I7112, I17142, g11096;
wire g7620, g4596, g3538, I6019, g4013, g6424, I16626, I10186, g6737, g10867, g2334;
wire g10894, g6809, I10685, g5743, g4413, g5890, I11289, I6052, g2548, I14373, I11309;
wire I5929, I13023, g8884, I16298, I13224, g7788, g6077, g11429, g5011, I16775, g3067;
wire I13571, g10315, g5856, g5734, g10819, g11428, g10910, g3290, I17362, g10202, I10334;
wire g10257, g4317, g8278, I4876, g3093, g1998, g5474, g10111, g7192, g5992, g7085;
wire g3256, I7746, g6634, I9188, I10762, g8667, g3816, g8143, I13816, I15548, I6504;
wire I9388, g8235, g8343, g6742, g11548, g6104, I14964, g10590, I9216, I6385, g6304;
wire I16856, g8566, g6499, I16261, g2202, g11504, g8988, g4775, I11752, g8134, g7941;
wire I15317, I6025, g2908, g8334, g9265, g6926, g2094, I12415, g11317, g10094, g3397;
wire g8548, g2518, g4060, g4460, I9564, I7468, g6273, I8885, g8804, I14543, I8414;
wire g10150, g10801, I9826, I10117, g7708, I13669, g10735, g10877, g11057, g7520, g8792;
wire I17347, I7677, I11668, g6044, g2593, g7031, g4739, I8903, g6444, g11245, g7431;
wire I15323, g6269, I15299, g7812, g11626, g9770, g10196, I11489, g10695, g5688, g11323;
wire I13489, g2965, I6406, I5475, I7716, g6572, g6862, g7376, I5949, g10526, g8313;
wire I12484, I14242, I9108, I15775, I13424, g4479, g9532, I9308, g6712, I8036, g4294;
wire I10123, g6543, g4840, I8436, g9553, I5292, I9883, I14123, g3723, g7765, g7286;
wire g4190, I5998, g4390, I10807, g10457, g3817, g7911, I5646, I10974, g8094, g2050;
wire g2641, I8831, I15232, I10639, I17516, g2450, I16432, g4501, g8518, g6729, g6961;
wire g8567, I10293, g4156, I11713, g7733, I5850, g7270, g9990, g6927, g3751, I9165;
wire I16461, I9571, I9365, g7610, g2179, g4942, g9029, g6014, g7073, I12799, g7796;
wire I12813, g6885, g9429, g22, g7473, I10391, I17209, g6660, I11255, g10256, I6173;
wire g11512, I13255, I14391, I16650, I6373, I6091, g5183, g7124, g7980, g7324, g10280;
wire g6903, g2777, I5919, I11188, g7069, I12805, I13188, g5779, I13678, I14579, g4954;
wire g4250, g4163, I5952, g2882, g7540, g8160, g4363, I11686, I16528, I7577, I5276;
wire g8360, I16843, I6007, g5423, I13460, I17453, I11383, g2271, g7377, g7206, g10157;
wire g11445, g6036, I5561, I13030, g2611, g4453, g8450, g6178, I6767, g11499, I8495;
wire g3368, g9745, I11065, I6535, g1987, g9338, g7287, g2799, g11498, I5986, g6135;
wire g5665, g9109, g6335, I15989, g9309, g3531, I8869, g5127, g3458, g6182, g6288;
wire I17274, g6382, I9662, g8179, g7849, g10876, g10885, g11056, g3743, g8379, g4912;
wire I14116, g2997, g11611, I12400, g2541, g11080, I7426, I9290, g5146, g10854, g6805;
wire g5633, g3505, g7781, I5970, g6749, I16708, g2238, g11432, I13837, g3411, I9093;
wire g7900, I16258, I4948, g2209, g7797, I9256, I8265, I9816, g5696, I15461, g6947;
wire I7984, I5224, I7280, I10237, g6798, I8442, I12538, g8271, g2802, g11342, I10340;
wire g1991, I5120, g3474, g9449, g6560, I14340, g5753, I8164, I15736, g10456, g5508;
wire g11199, I14684, g11650, g7144, I11617, g7344, g5072, I7636, I13915, g5472, g8981;
wire I9421, g8674, I5789, g5043, I11201, g10314, g7259, g5443, g6208, I7790, I16879;
wire g6302, g10307, I15365, I7061, g6579, g5116, g6869, g7852, g7923, I17164, I7387;
wire g10596, I11467, I11494, I13595, g8132, g6719, I12235, g8332, g10243, I11623, I12683;
wire I6388, g8680, g10431, I11037, g8353, I14130, I10362, g2864, I10165, I13782, g6917;
wire g4894, I6028, g10269, g8802, I6671, I6428, g7886, g4735, I17327, g6265, g3976;
wire I6247, g4782, I11155, g10156, I15708, I17537, I13418, I13822, g5697, I10006, g6442;
wire g9452, g7314, g5210, I17108, g11471, I7345, I16458, I8429, I9605, g4475, g5596;
wire g6164, I7763, I7191, g10734, I10437, g10335, g7650, g3326, I15244, g4292, g10930;
wire g11043, g6454, g11244, g4526, I5478, g6296, I11194, g3760, g7008, I13194, I13589;
wire g2623, I17381, I7536, I9585, g2076, g10131, g2889, I11524, I16598, g11069, g4084;
wire I11836, I5435, g4603, g5936, g7336, g8600, I15068, g7768, g4439, g11657, g5117;
wire g6553, g8714, g11068, I7858, I11477, g7594, g10487, g7972, g2175, I11119, g9025;
wire g2871, g10619, I12759, I7757, I16817, I9673, I14236, g7806, I10952, g3220, I8109;
wire g2651, I6217, g4583, g6412, I17390, g10279, g7065, I7315, g6389, I7642, I9168;
wire g6706, I9669, g7887, g7122, I15792, I9368, g7322, g4919, I10063, g6990, I7447;
wire g10278, g3977, I6861, g6888, I16656, I9531, g6171, g2184, I16295, I9458, g3161;
wire I11704, I12849, I6055, I17522, g2339, g7033, g10039, I10873, g6956, g5597, I14873;
wire I7654, I13809, I6133, g3051, g2838, g8076, g2024, I15458, I13466, I9505, g6281;
wire g8476, g3327, g2424, I8449, I12652, g9766, g2809, g5784, g4004, I9734, I13036;
wire I5002, I8865, g7550, g6297, I11560, g10187, I6196, I5824, g7845, I10834, g8871;
wire g8375, I15545, g3633, I15079, I8098, g2077, g2231, g7195, g11545, g11079, g11444;
wire g5937, g7395, I13642, g7337, g3103, I9074, g7913, I6538, g2523, I7272, g2643;
wire I9992, g10143, g5668, g11078, g6338, I15598, I10021, g5840, g4970, g8500, I7612;
wire g11598, I7017, g6109, I12406, g6309, g11086, g7807, I7417, g3732, I17252, g10169;
wire I7935, I9080, g8184, g10884, g6808, I15817, I9863, g8139, I16289, g8339, g2742;
wire g3944, g10168, I10607, g6707, I13630, g2304, g11322, g9091, g4320, I15977, g11159;
wire I10274, I11166, I11665, I16571, I13166, I7330, I8268, g8424, I5064, g8795, g10217;
wire g7142, I6256, g4277, g6201, g7342, I11008, g6957, I15353, g2754, g4906, g7815;
wire g11656, g4789, I7800, g10486, g11353, g8077, I15823, g6449, I13485, g2273, g8477;
wire g6575, g7692, I12613, g8523, I6381, g9767, g7097, I9688, g7726, I9857, I13454;
wire g2613, g7497, g9535, g6715, g2044, g7354, g10580, I10153, g2444, I5237, g5032;
wire g2269, g10223, I7213, g9261, I6421, g4299, I14409, I12463, g3697, g8099, I8385;
wire I14136, g8304, g3914, I9126, I13239, g10110, g11631, I9326, g2543, g6584, g11017;
wire g6539, g6896, g5568, g10321, I5089, I5731, I11238, I17213, g7783, g10179, g10531;
wire g7979, g3413, g5912, g7312, I7166, I5966, g10178, I7366, g4738, I13941, I13382;
wire g6268, I11519, I11176, g10186, g7001, g8273, g10676, g6419, I10891, I13185, g11289;
wire I7456, g1993, g3820, g7676, g4140, g6052, g11309, g4078, I12514, g8613, I16525;
wire I7348, g6452, I9383, I9608, I15308, g7329, g4478, g7761, g2014, g4907, g8444;
wire g2885, I9779, g2946, g4435, I9023, g8983, g4082, I12421, I8406, I5254, I14109;
wire g8572, g7727, I7964, g2903, I7260, I14537, I10108, g6086, g8712, g11495, I12012;
wire I9588, g7746, I8487, I5438, g3775, g7221, I17350, I14303, g6385, g6881, I12541;
wire g7703, I9665, I15752, g4915, g2178, g2436, I15374, g9028, g8729, g8961, I4900;
wire I11501, I16610, g9671, I17152, g3060, I13729, I13577, I10381, g4214, I16255, I14982;
wire g6425, I11728, g11643, g2135, I16679, g2335, g5683, I13439, I9346, I7118, g4310;
wire g2382, I7318, I12829, I16124, g10909, I12535, g5778, I10174, I15669, g10543, g3784;
wire I17413, g5894, g9826, g10117, g8660, g8946, g10908, g2916, I7843, g2022, g5735;
wire I15392, g7677, g2749, g3995, g3937, I10840, g9741, g4002, I7393, I16938, I6531;
wire I11348, I12344, I13083, g3479, g11195, g11489, g6131, g5661, g10747, I15559, g5075;
wire g8513, I15488, I15424, g6406, g10242, I8007, g5475, g4762, g2798, g5949, g7349;
wire I10192, g11424, I9240, g6635, I11566, g11016, g9108, g3390, g9308, g8036, g2560;
wire g5627, g8436, g8178, g6801, g6305, I6856, g4590, g7848, g5292, I10663, g8378;
wire g9883, I9043, g3501, I14522, I8535, I9443, g7747, g5998, g5646, g10974, g8335;
wire g2873, g6748, g2632, I6074, g2095, I11653, g2037, g8182, I4886, g4222, g5603;
wire I6474, I7625, g5039, I4951, g10293, g2653, g2208, g2302, I12029, g5850, g6226;
wire I10553, g3704, g8805, g10265, g2579, I5837, I7938, I9147, I13636, g8422, I10949;
wire I17302, g4899, I11333, I13415, g4464, g2719, g9448, I7909, I6080, I14326, g4785;
wire g11042, g10391, I6480, g5702, g6445, g2752, I14040, I14948, g9827, g6091, I10702;
wire g3810, g3363, I10904, g8798, g7119, g7319, g3432, I6569, g10579, g4563, g9774;
wire I7606, g8560, I14252, g6169, I15383, I16277, g6283, g7352, g2042, g4295, g10578;
wire I9013, g4237, g6407, I14564, g6920, g6578, g6868, g5616, I16595, g8873, g8632;
wire g8095, g2164, g6718, g2364, g2233, g9780, g4194, I16623, g8437, I10183, I7586;
wire g11065, g4394, I5192, I6976, g2054, g6582, I13609, I14397, g7386, g4731, I11312;
wire g5647, g2454, g8579, g8869, g7975, I13200, g6261, I11608, g2296, I11115, I12604;
wire g10116, I9117, g6793, g8719, g4557, I9317, g2725, g1974, I14509, g5546, g7026;
wire I5854, I8388, g4966, I12770, I14933, g7426, g9994, g9290, I11921, I17662, I12981;
wire g8752, g6227, g10041, g5503, I7710, g7614, g10275, g4242, g10493, g7325, I17249;
wire g4948, I7691, g9816, I17482, g10465, g1980, I8247, g7984, g2012, g11160, g8442;
wire I17710, g6203, I17552, I16853, I9581, g10035, g5120, I5031, g5320, g4254, I16589;
wire I11674, g10806, g7544, g8164, I13674, I15470, I5812, g8233, g11617, I6183, g11470;
wire I7659, g10142, g2888, I6924, g7636, I6220, I4891, g2171, g4438, I14452, g4773;
wire g7306, I13732, g8296, g2956, I15075, g8725, g7790, g9263, g3683, g11075, I5765;
wire I15595, I15467, I15494, I17356, g8532, I8308, g7187, I7311, g4769, g5987, I11692;
wire g7387, g11467, I9995, I12832, I4859, I10051, I10072, g4212, I9479, g6689, g10130;
wire g7756, g2297, g11623, g6388, g10193, I16616, g11037, I10592, g5299, I10756, I15782;
wire g7622, g3735, g7027, g7427, I17182, g10165, I13400, g10523, I17672, g3782, I13013;
wire g5892, I11214, g7904, g11419, g2745, g2639, g6030, g2338, g11352, I15418, I5073;
wire I13329, I11207, g7446, g3475, I6999, g11155, I7284, I15266, g8990, I9156, I12099;
wire I11005, I12388, I17331, I13005, g8888, g7403, g3627, g4822, g8029, g6564, I16808;
wire g8171, g7345, I17513, I8711, g2808, g3292, I10846, g8787, I12251, g7763, I16101;
wire g8956, g2707, I8827, g10437, I8133, g2759, I8333, I7420, g7637, I15589, g5078;
wire g3039, g2201, g3439, g7107, I7559, g7307, I12032, g8297, g10347, g5035, I6944;
wire I8396, g10253, I6240, I7931, g7359, g6108, g6308, I9810, g5082, g2449, I9032;
wire I11100, g5482, I14405, g10600, g11401, g10781, I4783, I6043, I9053, g8684, g3583;
wire g4895, g5876, g8138, I6443, I11235, g8338, g10236, g7757, g2604, g4062, g2098;
wire I11683, g5656, g7416, g4620, g10351, g4462, I15864, I5399, g6589, I12871, g10175;
wire g10821, I7630, I15749, g2833, I6034, g7522, I8418, g7811, g7315, g11616, I17149;
wire I6565, g7047, I7300, g11313, I12360, I8290, g10063, I17387, g8707, g6165, g10264;
wire g6571, g6365, g6861, g5214, g10137, g6048, I11515, g9772, I11882, I5510, g2539;
wire g2896, I6347, I15704, I5245, g6448, g9531, I15305, g6711, g6055, I12162, I17104;
wire g10873, g11053, I8256, g9890, I10282, g3404, g6133, g11466, g5663, I10302, I6914;
wire g9505, g2162, I7973, I15036, g2268, g8449, g4192, I10105, g4298, g3764, I12451;
wire g6846, g11036, I12472, g8575, g3546, I14105, g4485, I6013, g5402, g6196, g7880;
wire g6396, g7595, g6803, g7537, g5236, I17368, g8604, g10208, I16239, g11642, g8498;
wire I11584, g1972, I8421, g9474, g7272, I13206, g10542, g6509, g11064, I15733, g7612;
wire g7243, g2086, I11759, I11725, I12776, g5657, g10913, I16941, g2728, I13114, g6418;
wire I11082, g7982, g4520, g5222, I17228, g11630, g2185, g4219, g6290, I7151, g2881;
wire I7351, I16518, I6601, I7648, I12825, g10320, g10905, g7629, I15665, g7328, g2070;
wire g10530, g3906, I17716, g7330, g10593, I4866, g8362, I13744, g2025, I11345, g10346;
wire I8631, g5899, g8419, g4958, g6256, g4176, g6816, g10122, g4376, g4005, g10464;
wire I10027, I15476, I15485, g7800, g10034, g6181, I11804, I14249, g11454, g6847, g10292;
wire I9475, I10248, g6685, g6197, g6700, I17112, I10710, g6397, I10003, g7213, I10204;
wire I14552, I5336, g2131, g8486, I6784, g2006, g2331, I16577, g4733, g2406, g5844;
wire I13332, g6263, g4270, I11135, I7372, g10136, g2635, I16439, I17742, I12318, g11074;
wire g6950, g11239, I10081, I17096, g4225, I15238, g2087, g11594, g3945, I7143, I5943;
wire g2801, g5089, I13406, I9084, g3738, I13962, I14786, g7512, g8025, g9760, I6294;
wire I17681, g8425, g3709, g4124, g4324, g2748, g6562, g7366, g10164, I11833, I11049;
wire I15675, g4469, g5705, g5471, g2755, g11185, g7056, I17730, g3907, g10891, g2226;
wire I6501, I10090, g6723, I13048, g6257, I14090, g11518, g4177, I6156, g6101, g7148;
wire g6817, g7649, g5948, g6301, g7348, I6356, g4377, g4206, I10651, g3517, g10575;
wire I14182, I14672, g7355, g2045, g7851, I17549, g3876, g8131, g10327, g8331, g2173;
wire I12120, g2373, g4287, I9276, g10537, I10331, g7964, g8635, g6751, I12562, I8011;
wire I11947, g8105, g2169, I5395, I14449, g10283, g2369, I5913, I11106, g8487, g2602;
wire I11605, g4199, g6585, g2007, g5773, g10492, g4399, g7463, g2407, I6163, g2920;
wire I14961, g2578, g2868, g3214, g4781, g6041, I6363, I7202, I15729, I13812, I9647;
wire g4898, g6441, I13463, g9451, g4900, I6432, g11501, g3110, g11577, g7279, g5836;
wire g4510, g11439, g3663, I12427, g10091, g9346, I12366, g2261, g7619, g7318, g2793;
wire g4291, g7872, g11438, g10174, g10796, I16664, g9103, I8080, g2015, g6368, g8445;
wire I7776, g7057, g2227, g4344, I5142, I7593, I5248, g7989, I9224, I15284, g3762;
wire I12403, I12547, g4207, g11083, g11348, g10390, I16484, g9732, I5815, I9120, g11284;
wire I9320, g2246, g5822, g4819, g3877, g9508, I12226, g8007, I7264, g11622, g2203;
wire g7686, g10192, I10620, I5497, I6929, I12481, I13421, I16200, g8868, I5960, I7360;
wire I14097, I9617, g6856, g6411, g6734, I9789, I10343, g8535, I7450, I10971, g7321;
wire g8582, g7670, I17261, g4215, I7996, g11653, g2502, g4886, g4951, I16799, g7232;
wire I12490, g10553, g8015, I15415, g5895, g7938, I8126, g7813, I5979, g4314, I5218;
wire g5062, I13788, g9347, I12376, g10326, g5620, g7909, g2689, I12103, I11829, g6863;
wire I16184, I16805, g10536, g8664, g10040, I10412, I12354, g2216, g9533, g6713, I14412;
wire g7519, I13828, g10904, g2028, I14133, g10252, g8721, g6569, g10621, g7606, I6894;
wire I13344, I10228, g2247, I14228, g4336, g3394, I5830, g2564, g7687, g4768, g11576;
wire I10716, I13682, g3731, I15554, g2826, I6661, g6688, I11173, g10183, g6857, g5192;
wire g5085, I5221, g9820, g4943, I12190, I7674, g11200, g10062, g3705, I16214, I17271;
wire I12520, g2638, g4065, I8161, g4887, g4228, g4322, g7570, g2108, g5941, I14379;
wire g2609, g4934, g7341, I11029, g10851, g10872, g11052, I5932, I10958, g6400, I14112;
wire I10378, g7525, I7680, I14958, g2883, g8671, I6484, I6439, I9915, g3254, g9775;
wire I17736, I15798, g3814, g5708, I10096, g2217, g2758, g5520, I14944, I17198, I15184;
wire g4096, g8564, g3038, g4496, I8303, g11184, g5252, g7607, I17528, I6702, g3773;
wire g5812, g3009, I14681, g2165, g6183, g2571, g7659, g2861, g7358, g4195, g5176;
wire g6220, I5716, g10574, I17764, I5149, g4395, g10047, g4337, g4913, I17365, I14802;
wire g10205, g2055, g3769, g10912, g10311, g2455, g9739, g2827, I6952, I14793, g3212;
wire I9402, I12339, I8240, g1975, I5198, I12296, g7311, g2774, I6616, g3967, I17161;
wire g6588, I4935, I12644, g2846, I9762, I10549, g9079, I13648, g10051, I14690, g6161;
wire I14549, g7615, g6361, g2196, g4266, I7600, g9668, g2396, g10592, I15400, g2803;
wire g5733, I17225, g11400, g6051, I11770, g5270, g7374, I11563, I8116, g6127, g6451;
wire g8758, g8066, g8589, I15329, g7985, I17258, g4142, g2509, I16407, I15539, I6546;
wire g5073, g10350, g11207, g1984, I10317, g7284, g11539, g6146, g10820, g4081, g7545;
wire g9356, g8571, I8147, g2662, g5124, g2018, g5980, g2067, g7380, g8448, g6103;
wire I10129, I9930, I11767, I11794, g8711, g7591, g6303, g2418, I11845, g5069, I13794;
wire I10057, g4726, g2994, g5469, g7853, g4354, I5258, g7020, I5818, g8133, g8333;
wire g7420, I15241, I11898, g5177, g6732, I12867, I17657, I13633, g11241, I16206, I10299;
wire g2256, I11191, I11719, g7559, I14323, g10691, g7794, I7076, I13191, I14299, I7889;
wire g8196, g6944, g8803, I6277, g6072, I15771, I9237, I17337, g2181, g8538, g2381;
wire g9432, I15235, I6789, I16114, g4783, g6043, I12910, I7375, g2847, g8780, g6443;
wire I12202, g8509, g9453, g4112, g7905, g2197, I7651, g4312, I8820, I11440, g10929;
wire I12496, g2021, I9194, g7628, I9394, g6116, g2421, g7630, g4001, I12978, I14232;
wire g10928, g8067, I9731, g5898, g8418, g6434, g4676, g5900, g6565, I5821, I6299;
wire I11926, g8290, I12986, g4129, g5797, g4329, I14697, g4761, g11515, I7384, I13612;
wire g5245, I7339, I13099, I12384, g8093, I13388, g6681, I11701, I11534, g10787, g5291;
wire g3392, I11272, g10282, g7750, g3485, g2562, g6697, g5144, g4592, g6914, I17444;
wire g5344, g6210, I12150, g4746, g8181, g10827, g6596, I6738, g4221, g8381, g2101;
wire g2817, g3941, g7040, g6413, I10831, g7440, g8197, g8700, I10445, I7523, I11140;
wire I12196, g2605, g11441, I9150, I10499, g8421, g7123, g5088, g11206, g7323, I14499;
wire I6907, I12526, g10803, I7205, I9773, I15759, I11061, I15725, g5701, g3708, g4953;
wire g2751, g3520, g8950, I16500, g3219, I6517, I6690, I9409, I15114, I5427, g4468;
wire I15082, g6117, I14989, I17158, g3252, g10881, I7104, g11435, I6876, I9769, g11082;
wire g3812, I7099, I12457, I10924, g5886, g11107, I9836, I14080, g7351, g2041, g7648;
wire g7530, I11360, g8562, I15744, I13360, I17353, g3405, g5114, I5403, g9778, g5314;
wire I11447, g11345, g9894, g8723, g4716, I11162, I16613, g11399, g3765, I10753, I10461;
wire I5391, g3911, I9229, g7010, g6581, g10890, g5650, g7410, g9782, g11398, I15804;
wire I16947, I5695, g10249, g2168, g2669, g6060, I16273, g2368, I11629, g11652, I9822;
wire g9661, g4198, g4747, I11472, I10736, g4398, I13451, g3733, I7444, g10248, g2772;
wire I7269, I15263, I10198, I12300, g10552, g8751, I15332, g10204, g2743, g4241, g2890;
wire g5768, I10843, g8585, I5858, g5594, I14528, g3473, g7278, I14330, g9526, I4938;
wire I8250, I11071, I15406, I15962, g2011, g6995, g7618, g3980, g8441, g11406, g5943;
wire g7343, g2411, I10132, g10786, g3069, I13776, I13785, g1982, g4524, g6294, I15500;
wire I5251, I6590, g3540, I7729, g5887, g10356, I5047, g5122, g11500, g6190, g2074;
wire g4319, g7693, g11049, I11950, I16514, g10826, I9062, g7334, g10380, g3206, I13825;
wire I13370, I9620, g4258, I16507, g4352, I11858, g11048, g4577, g4867, I14709, g5033;
wire g10233, g6156, g4717, I7014, I12511, g10182, g7555, g7804, I7414, I10087, g9919;
wire g2080, I7946, I10258, I14087, g7792, g2480, I11367, I11394, g5096, g6942, g8890;
wire g2713, I13367, I13394, g4211, g4186, g6704, I17687, g4386, g10932, I8929, g5845;
wire g4975, g2569, I7513, g8011, I17752, g5195, g5395, g5891, I9842, I17374, g7113;
wire g11106, g7313, I11420, g4426, g10897, I12916, I10069, g6954, g6250, g4170, g6810;
wire g4614, g9527, g4370, I12550, I7378, I10810, I11318, g4125, I15371, g6432, g7908;
wire I13227, g6053, I14955, I17669, g8992, g9764, I16920, g11033, g3291, I12307, I5935;
wire I6844, g6453, I9854, I14970, g4280, I7182, I7288, g4939, I11540, I5982, g3144;
wire I11058, I15795, g3344, I16121, g6568, I10171, g4083, g8080, I4879, g4544, g3207;
wire g8573, I7916, I7022, I13203, g8480, g7776, g2000, I7749, I6557, g8713, I17525;
wire g2126, g4636, I15514, I17424, g3694, g6157, I6071, I14967, I12773, I16682, I17558;
wire I15507, g5081, I12942, g3088, g5815, g8569, g4306, g7965, I12268, g5481, g11507;
wire I12156, g4790, I12655, g5692, I15421, g1964, g10387, g97, g7264, I12180, g10620;
wire g4187, g4061, g10148, g11421, g4387, g4461, I6955, g7360, g11163, g10104, I11146;
wire g4756, I17713, I13738, I13645, g8688, I12335, g7521, g10343, I14010, I14918, g8976;
wire g2608, I9829, I16760, g2220, g4427, I12930, g7450, I12993, I15473, I13290, g2779;
wire I6150, g9987, g11541, I17610, I11698, g4200, g9771, I12694, I12838, g11473, g2023;
wire I10078, I17255, g4514, I10598, g5783, g4003, g7724, I15359, I6409, g8126, I7719;
wire g5112, g7379, g5218, g8326, I17188, I17124, g5267, I17678, I11427, I12487, I15829;
wire I13427, g9892, I8039, I7752, g4763, I12502, g4191, I11632, g7878, g10850, g8760;
wire g11434, g4391, g1989, I10322, g7289, g7777, g7658, g5401, g3408, I10159, g10133;
wire g5676, g2451, I10901, g4637, I12279, I5348, g3336, I15344, g6778, g7882, g3768;
wire g10896, I13403, g11344, g4307, g4536, g10228, g4159, g2346, g4359, I12469, g6735;
wire g8183, g8608, g8924, g5830, g7611, g8220, I12286, I14561, g5727, g2103, I8919;
wire g3943, I9177, I7233, I10144, g9340, I14295, I9377, I17219, g7799, g4757, I16604;
wire I7054, I11572, g8423, g6475, g4416, g7981, g6949, g3228, g8977, g2732, I9287;
wire g9082, g10310, g8588, g7997, g2753, I12601, g6292, I11127, g4315, g4811, g2508;
wire g8361, g10379, I10966, g2240, I8004, g2072, g3433, I6921, I5279, g7332, g10050;
wire I9199, g10378, I8647, I9399, g5624, g7680, g11506, g7353, g2043, g6084, g8327;
wire I14364, g4874, g6039, g5068, I11956, g3096, I13956, I13376, I13385, I11103, g3496;
wire g7744, I11889, I17470, g7802, I5652, g8146, I5057, I11354, g2116, g8346, I5843;
wire I13354, I8503, I5989, I9510, I11824, g2034, g5677, g8103, g3395, g2434, g3337;
wire g3913, I10289, I17277, I12168, I11671, g9310, g6583, g6702, g4880, g5866, g8696;
wire I5549, I7029, I14309, g2347, I7429, g10802, g5149, I9144, I14224, g6919, I10308;
wire I12363, I7956, g7901, g4272, I8320, g10730, I12478, I12015, g6276, g11649, g9824;
wire g4243, g3266, I9259, g8240, g2914, g5198, g5747, I15491, g2210, g4417, I10495;
wire g8472, g6561, g11648, g4935, g9762, I17419, I12556, I15604, I10816, I9923, g2013;
wire g8443, g7600, I12580, g7574, I6085, g10548, I17155, g3142, g5241, g6527, I12223;
wire g4328, I14687, I17170, I14976, g8116, g3255, I7639, g8316, g3815, I11211, I10374;
wire g6764, I7109, I5909, I16534, I10643, I11088, I11024, g9556, I16098, g10317, g8565;
wire g2820, g3097, I9886, I6941, g3726, g7580, g6503, g5644, I5740, g6970, g8347;
wire I15395, g2317, I8892, g10129, g9930, I9114, g6925, I17194, I7707, g11395, g1962;
wire g10057, g2601, g10128, g5818, g8697, I6520, I14668, g4213, g11633, I11659, I12186;
wire g6120, I10195, I6031, I12953, g10323, g11191, g2775, g7076, I6812, g3783, g7476;
wire I6958, g5893, g6277, I14525, I14424, g3112, g3267, g10775, I16766, I12936, I15832;
wire I8340, I11296, g2060, g6617, I14558, g6789, I17749, I11644, I17616, I16871, I11338;
wire I13338, I9594, g4166, g11440, g4366, g5426, I15861, I16360, I6911, I13969, I7833;
wire g7285, g3329, I15247, g11573, I5525, I5710, g3761, g5614, I12762, I17704, g4056;
wire g7500, I10713, g8317, I15389, g4456, I14713, g6299, g5821, g3828, g10697, g6547;
wire I13197, g11389, g11045, I6733, I9065, I17466, g8601, g10261, g2937, g3727, g2079;
wire g5984, I10610, g10880, I15701, g4355, g11388, g7339, g2479, I10042, I15272, I16629;
wire g2840, I10189, g7024, I16220, g2190, g4260, g2390, g7795, I9433, I17642, I10678;
wire g7737, g7809, g3703, I14188, I14678, g5106, g4463, I9096, g2156, g7672, I14939;
wire g2356, g7077, g6709, I17733, g9814, g5790, I9550, I10030, g7477, I10093, I9845;
wire g3624, g6140, g6340, I5111, I11581, I11450, I12568, g9350, g10499, I5311, g3068;
wire I13714, I11315, g8784, g2942, g8739, I12242, g4279, I11707, g7205, g9773, I7086;
wire I13819, g11061, g10498, g9009, g6435, g4167, g5027, g6517, g6082, I12123, g4318;
wire g4367, I16859, g4872, g7634, I5174, I16950, g8079, I16370, g6482, I11055, g10056;
wire I9807, g8479, I7185, I12751, g9769, g4057, g5904, g7304, g5200, g10080, g8294;
wire I13978, g4457, g2163, I8877, g2363, I7070, g5446, I11590, I16172, g4193, g3716;
wire g11360, g4393, I10837, g2432, I12293, g10271, I12638, g11447, I13741, I15162, g4549;
wire I17555, I6898, I12265, g11162, g7754, g10461, g5191, g8156, I9248, g3747, I11094;
wire g1973, g5391, g8356, g10342, g3398, g6214, g7273, I5020, I6510, g9993, g10145;
wire g10031, g6110, g5637, g6310, g11629, g9822, g10199, g11451, g11472, g7044, g10887;
wire g2912, I13735, g1969, g4121, g5107, g8704, g4321, g2157, g11628, g10198, I7131;
wire I7006, g7983, I10201, g5223, I11695, g10528, g10696, g4232, I12835, I13695, g10330;
wire g5858, g10393, I10075, I7766, g8954, I16540, g6236, I6694, g7543, I12586, g11071;
wire g8363, I7487, I8237, g5416, I14494, g3119, g10132, I17519, g10869, I6088, I17176;
wire I17185, I10623, I12442, I17675, I17092, I16203, g4519, g5251, g6590, g6877, I4777;
wire g10868, g5811, g5642, g3352, I9783, g2626, g7534, g7729, g7961, g5047, I13457;
wire I10984, g9895, g6657, g10161, g4552, g4606, I15858, g8568, I8089, I10352, g6556;
wire I14352, g7927, I10822, g5874, I9001, g10259, I14418, g10708, I16739, I12430, g3186;
wire g5654, I12493, g10471, g7414, I9293, g3386, g10087, g8357, I9129, g7946, g10258;
wire g3975, I7173, I9329, I5973, g4586, g11394, g6464, g7903, g2683, I11689, I6870;
wire g3274, g3426, g5880, I12035, I13280, g2778, g10244, I9727, I7369, g3370, I10589;
wire I13624, I14194, g11420, g6563, I7920, g5272, g11319, g7036, g9085, g10069, I7459;
wire I9221, g4525, g7436, g8626, g6295, I12517, I13102, g6237, g11446, g10774, I17438;
wire I10477, I16366, g5417, g2075, I14477, g10879, I16632, g11059, g6844, g7335, g2475;
wire I14119, g1988, g3544, g2949, g7288, g11540, g5982, g10878, I7793, I10864, g3636;
wire g5629, I9953, g6089, I12193, g10171, g6731, I9068, g7805, I5655, g7916, g11203;
wire g5542, g7022, g3306, g2998, g2646, g4158, g7422, g7749, I6065, g6557, I12165;
wire I12523, g10792, g11044, g3790, I15281, g2084, g2603, I8967, g6705, g2039, I9677;
wire g3387, I10305, g5800, I5410, g3461, I15377, g6242, g2850, g9431, g7798, g11301;
wire g10459, g9812, g3756, g4587, I12475, g11377, I9866, g6948, g3622, g9958, g7560;
wire g4275, g4311, g10458, g8782, g3427, I15562, I9349, g6955, I10036, g4615, g5213;
wire g11645, I10177, I10560, I11456, I14101, I9848, I15290, g6254, g8475, g4174, g6814;
wire g9765, I17636, I15698, g10545, g2919, g7037, g10079, g10444, I9699, g6150, I14642;
wire g7437, I16784, I5667, I6395, I6891, g8292, g2952, I16956, g3345, I16376, I13314;
wire g4284, g7579, g8526, g10598, g3763, I10733, g4545, I11076, I11085, g3391, g9733;
wire I15427, I16095, g4180, g5490, g9270, g4380, g11427, g5166, I11596, g4591, I15632;
wire g11366, g3637, I7216, g7752, g11632, g8484, I16181, I10630, g8439, g2004, I10693;
wire g6836, I12372, g7917, g2986, g3307, g9473, I7671, g2647, g10159, g4420, g10125;
wire g10532, g10901, I10009, g5649, g3359, I15403, g1965, g4507, g5348, g6967, I5555;
wire I11269, g9980, g2764, I8462, g11403, g10158, g11547, g7042, I11773, g10783, g4794;
wire I11942, I13773, I5792, g7442, g8702, I13341, I12790, g7786, g2503, g3757, I9352;
wire I17312, g10353, g3416, g6993, I11180, I16190, I14485, g7364, I6815, I9717, I15551;
wire I14555, g3522, g8952, g11572, I11734, g8276, g3811, g2224, I6097, g5063, I10914;
wire g7454, I6726, I14570, I9893, I13335, g7770, I14914, g4515, g4204, I15127, I16546;
wire g8561, g2320, I10907, g7725, I8842, g7532, I7308, g3874, I8192, I12208, I8298;
wire I8085, I13965, g8004, g6921, g8986, I5494, I13131, I14239, I15956, g2617, g2906;
wire I14567, g2789, g5619, g5167, I15980, g11103, g9900, g11095, g3880, g4973, g7389;
wire g7888, g4969, g8224, g2892, g5686, g10308, g4123, g8120, g6788, g5598, g9694;
wire g10495, g2945, g11190, g8789, g9852, g5625, g4875, g9701, g7138, g10752, g11211;
wire g11024, g8547, g10669, g7707, g4884, g4839, g9870, g6640, g9650, g5687, g7957;
wire g3512, g8244, g7449, g4235, g4343, g11296, g9594, g6829, g4334, g9943, g5525;
wire g4548, g8876, g6733, g4804, g10705, g9934, g6225, g6324, g10686, g6540, g8663;
wire g11581, g6206, g4518, g3989, g7730, g5174, g7504, g7185, g2563, g7881, g11070;
wire g9859, g8877, g11590, g6199, g9266, g5545, g5180, g5591, g8556, g11094, g5853;
wire g6245, g4360, g8930, g5507, g11150, g8464, g9692, g4996, g7131, g11019, g9960;
wire g11196, g11018, g6819, g10595, g10494, g10623, g4878, g5204, g8844, g6701, g10782;
wire g5100, g4882, g8731, g6215, g6886, g3586, g8557, g8966, g8071, g11597, g9828;
wire g2918, g9830, g8955, g9592, g5123, g7059, g8254, g7459, g11102, g7718, g7535;
wire g9703, g5528, g5151, g9932, g5530, g3506, g8769, g6887, g6228, g6322, g3111;
wire g8967, g5010, g3275, g10809, g2895, g7721, g9866, g9716, g10808, g3374, g4492;
wire g8822, g10560, g11456, g9848, g4714, g6550, g5172, g10642, g3284, g9699, g9855;
wire g5618, g6891, g7940, g11085, g4736, g4968, g8837, g9644, g5804, g8462, I6330;
wire g11156, g6342, g9867, g9717, g4871, g10454, g4722, g7741, g4500, g9386, g8842;
wire g9599, g9274, g5518, g9614, g4838, g9125, g7217, g11557, g2911, g11210, g7466;
wire g9939, g11279, g10518, g4477, g8708, g7055, g5264, g6329, g6828, g8176, g6830;
wire g8005, g4099, g11601, g11187, g6746, g6221, g8765, g9622, g11143, g9904, g8733;
wire g8974, g6624, g11169, g8073, g9841, g5882, g8796, g11168, g4269, g5271, g10348;
wire g5611, g8069, g9695, g10304, g8469, g4712, g6576, g10622, g11015, g5674, g9359;
wire g9223, g11556, g9858, g5541, g4534, g6198, g6747, g6699, g6855, g3804, g5680;
wire g9642, g5744, g10333, g8399, g9447, g4903, g11178, g8510, g8245, g6319, g11186;
wire g3908, g2951, g6352, g9595, g4831, g5492, g9272, g10312, g6186, g9612, g9417;
wire g9935, g8701, g10745, g11216, g9328, g11587, g6821, g6325, g4560, g7368, g6083;
wire g6544, g5476, g7743, g4869, g5722, g6790, g8408, g10761, g7734, g8136, g6187;
wire g4752, g9902, g8768, g5500, g2496, g6756, g8972, g6622, g11639, g9366, g11230;
wire g10328, g5024, g4364, g9649, g5795, g5737, g6841, g4054, g6345, g11391, g9851;
wire g6763, g4770, I16142, g9698, g4725, g5477, g9964, g5523, g4553, g8550, g8845;
wire g2081, g6359, g11586, g11007, g5104, g5099, g6757, g5499, g4389, g6416, g9720;
wire g4990, g9619, I6630, g6047, g9652, g10515, g9843, g5273, g11465, g5044, g11237;
wire g9834, g6654, g5444, g3714, g11340, g9598, g8097, g8726, g6880, g4338, g5543;
wire g8960, g4109, g10759, g9938, g10758, g4759, g9909, g7127, g11165, g6234, g6328;
wire g8401, g11006, g4865, g4715, g4604, g5513, g11222, g4498, g6554, g7732, g9586;
wire g5178, g4584, g7472, g11253, g5182, g9860, g8703, g11600, g9710, g9645, g11236;
wire g4162, g6090, g9691, g11372, g6823, g11175, g8068, g9607, g9962, g6348, g9659;
wire g9358, g3104, g4486, g9587, g5632, g9111, g4881, g11209, g8848, g4070, g6463;
wire g8699, I5689, g7820, g11021, g5917, g6619, g6318, g6872, g11320, g10514, g4006;
wire g9853, g11274, g6193, g8119, g9420, g5233, g7581, g6549, g11464, g4801, g6834;
wire g4487, g2939, g7060, g5770, g5725, g11641, g2544, g11292, g5532, g11153, g9905;
wire g7739, g6321, g8386, g8975, g2306, g6625, g7937, g10788, g10325, g8170, g5706;
wire g2756, g8821, g10946, g4169, g5029, g11164, g4007, g4059, g4868, g5675, g4718;
wire g10682, g6687, g7704, g4582, g4261, g3422, g5745, g8387, g7954, g11283, g8461;
wire g10760, g11492, g7032, g8756, g9151, g6341, g10506, g9648, g7453, g6525, g6645;
wire g5707, g8046, g11091, g11174, g9010, g8403, g5201, g8841, g6879, g8763, g4502;
wire g9839, g6358, g5575, g4940, g8107, g10240, g11192, g9618, g5539, g8416, g9693;
wire g11553, g8047, g5268, g9555, g6180, g6832, g10633, g7894, g8654, g9621, g6794;
wire g9313, g4883, g3412, g7661, g2800, g3389, g3706, g9908, g3429, g6628, g5470;
wire g7526, g5897, g5025, g6204, g4048, g8935, g3281, g9593, g4827, g10701, g10777;
wire g8130, g9965, g3684, g11213, g5006, g9933, g8554, g9641, g6123, g6323, g10766;
wire g6666, g4994, g5755, g11592, g6351, g6875, g4816, g9658, g6530, g8366, g9835;
wire g6655, g5445, g5173, g7970, g3098, g5491, g9271, g11152, g9611, g6410, g10451;
wire g4397, g7224, g5602, g4421, g6884, g6839, g8698, g8964, g8260, g11413, g4950;
wire g5535, g7277, g8463, g3268, g10785, g6618, g6235, g10950, g4723, g8720, g6693;
wire g11020, g11583, g8118, g8167, g6334, g7892, g8652, g5721, g10367, g9901, g6792;
wire g11282, g7945, g8971, g11302, g4585, g6621, g5502, g11105, g7709, g8598, g7140;
wire g9600, g9864, g11640, g5188, g7435, g7876, g5030, g4058, g6776, g4890, g2525;
wire g10301, g4505, g9623, g10739, g11027, g10738, g8687, g6360, g9871, g5108, g11248;
wire g4992, g11552, g9651, g11204, g7824, g4480, g6179, g8710, g7590, g9384, g3407;
wire g9838, g3718, g10661, g11380, g8879, g7930, g8962, g10715, g8659, g3015, g9643;
wire g9205, g5538, g4000, g4126, g4400, g2794, g4760, g6238, g10784, g8174, g6332;
wire g5067, g5418, g10297, g6353, g11026, g11212, g6744, g5493, g10671, g4383, g5256;
wire g4220, g8380, g7071, g4779, g9613, g7705, g9269, g5181, g4977, g7948, g11149;
wire g9862, g11387, g7955, g4161, g11148, g9712, g8931, g11097, g5421, g11104, g5263;
wire g6092, g4999, I6338, g7409, g4103, I6309, g6580, g5631, g9414, g9660, g9946;
wire g5257, g4732, g3108, g4753, g9903, g10625, g5605, g6623, g11228, g11011, g6889;
wire g8040, g7822, g8123, g11582, g4316, g10969, g5041, g9335, g9831, g4565, g9422;
wire g8648, g8875, g5168, g7895, g8655, g3396, g4914, g9947, g5772, g6838, g5531;
wire g6795, g10503, g8010, g8410, g6231, g10581, g10450, g2804, g3418, g4820, g9653;
wire g6205, g10818, g8172, g10496, g5074, g9869, g9719, g10741, g3381, g5863, g8693;
wire g5480, g4581, g3685, g5569, g8555, g3263, g9364, g4784, g9454, I6331, g11299;
wire g6983, g7958, g4995, g4079, g2264, g2160, g3257, g3101, g5000, g3301, g5126;
wire I5084, g9412, g9389, g2379, g10706, I16145, g10597, g8965, g5608, g5220, g10624;
wire g10300, g5023, g4432, g4053, g8050, g5588, g6679, g9963, g3772, g5051, g6831;
wire g2981, g8724, g4157, g9707, g8878, g2132, g10763, g8289, g7898, g11271, g11461;
wire g5732, g11145, g11031, g9865, g5944, g9715, g9604, g8799, g11198, g6873, g6632;
wire g6095, g3863, g9833, g6653, g6102, g7819, g11393, g2511, g7088, g9584, g9896;
wire g8209, g6752, g4778, g11161, g9268, g5681, g7951, g9419, g10268, g5533, g9052;
wire g6786, g10670, g11087, g4949, g6364, g7825, g3400, g4998, g10667, g7136, g6532;
wire g9385, I5690, g4484, g9897, g9425, g3383, g5601, g7943, g11171, g3423, g7230;
wire g4952, g8736, g6787, g8968, g10306, g9331, g11459, g4561, g11425, g11458, g5739;
wire g7496, g4986, g11010, g3999, g8175, g8722, g4764, g7137, g7891, g8651, g5479;
wire g11599, g6684, g6745, g6639, g10937, g3696, g4503, g6791, g5190, g5390, g8384;
wire g4224, g5501, g9173, g6759, g8838, g8024, g10666, g11158, g9602, g5704, g4617;
wire g11561, g9868, g11295, g11144, g9718, g3434, g4987, g4771, g5250, g6098, g9582;
wire g6833, g3533, g4892, g8104, g9415, g8499, g9664, g10740, g2534, g8754, g9721;
wire g6162, g4991, g6362, I6631, g10685, g4340, g11023, g8044, g11224, g11571, g4959;
wire g10334, g5626, g9940, g4876, g6728, g6730, g9689, g10762, g6070, g9428, g9030;
wire g9430, g8927, g7068, g8014, g11392, g5782, g9910, g4824, g6331, g4236, g11559;
wire g9609, g11558, g6087, g4877, g5526, g10751, g10772, g8135, g11544, g5084, g8382;
wire g10230, g5484, g7241, g3942, g10638, g4064, g9365, g9861, g8749, g11255, g11189;
wire g10510, g8947, g2917, g5919, g11188, g9846, g7818, g11460, g5276, g11030, g11093;
wire g7893, g8653, g10442, g6535, g8102, I5085, g5004, g3912, g7186, g4489, g9662;
wire g9418, g11218, g4471, g10746, g7125, g7821, g6246, g9256, g8042, g10237, g7939;
wire g8786, g10684, g11455, g8364, g2990, g9847, g8054, g5617, g6502, g5789, g4009;
wire g11277, g6940, g7061, g11595, g5771, g8553, g4836, g5547, g6216, g4967, g6671;
wire g7200, g3661, g7046, g4229, g8389, g6430, g8706, g4993, g6247, g9257, g11170;
wire g7145, g5738, g6826, g7191, g3998, g6741, g5478, g11167, g11194, g11589, g6638;
wire g4921, g7536, g9585, g2957, g11588, g5690, g6883, g4837, g8963, g8791, g6217;
wire I6316, g11022, g5915, g4788, g8759, g5110, g11254, g6827, g8957, g6333, g8049;
wire g4392, g9856, g9411, g5002, g11101, g11177, g11560, g8098, g3970, g4941, g10453;
wire g5877, g6662, g7935, g6067, I6317, g9863, I5886, g6994, g9713, g4431, g4252;
wire g11166, g7130, g11009, g7542, g8019, g11008, g3516, g8052, g3987, g4765, g11555;
wire g9857, g8728, g8730, g8185, g5194, g8385, g4610, g7902, g4073, g8070, g5731;
wire g11238, g4473, g8470, g5489, g3991, I5887, g7823, g4069, g11519, g11176, g11092;
wire g11154, g9608, g11637, g2091, g8406, g5254, g7260, g5150, g8766, g9588, g8801;
wire g7063, g10303, g5009, g9665, g8748, g11215, g10750, g5769, g8755, g6673, g5212;
wire g7720, g5918, g8045, g8173, g11349, g7843, g9696, g6772, g6058, g6531, g6743;
wire g6890, g7549, g8169, g11304, g9944, g9240, g8059, g8718, g8767, g9316, g7625;
wire g8793, g2940, g4114, g11636, g10949, g4870, g3563, g10948, g8246, g5788, g4008;
wire g9596, g5249, g11585, g3089, g4972, g11554, g7586, g10673, g4806, g5485, g9936;
wire g2910, g9317, g10933, g8388, g4465, g7141, g10508, g4230, g10634, g9601, g6126;
wire g6326, g7710, g8028, g6760, g5640, g5031, g4550, g7879, g7962, g9597, g10452;
wire g4891, g5005, g6423, g8108, g4807, g5911, g9937, g9840, g10780, g8217, g11013;
wire g9390, g11214, g6327, g4342, g5796, g5473, g6346, g6633, g11005, g8365, g8048;
wire g4481, g4097, g8055, g4497, g9942, g6696, g10731, g8827, g5540, g4960, g8846;
wire g6508, g6240, g7931, g5287, g6472, g11100, g11235, g5199, g6316, g7515, g10583;
wire g5781, g8018, g4401, g8994, g2950, g5510, g6347, g9357, g4828, g11407, g4727;
wire g10357, g10743, g5259, g5694, g10769, g11584, g4932, g10768, g6820, g4068, g6317;
wire g5215, g4576, g4866, g6775, g3829, g10662, g8101, g5825, I6310, g7884, g5008;
wire g3974, g9949, g2531, g9292, g10778, g8041, g6079, g7235, g9603, g6840, g9850;
wire g7988, g5228, g7134, g5934, g5230, g8168, g9583, g10672, g3287, g8772, g4893;
wire g10331, g8505, g10449, g11273, g8734, g5913, g10448, g6163, g6363, g7202, g11463;
wire g8074, g4325, g8474, g11234, g5266, g4483, g5248, g11514, g5255, g4106, g2760;
wire g5097, g5726, g5497, g5354, g7933, g9617, g9906, g11012, g7050, g10971, g4904;
wire g10369, g8400, g4345, g2161, g5001, g9945, g7271, g9709, g4223, g10716, g11291;
wire g6661, g11173, g6075, g8023, g9907, g10582, g5746, g5221, g9959, g7674, g9690;
wire g6627, g5703, g4522, g4115, g7541, g10627, g4047, g6526, g2944, g6646, g7132;
wire g11029, g8051, g8127, g7209, g11028, g6439, g10742, g9110, g10681, g4537, g9663;
wire g5349, g8732, g3807, g8753, g5848, g8508, g8072, g5699, g11240, g5398, g6616;
wire g10690, g8043, g9590, g4128, g6404, g6647, g10504, g9657, g4542, g4330, g3497;
wire g5524, g8147, g4554, g9899, g5258, g7736, g6224, g10626, g6320, g7623, g10299;
wire g7889, g10298, g8413, g3979, g4902, g5211, g4512, g7722, g9844, g4490, g4823;
wire g6516, g5026, g8820, g10737, g8936, g10232, g6771, g5170, g8117, g4529, g4348;
wire g9966, g5280, g7139, g11099, g6892, g9705, g10512, g11098, g8775, g5083, g5544;
wire g11272, g5483, g9948, g4063, g11462, g6738, g8060, g6244, g11032, g10445, g9150;
wire g10316, g5756, g4720, g9409, g8995, g6876, g4989, g9836, g6656, g5514, g8390;
wire g5003, g9967, g5145, g4834, g4971, g10753, g5695, g7613, g10736, g11220, g7444;
wire g5536, g6663, g4670, g6824, g4253, g8250, g8163, g10764, g5757, g10365, g8032;
wire g11591, g8053, g11147, g5522, g5115, g9837, g9620, g11151, g11172, g7885, g6064;
wire g8929, g5595, g5537, g9842, g4141, g4341, g9192, g7679, g7378, g5612, g3939;
wire g7135, g10970, g11025, g9854, g7182, g9941, g6194, g5128, g4962, g4358, g8683;
wire g4506, g6471, g8778, g11281, g8735, g11146, g3904, g8075, g9829, g8949, g7632;
wire g11290, g6350, g10599, g5902, I6337, g2276, g6438, g5512, g5090, g7719, g2561;
wire g3695, g8603, g8039, g9610, g3536, g5529, g5148, g9124, g9324, g4559, g10561;
wire g5698, g11226, g10295, g5260, g10680, g6822, g4905, g11551, g3047, g9849, g5279;
wire g8404, g5720, g5318, g8764, g11376, g11297, g9898, g6895, g7189, g9510, g7297;
wire g9088, g9923, g6485, g8771, g5813, g7963, g10643, g9886, g9951, g11625, g8945;
wire g10489, g10559, g10558, g11338, g8435, g10544, g6911, g10865, g3698, g8214, g6124;
wire g6469, g5587, g6177, I14585, g9891, g9913, I5600, g11257, g8236, g7385, g6898;
wire g6900, g4264, g9726, g6088, g6923, g8194, g9676, g11256, g3860, g11280, g9727;
wire g4997, g11624, g11300, g4238, g8814, g10401, g8773, g11231, g10864, g9624, g9953;
wire g6122, g6465, g6934, g7664, g7246, g7203, g6096, g9747, g11314, g10733, g8921;
wire I15054, g11269, g5555, g11268, g10485, g10555, g6481, g10712, g11335, g8249, g7638;
wire g10567, g11487, I15210, I5805, g8941, g11443, g4231, g11278, I15039, g11286, g8431;
wire g7133, g11306, g8252, g8812, g7846, g3875, g5996, g6592, g8286, g10501, g10728;
wire g8270, g7290, g6068, g6468, g11217, g11478, g9536, g5981, g11486, g8377, g8206;
wire g11580, g8287, g11223, g9522, g8199, g5802, g11321, g6524, g10664, g7257, g7301;
wire g10484, g10554, g8259, g11334, g8819, g8923, g8488, g7441, g6026, g10799, g10798;
wire g10805, g10732, g6061, g9512, g10013, g8806, g8943, g11293, g11265, g8887, g5838;
wire g6514, g8322, g8230, g5809, g8433, g11579, g10771, g11615, g9367, g9872, g6522;
wire g8266, g10414, g11275, g11430, g8248, g9686, g8815, g7183, g5983, g8154, g6537;
wire g4309, g10725, g6243, I6351, g9519, g9740, g8267, g10744, g6542, g7303, g10652;
wire g5036, g7240, g8221, g6902, I14776, g10500, g4052, I14858, g6529, g11264, I15209;
wire g8241, g10795, g11607, g8644, g4682, g8818, g2984, g9931, g3414, g9515, g10724;
wire g7294, g5189, g8614, g3513, g6909, I5571, g4283, g8939, g2514, g11327, g8187;
wire g11606, g11303, g5309, g9528, g8200, g2522, g2315, g6506, g10649, g8159, g7626;
wire g10770, g9566, g11483, g8811, g8642, g6545, g10767, g11326, g10898, g11252, g10719;
wire g4609, g6507, g10718, g10521, g7075, g7292, g10861, g8417, g6515, I14855, I15205;
wire I15051, g9724, g6528, g8823, g7503, g8148, g8649, g3584, g10776, g9680, g10859;
wire I14866, g7299, g10858, g8193, g9511, g7738, g7244, g3425, g7478, g9714, g10025;
wire g6908, g5028, g8253, g8938, g8813, g9736, g9968, g8552, g5910, g11249, g11482;
wire g9722, I15204, g7236, I14596, g8645, g11647, g6777, g9737, I16149, g11233, g8607;
wire I16148, g8158, g5846, g5396, g5803, g11331, g7295, g6541, g8615, g9742, g9926;
wire g9754, g8284, g2204, g7471, g7242, g5847, g6901, g8559, g9729, g10860, g9927;
wire g10497, g9885, g2528, g11229, g8973, g10658, g10339, I5363, g11310, g6500, g10855;
wire g9916, g10411, g11603, I5357, g9560, g6672, g9873, g6523, g10707, I5626, g9579;
wire g7298, g6551, g6099, g8282, g9917, I15057, g7219, g10019, g5857, g9725, g11298;
wire g10402, g2521, I14751, g10866, g6534, g11232, g9706, g10001, g8776, g7225, g9888;
wire g11261, g9956, g10923, g8264, g6513, I14835, g8641, g5361, g11316, I16161, g6916;
wire g8777, g2353, g7510, g9957, g2744, g7245, g7291, g8611, I15199, g10550, g11330;
wire g10721, g8153, g10773, g3688, I15225, g6042, g10655, g11259, g11225, g5914, g11258;
wire g6054, g9728, g9730, g5820, g8574, g11602, g10502, g10557, I15171, g11337, g7465;
wire g8262, g8889, g7096, g5995, g8285, g10791, g2499, I14607, g6049, g9920, g10556;
wire g8643, g5810, g11336, g8742, g8926, g7218, I15224, g7293, g11288, g10800, g11308;
wire g8269, g10417, g10936, g9388, g6185, g6470, g6897, g8885, g11260, g11488, g6105;
wire g10807, g10639, g4556, g8288, g6755, I14862, I16160, I15042, g11610, g9711, g6045;
wire g11270, g7258, g6059, g10007, g11267, g11294, g9509, g7211, g5404, g4089, I15219;
wire g11219, g6015, g10720, g8265, g5224, g9700, g7106, g8770, g11201, g9950, g9723;
wire g2309, g11266, g10727, g10863, g8429, g9751, g8281, g6910, g8639, g9673, g11285;
wire g11305, I15177, g9734, I14827, g5824, g8715, g5762, g6538, g5590, g10726, g3120;
wire g9573, g4640, g6093, g8162, g8268, g9569, g11485, g10797, I14779, g10408, g10635;
wire g2305, I15176, g3435, g9924, g10711, g5814, g5038, I15215, g8226, g7367, g7457;
wire g5229, g5993, g8283, g7971, g8602, g8920, g10663, g6074, g8261, g10862, g5837;
wire g11333, g6080, g6480, g7740, g10702, g9697, g8203, g9914, g10564, g11484, g5842;
wire I15200, g11609, I14582, g8940, g11312, g11608, g6000, g8428, g8430, g9922, g8247;
wire g3438, I5576, g6924, g5405, g8638, g8609, g9995, g8883, I15214, g2538, g11329;
wire g4255, g11328, g9704, I5352, g8774, g9954, g10405, g9363, g5849, I5599, g7204;
wire g7300, g4293, g9912, g6533, g8816, g9929, g5819, I14831, g5852, g8263, g3431;
wire g9683, g8631, g6922, g8817, g9735, g8605, g11263, g6739, g11332, g7143, g6479;
wire I15048, g6501, g9702, g11221, g9952, g11613, g7621, g3399, g11605, g4274, I14602;
wire I15033, g10717, I5629, g9925, g3819, g6912, g10723, g6929, g10646, g9516, g6626;
wire I6350, g11325, I5366, I5649, g6894, g9738, g8383, g8779, g8161, g8451, g9915;
wire g2316, g5576, g10857, g10793, g7511, g8944, g10765, g10549, g7092, g11604, g8434;
wire g6546, g3354, g9928, g11262, g9785, g5867, g8210, g10533, g9563, g6906, g7375;
wire g7651, I5570, g9731, g11247, I15045, g10856, g9557, g7184, g11612, g7384, g11324;
wire g8922, I5358, g9955, g2501, g7231, g6078, g6478, g6907, g6035, g8937, g7742;
wire g10722, g9918, g5403, g7926, g6915, g5841, I15220, g10529, g11246, g6002, g7712;
wire g8810, g9921, g8432, I15172, I14822, g6928, g8157, g6930, g7660, g6899, g9392;
wire g11318, I16427, g11227, g11058, I5351, g9708, g6071, g9911, g7102, g7302, g6038;
wire g4239, g8646, g9974, g5823, g6918, g7265, I5804, g5851, g11481, g10336, g7296;
wire g4300, g8647, g8546, g2516, g2987, I5593, g8970, I10519, I11279, g7990, I11278;
wire g3978, I5264, I8640, I6761, I17400, I5450, I16060, I6746, I11975, I12136, I11937;
wire g2959, I5878, g2517, g5552, I6468, I8796, g10392, I5611, g8738, I6716, g2310;
wire I7685, g3056, I12108, g3529, I6747, g2236, g7584, I15870, I16067, I7562, I13531;
wire I8797, I17584, I11936, I15257, g8402, g8824, I6186, g11496, I16001, I6125, I11909;
wire I12040, I13909, g3625, I11908, g10470, I13908, g3813, I8650, g6207, I16066, g2948;
wire I11242, g10467, I6187, g6488, I5500, I11974, I12062, g5300, I5184, I13293, I6200;
wire I13265, I5024, I7863, g8705, g8471, I15256, I6145, I13992, I11510, g10853, I5231;
wire I12047, I10771, g10477, g7582, I5104, g8409, I6447, I4956, I5613, I8481, g5278;
wire I6880, I15431, g5548, g7671, I12020, g10665, I16469, I5014, I13523, I16039, I16468;
wire I12046, g4476, g10476, I16038, I8676, I12113, I8761, g3204, I15993, I5036, I14263;
wire g8298, I5135, g2405, I7034, I15443, I6166, I8624, I16015, I8677, I8576, I14613;
wire I8716, g3530, g8405, g4104, I12003, g2177, g3010, g5179, I17395, g7067, g7994;
wire I6167, I5265, I6989, I13274, I10507, I13530, I5164, g9107, I9559, I8577, g2510;
wire g8177, I8717, I5296, g5209, g7950, g2088, I16000, I5371, g2215, g7101, I5675;
wire I8544, g6577, I5297, I13537, I13283, g4749, I11982, I8514, I13091, g2943, I15908;
wire I6879, I8763, I5449, g8825, I16007, I5865, I5604, g2433, I6111, g2096, I13522;
wire I10770, g6027, g7992, I5539, I17394, I13553, I8642, g7573, g11416, g6003, g8934;
wire I15992, I7683, I4910, g3209, I6794, I10521, I5486, I15442, g6858, I5185, g5304;
wire g2354, I15615, I17281, I5470, I11509, I5025, I11508, I15430, I14612, g4675, I14272;
wire g2979, I17290, g5269, g4297, I12002, I5006, I12128, I5105, I6323, g7588, I6666;
wire g3623, I5373, I8529, I5283, I7224, I5007, I5459, I17297, g8746, I6143, I5015;
wire g8932, I16073, I6988, g3205, I8652, I9558, I5203, g7533, g3634, I6792, g3304;
wire I12145, g7596, I13302, I5502, I9574, g3273, I8670, I7035, I15453, I8625, I7876;
wire I14203, I15607, g2274, I8740, I17296, g10507, g2325, I8606, I12087, I13249, I13248;
wire I13552, g2106, I12069, g9204, I12068, I17503, I7877, I5165, g6740, I6289, I6777;
wire g5171, I15891, I13090, g11474, g7942, I5538, I7563, I13513, g2107, g2223, I13505;
wire I6209, I12086, I8545, I8180, g2115, I8591, I10931, I17402, g8307, I12144, I10520;
wire I5263, g8757, I6714, I14211, I8515, g2272, I9946, I8750, I5605, g8880, I16051;
wire I16072, g10440, g8612, I15872, I8528, g8629, g8542, I9947, I6838, g7583, g4803;
wire I17307, g4538, I15452, I13857, I14202, I13765, g2260, g7986, g5226, g8512, I16046;
wire I13504, g10447, g2167, I8804, g10472, I17487, I4995, I12093, g7987, g5227, I5126;
wire g2321, g7547, I17306, g6548, I11995, I7225, I11261, g8843, g2938, I4942, g10394;
wire g8549, g3070, I4954, I5023, g10446, I16081, I8641, I6178, I12075, I5127, I5451;
wire g4168, I6288, I8179, I4912, I6805, g3766, g3087, I17486, I4929, I15890, I16331;
wire I9575, I13887, g5308, I13529, I6208, g5217, I5316, g2111, g10366, I5034, I13869;
wire I13868, I15999, I13259, g3261, g10481, g2180, g4976, g8506, g2380, I13258, I5013;
wire g5196, I10930, I6770, g11449, g11448, I15717, I5317, I14210, I17569, I13878, g8545;
wire g2515, I14443, g7557, g8180, I14279, I17568, I13886, I7322, I6990, I14278, I7033;
wire I9006, g8507, I5460, g4588, I4986, g3247, I8651, I13545, g8628, I6138, I12074;
wire g8630, I13078, I6109, g8300, I5501, I17586, I12092, I13901, I8795, I6201, I14217;
wire I9007, I13561, I15716, I6449, I13295, I4987, I6715, I17493, I12215, g2372, g7062;
wire g2988, I13309, g8839, g2555, g3662, I13308, g2792, g4117, I8543, g11549, I6881;
wire I12138, I8729, I14216, g10384, I13260, g2776, I8513, I13559, I8178, g3631, I6487;
wire I16080, I13893, I12115, I6748, I13544, I5484, I4928, I6226, I8805, I4930, I15880;
wire I14265, I16031, g3585, g3041, g8933, I16330, I13267, I13294, g10231, I14442, I6793;
wire I4966, I8752, I15432, I12214, g10511, g3011, g5103, I16087, g3734, I6664, g8882;
wire I4955, I8786, g3992, g10480, I11915, I8770, I5516, g8541, I6188, g5147, g8744;
wire I5892, g8558, I15258, I13266, I8787, I6826, I17283, g5013, I17492, g8511, I16079;
wire I5035, I5517, I7223, I16086, g5317, I15879, I15878, I12114, I12107, g2500, I15994;
wire g7934, g10469, I14264, I6448, I13285, g10468, I6827, g8623, I13900, g2795, I8575;
wire I14209, I13560, I8715, I8604, I16017, I4941, g2205, g3753, I6467, I14614, g2104;
wire g2099, I16023, g10479, g8737, g5942, g10478, I12004, I4911, I11914, g7960, I5295;
wire I12106, I8728, g3681, I11907, I13907, I8730, g8551, I4980, g2961, g6019, I16016;
wire I11935, I8678, I17051, g4482, g7592, g3460, g7932, g7624, g7953, g8414, I6168;
wire I5229, I6772, I16030, I13284, I16065, g2947, I7321, g2437, g2102, I17282, I5620;
wire I8664, g7524, g7717, I16467, I4972, I13554, I16037, g8302, I4943, I5485, g5527;
wire I10509, g7599, I10508, I6126, I8671, I6760, g3626, I11973, g2389, I15617, g5277;
wire I5005, I6779, I6665, I8589, g8412, g2963, I12045, I16053, g2109, g11418, I13539;
wire g10475, I5324, I13538, I5469, I5540, I17505, I11241, I8803, I12061, I8780, g8745;
wire I4979, g8109, g8309, g6758, I16009, I15616, I8662, I16008, I13515, I13991, g11276;
wire I15900, g2419, I16074, I10769, I7323, g7978, I7875, I8562, I15892, g3771, I8605;
wire g10153, g5295, I8751, I15907, I5136, I11263, I14204, g8881, g2105, g5557, I5230;
wire I8669, g10474, I8772, g2445, g8006, I10932, I17504, I5137, g8305, I5891, I13273;
wire I8480, g4144, I15906, I5342, I13514, g8407, g4088, g4488, g7598, g3222, I16052;
wire I12127, g10483, g8415, g11415, g6573, I5676, I6778, g9413, I8779, I5592, g8502;
wire I15609, I15608, g3071, g10509, I17461, I13506, I5468, g5219, I5677, g8826, I17393;
wire I5866, I12126, I4978, g7587, g5286, g8308, I7864, I11981, I12060, g5225, g11538;
wire I13767, g10396, I11262, I13990, I6224, I5867, g2493, I5893, g3062, I13521, I5186;
wire I6771, I5325, I17459, I9557, g11414, I12067, I12094, I4964, I13272, I9948, g10302;
wire I16332, I5106, g8847, g2257, I12019, I15441, I11997, I8739, I5461, I13766, I8479;
wire I17295, I14271, I4971, g8301, I6110, g10482, g10779, I6762, I17289, I5315, I17288;
wire I13859, g7548, I13858, I11996, g8743, I5880, g10513, g8411, I8626, g10505, I5612;
wire g4821, I12076, I12085, g7567, I5128, I6489, g7593, I8778, g10149, I13902, I13301;
wire g3215, g7996, I4985, I14444, g8000, I5166, I17460, g3008, I6836, I5529, g10229;
wire I13661, I13895, g2303, I12039, g5592, I12038, g3322, I8561, I8527, I12143, I5619;
wire g10386, I11980, I6837, I4973, I13888, g7558, I17494, g11491, I16045, I7684, g4130;
wire I8771, I13546, I13089, g2117, g5119, g5319, I15899, I5606, I15898, I16032, I17401;
wire I13659, I8738, I13250, I15718, I9008, I6176, I7865, g5274, I5341, I17305, I17053;
wire g5125, I12216, I6225, I5879, g3221, I14270, I6124, I6324, I13867, I13894, I6469;
wire I8663, g7523, I6177, g5187, I6287, I8762, I15871, g8840, g2250, I8590, I6199;
wire I14218, g8190, I5284, I17485, I4965, I5591, g8501, I15451, g8942, I13877, g7269;
wire I4996, I6144, I17567, g7572, I6207, I14277, I16059, I16025, I8563, g3524, I16058;
wire I5204, I6488, g3818, I16044, g3717, I13077, g10043, I11280, I6825, I4997, I13300;
wire I5323, I6136, g5935, I5528, I6806, I5530, g10886, g3106, I13876, I6322, g3061;
wire g2439, g7947, I9576, I13660, g3200, g4374, I11916, I5372, g3003, g8627, I5618;
wire I6137, I5343, I5282, I13307, I13076, I6807, I11243, I17585, I12137, I7564, g2970;
wire g10144, I8788, g7054, I17052, g2120, g8616, I5202, I16088, I16024, g11490, I5518;
wire g5118, I12021, g6392, g5938, g2478, g10374, g4278, g10424, g10383, g3118, g9815;
wire g11077, g9746, g3879, g10285, g11480, g4076, g10570, g10239, g10594, g9426, g10382;
wire g4672, g5360, g9387, g10438, g4613, g9391, g4572, g9757, g9416, g9874, g9654;
wire g9880, g4873, g2807, g10441, g4639, g10435, g10849, g9606, g9879, g9506, g6155;
wire g6355, g9615, g10371, g9591, g10359, g10434, g10358, g9750, g10291, g4227, g9655;
wire g9410, g9667, g10563, g9776, g10324, g4455, g9878, g10360, g9882, g10370, g4605;
wire g10420, g10562, g10427, g5780, g10385, g10376, g10426, g4601, g5573, g9808, g5999;
wire g9759, g6037, g10287, g5034, g9362, g9881, g10443, g10286, g4276, g4616, g10363;
wire g2862, g10373, g10423, g9758, g9589, g9803, g10430, g9421, g10362, g2791, g9817;
wire g9605, g10372, g9669, g10422, g10436, g5556, g4286, g4974, g9779, g9423, g5350;
wire g9361, g2459, g10381, g4259, g10522, g5392, g4122, g6023, g3462, g4218, g4267;
wire g4677, g9646, g2863, g9616, g6032, g9647, g5859, g10433, g10368, g4251, g9876;
wire g9656, g8303, g10429, g10428, g4234, g9877, g5186, g9489, g4619, g10432, g5345;
wire g5763, g10375, g4879, g4607, g10425, g3107, g10322, g4630, g10364, g9781;
wire line1, line2, line3, line4, line5, line6, line7, line8, line9, line10, line11;
wire line12, line13, line14, line15, line16, line17, line18, line19, line20, line21, line22;
wire line23, line24, line25, line26, line27, line28, line29, line30, line31, line32, line33;
wire line34, line35, line36, line37, line38, line39, line40, line41, line42, line43, line44;
wire line45, line46, line47, line48, line49, line50, line51, line52, line53, line54, line55;
wire line56, line57, line58, line59, line60, line61, line62, line63, line64, line65, line66;
wire line67, line68, line69, line70, line71, line72, line73, line74, line75, line76, line77;
wire line78, line79, line80, line81, line82, line83, line84, line85, line86, line87, line88;
wire line89, line90, line91, line92, line93, line94, line95, line96, line97, line98, line99;
wire line100, line101, line102, line103, line104, line105, line106, line107, line108, line109, line110;
wire line111, line112, line113, line114, line115, line116, line117, line118, line119, line120, line121;
wire line122, line123, line124, line125, line126, line127, line128, line129, line130, line131, line132;
wire line133, line134, line135, line136, line137, line138, line139, line140, line141, line142, line143;
wire line144, line145, line146, line147, line148, line149, line150, line151, line152, line153, line154;
wire line155, line156, line157, line158, line159, line160, line161, line162, line163, line164, line165;
wire line166, line167, line168, line169, line170, line171, line172, line173, line174, line175, line176;
wire line177, line178, line179, line180, line181, line182, line183, line184, line185, line186, line187;
wire line188, line189, line190, line191, line192, line193, line194, line195, line196, line197, line198;
wire line199, line200, line201, line202, line203, line204, line205, line206, line207, line208, line209;
wire line210, line211, line212, line213, line214, line215, line216, line217, line218, line219, line220;
wire line221, line222, line223, line224, line225, line226, line227, line228, line229, line230, line231;
wire line232, line233, line234, line235, line236, line237, line238, line239, line240, line241, line242;
wire line243, line244, line245, line246, line247, line248, line249, line250, line251, line252, line253;
wire line254, line255, line256, line257, line258, line259, line260, line261, line262, line263, line264;
wire line265, line266, line267, line268, line269, line270, line271, line272, line273, line274, line275;
wire line276, line277, line278, line279, line280, line281, line282, line283, line284, line285, line286;
wire line287, line288, line289, line290, line291, line292, line293, line294, line295, line296, line297;
wire line298, line299, line300, line301, line302, line303, line304, line305, line306, line307, line308;
wire line309, line310, line311, line312, line313, line314, line315, line316, line317, line318, line319;
wire line320, line321, line322, line323, line324, line325, line326, line327, line328, line329, line330;
wire line331, line332, line333, line334, line335, line336, line337, line338, line339, line340, line341;
wire line342, line343, line344, line345, line346, line347, line348, line349, line350, line351, line352;
wire line353, line354, line355, line356, line357, line358, line359, line360, line361, line362, line363;
wire line364, line365, line366, line367, line368, line369, line370, line371, line372, line373, line374;
wire line375, line376, line377, line378, line379, line380, line381, line382, line383, line384, line385;
wire line386, line387, line388, line389, line390, line391, line392, line393, line394, line395, line396;
wire line397, line398, line399, line400, line401, line402, line403, line404, line405, line406, line407;
wire line408, line409, line410, line411, line412, line413, line414, line415, line416, line417, line418;
wire line419, line420, line421, line422, line423, line424, line425, line426, line427, line428, line429;
wire line430, line431, line432, line433, line434, line435, line436, line437, line438, line439, line440;
wire line441, line442, line443, line444, line445, line446, line447, line448, line449, line450, line451;
wire line452, line453, line454, line455, line456, line457, line458, line459, line460, line461, line462;
wire line463, line464, line465, line466, line467, line468, line469, line470, line471, line472, line473;
wire line474, line475, line476, line477, line478, line479, line480, line481, line482, line483, line484;
wire line485, line486, line487, line488, line489, line490, line491, line492, line493, line494, line495;
wire line496, line497, line498, line499, line500, line501, line502, line503, line504, line505, line506;
wire line507, line508, line509, line510, line511, line512, line513, line514, line515, line516, line517;
wire line518, line519, line520, line521, line522, line523, line524, line525, line526, line527, line528;
wire line529, line530, line531, line532, line533, line534;
DFFX1 gate1(.Q (g1289), .QB (line1), .D(g5660), .CK(clk));
DFFX1 gate2(.Q (g1882), .QB (line2), .D(g9349), .CK(clk));
DFFX1 gate3(.Q (g312), .QB (line3), .D(g5644), .CK(clk));
DFFX1 gate4(.Q (g452), .QB (line4), .D(g11257), .CK(clk));
DFFX1 gate5(.Q (g123), .QB (line5), .D(g8272), .CK(clk));
DFFX1 gate6(.Q (g207), .QB (line6), .D(g7315), .CK(clk));
DFFX1 gate7(.Q (g713), .QB (line7), .D(g9345), .CK(clk));
DFFX1 gate8(.Q (g1153), .QB (line8), .D(g6304), .CK(clk));
DFFX1 gate9(.Q (g1209), .QB (line9), .D(g10873), .CK(clk));
DFFX1 gate10(.Q (g1744), .QB (line10), .D(g5663), .CK(clk));
DFFX1 gate11(.Q (g1558), .QB (line11), .D(g7349), .CK(clk));
DFFX1 gate12(.Q (g695), .QB (line12), .D(g9343), .CK(clk));
DFFX1 gate13(.Q (g461), .QB (line13), .D(g11467), .CK(clk));
DFFX1 gate14(.Q (g940), .QB (line14), .D(g8572), .CK(clk));
DFFX1 gate15(.Q (g976), .QB (line15), .D(g11471), .CK(clk));
DFFX1 gate16(.Q (g709), .QB (line16), .D(g8432), .CK(clk));
DFFX1 gate17(.Q (g1092), .QB (line17), .D(g6810), .CK(clk));
DFFX1 gate18(.Q (g1574), .QB (line18), .D(g7354), .CK(clk));
DFFX1 gate19(.Q (g1864), .QB (line19), .D(g7816), .CK(clk));
DFFX1 gate20(.Q (g369), .QB (line20), .D(g11439), .CK(clk));
DFFX1 gate21(.Q (g1580), .QB (line21), .D(g7356), .CK(clk));
DFFX1 gate22(.Q (g1736), .QB (line22), .D(g6846), .CK(clk));
DFFX1 gate23(.Q (g39), .QB (line23), .D(g10774), .CK(clk));
DFFX1 gate24(.Q (g1651), .QB (line24), .D(g11182), .CK(clk));
DFFX1 gate25(.Q (g1424), .QB (line25), .D(g7330), .CK(clk));
DFFX1 gate26(.Q (g1737), .QB (line26), .D(g1736), .CK(clk));
DFFX1 gate27(.Q (g1672), .QB (line27), .D(g11037), .CK(clk));
DFFX1 gate28(.Q (g1077), .QB (line28), .D(g6805), .CK(clk));
DFFX1 gate29(.Q (g1231), .QB (line29), .D(g8279), .CK(clk));
DFFX1 gate30(.Q (g4), .QB (line30), .D(g8079), .CK(clk));
DFFX1 gate31(.Q (g774), .QB (line31), .D(g7785), .CK(clk));
DFFX1 gate32(.Q (g1104), .QB (line32), .D(g6815), .CK(clk));
DFFX1 gate33(.Q (g1304), .QB (line33), .D(g7290), .CK(clk));
DFFX1 gate34(.Q (g243), .QB (line34), .D(g7325), .CK(clk));
DFFX1 gate35(.Q (g1499), .QB (line35), .D(g8447), .CK(clk));
DFFX1 gate36(.Q (g1044), .QB (line36), .D(g7789), .CK(clk));
DFFX1 gate37(.Q (g1444), .QB (line37), .D(g8987), .CK(clk));
DFFX1 gate38(.Q (g757), .QB (line38), .D(g11179), .CK(clk));
DFFX1 gate39(.Q (g786), .QB (line39), .D(g8436), .CK(clk));
DFFX1 gate40(.Q (g1543), .QB (line40), .D(g7344), .CK(clk));
DFFX1 gate41(.Q (g552), .QB (line41), .D(g11045), .CK(clk));
DFFX1 gate42(.Q (g315), .QB (line42), .D(g5645), .CK(clk));
DFFX1 gate43(.Q (g1534), .QB (line43), .D(g7341), .CK(clk));
DFFX1 gate44(.Q (g622), .QB (line44), .D(g9338), .CK(clk));
DFFX1 gate45(.Q (g1927), .QB (line45), .D(g9354), .CK(clk));
DFFX1 gate46(.Q (g1660), .QB (line46), .D(g11033), .CK(clk));
DFFX1 gate47(.Q (g278), .QB (line47), .D(g7765), .CK(clk));
DFFX1 gate48(.Q (g1436), .QB (line48), .D(g8989), .CK(clk));
DFFX1 gate49(.Q (g718), .QB (line49), .D(g8433), .CK(clk));
DFFX1 gate50(.Q (g76), .QB (line50), .D(g7775), .CK(clk));
DFFX1 gate51(.Q (g554), .QB (line51), .D(g11047), .CK(clk));
DFFX1 gate52(.Q (g496), .QB (line52), .D(g11333), .CK(clk));
DFFX1 gate53(.Q (g981), .QB (line53), .D(g11472), .CK(clk));
DFFX1 gate54(.Q (g878), .QB (line54), .D(g4896), .CK(clk));
DFFX1 gate55(.Q (g590), .QB (line55), .D(g5653), .CK(clk));
DFFX1 gate56(.Q (g829), .QB (line56), .D(g4182), .CK(clk));
DFFX1 gate57(.Q (g1095), .QB (line57), .D(g6811), .CK(clk));
DFFX1 gate58(.Q (g704), .QB (line58), .D(g9344), .CK(clk));
DFFX1 gate59(.Q (g1265), .QB (line59), .D(g7302), .CK(clk));
DFFX1 gate60(.Q (g1786), .QB (line60), .D(g7814), .CK(clk));
DFFX1 gate61(.Q (g682), .QB (line61), .D(g8429), .CK(clk));
DFFX1 gate62(.Q (g1296), .QB (line62), .D(g7292), .CK(clk));
DFFX1 gate63(.Q (g587), .QB (line63), .D(g6295), .CK(clk));
DFFX1 gate64(.Q (g52), .QB (line64), .D(g7777), .CK(clk));
DFFX1 gate65(.Q (g646), .QB (line65), .D(g8065), .CK(clk));
DFFX1 gate66(.Q (g327), .QB (line66), .D(g5649), .CK(clk));
DFFX1 gate67(.Q (g1389), .QB (line67), .D(g6836), .CK(clk));
DFFX1 gate68(.Q (g1371), .QB (line68), .D(g7311), .CK(clk));
DFFX1 gate69(.Q (g1956), .QB (line69), .D(g1955), .CK(clk));
DFFX1 gate70(.Q (g1675), .QB (line70), .D(g11038), .CK(clk));
DFFX1 gate71(.Q (g354), .QB (line71), .D(g11508), .CK(clk));
DFFX1 gate72(.Q (g113), .QB (line72), .D(g7285), .CK(clk));
DFFX1 gate73(.Q (g639), .QB (line73), .D(g8063), .CK(clk));
DFFX1 gate74(.Q (g1684), .QB (line74), .D(g11041), .CK(clk));
DFFX1 gate75(.Q (g1639), .QB (line75), .D(g8448), .CK(clk));
DFFX1 gate76(.Q (g1791), .QB (line76), .D(g8080), .CK(clk));
DFFX1 gate77(.Q (g248), .QB (line77), .D(g7323), .CK(clk));
DFFX1 gate78(.Q (g1707), .QB (line78), .D(g4907), .CK(clk));
DFFX1 gate79(.Q (g1759), .QB (line79), .D(g5668), .CK(clk));
DFFX1 gate80(.Q (g351), .QB (line80), .D(g11507), .CK(clk));
DFFX1 gate81(.Q (g1957), .QB (line81), .D(g1956), .CK(clk));
DFFX1 gate82(.Q (g1604), .QB (line82), .D(g7364), .CK(clk));
DFFX1 gate83(.Q (g1098), .QB (line83), .D(g6812), .CK(clk));
DFFX1 gate84(.Q (g932), .QB (line84), .D(g8570), .CK(clk));
DFFX1 gate85(.Q (g126), .QB (line85), .D(g5642), .CK(clk));
DFFX1 gate86(.Q (g1896), .QB (line86), .D(g8282), .CK(clk));
DFFX1 gate87(.Q (g736), .QB (line87), .D(g8435), .CK(clk));
DFFX1 gate88(.Q (g1019), .QB (line88), .D(g7807), .CK(clk));
DFFX1 gate89(.Q (g1362), .QB (line89), .D(g7305), .CK(clk));
DFFX1 gate90(.Q (g745), .QB (line90), .D(g2639), .CK(clk));
DFFX1 gate91(.Q (g1419), .QB (line91), .D(g7332), .CK(clk));
DFFX1 gate92(.Q (g58), .QB (line92), .D(g7779), .CK(clk));
DFFX1 gate93(.Q (g32), .QB (line93), .D(g11397), .CK(clk));
DFFX1 gate94(.Q (g876), .QB (line94), .D(g878), .CK(clk));
DFFX1 gate95(.Q (g1086), .QB (line95), .D(g6808), .CK(clk));
DFFX1 gate96(.Q (g1486), .QB (line96), .D(g8444), .CK(clk));
DFFX1 gate97(.Q (g1730), .QB (line97), .D(g10881), .CK(clk));
DFFX1 gate98(.Q (g1504), .QB (line98), .D(g7328), .CK(clk));
DFFX1 gate99(.Q (g1470), .QB (line99), .D(g8440), .CK(clk));
DFFX1 gate100(.Q (g822), .QB (line100), .D(g8437), .CK(clk));
DFFX1 gate101(.Q (g583), .QB (line101), .D(g6291), .CK(clk));
DFFX1 gate102(.Q (g1678), .QB (line102), .D(g11039), .CK(clk));
DFFX1 gate103(.Q (g174), .QB (line103), .D(g8423), .CK(clk));
DFFX1 gate104(.Q (g1766), .QB (line104), .D(g7810), .CK(clk));
DFFX1 gate105(.Q (g1801), .QB (line105), .D(g8450), .CK(clk));
DFFX1 gate106(.Q (g186), .QB (line106), .D(g7317), .CK(clk));
DFFX1 gate107(.Q (g959), .QB (line107), .D(g11403), .CK(clk));
DFFX1 gate108(.Q (g1169), .QB (line108), .D(g6314), .CK(clk));
DFFX1 gate109(.Q (g1007), .QB (line109), .D(g7806), .CK(clk));
DFFX1 gate110(.Q (g1407), .QB (line110), .D(g8993), .CK(clk));
DFFX1 gate111(.Q (g1059), .QB (line111), .D(g7794), .CK(clk));
DFFX1 gate112(.Q (g1868), .QB (line112), .D(g7817), .CK(clk));
DFFX1 gate113(.Q (g758), .QB (line113), .D(g6797), .CK(clk));
DFFX1 gate114(.Q (g1718), .QB (line114), .D(g6337), .CK(clk));
DFFX1 gate115(.Q (g396), .QB (line115), .D(g11265), .CK(clk));
DFFX1 gate116(.Q (g1015), .QB (line116), .D(g7808), .CK(clk));
DFFX1 gate117(.Q (g38), .QB (line117), .D(g10872), .CK(clk));
DFFX1 gate118(.Q (g632), .QB (line118), .D(g5655), .CK(clk));
DFFX1 gate119(.Q (g1415), .QB (line119), .D(g7335), .CK(clk));
DFFX1 gate120(.Q (g1227), .QB (line120), .D(g8278), .CK(clk));
DFFX1 gate121(.Q (g1721), .QB (line121), .D(g10878), .CK(clk));
DFFX1 gate122(.Q (g882), .QB (line122), .D(g883), .CK(clk));
DFFX1 gate123(.Q (g16), .QB (line123), .D(g4906), .CK(clk));
DFFX1 gate124(.Q (g284), .QB (line124), .D(g7767), .CK(clk));
DFFX1 gate125(.Q (g426), .QB (line125), .D(g11256), .CK(clk));
DFFX1 gate126(.Q (g219), .QB (line126), .D(g7310), .CK(clk));
DFFX1 gate127(.Q (g1216), .QB (line127), .D(g1360), .CK(clk));
DFFX1 gate128(.Q (g806), .QB (line128), .D(g7289), .CK(clk));
DFFX1 gate129(.Q (g1428), .QB (line129), .D(g8992), .CK(clk));
DFFX1 gate130(.Q (g579), .QB (line130), .D(g6287), .CK(clk));
DFFX1 gate131(.Q (g1564), .QB (line131), .D(g7351), .CK(clk));
DFFX1 gate132(.Q (g1741), .QB (line132), .D(g5662), .CK(clk));
DFFX1 gate133(.Q (g225), .QB (line133), .D(g7309), .CK(clk));
DFFX1 gate134(.Q (g281), .QB (line134), .D(g7766), .CK(clk));
DFFX1 gate135(.Q (g1308), .QB (line135), .D(g11627), .CK(clk));
DFFX1 gate136(.Q (g611), .QB (line136), .D(g9930), .CK(clk));
DFFX1 gate137(.Q (g631), .QB (line137), .D(g5654), .CK(clk));
DFFX1 gate138(.Q (g1217), .QB (line138), .D(g9823), .CK(clk));
DFFX1 gate139(.Q (g1589), .QB (line139), .D(g7359), .CK(clk));
DFFX1 gate140(.Q (g1466), .QB (line140), .D(g8439), .CK(clk));
DFFX1 gate141(.Q (g1571), .QB (line141), .D(g7353), .CK(clk));
DFFX1 gate142(.Q (g1861), .QB (line142), .D(g7815), .CK(clk));
DFFX1 gate143(.Q (g1365), .QB (line143), .D(g7307), .CK(clk));
DFFX1 gate144(.Q (g1448), .QB (line144), .D(g11594), .CK(clk));
DFFX1 gate145(.Q (g1711), .QB (line145), .D(g6335), .CK(clk));
DFFX1 gate146(.Q (g1133), .QB (line146), .D(g6309), .CK(clk));
DFFX1 gate147(.Q (g1333), .QB (line147), .D(g11635), .CK(clk));
DFFX1 gate148(.Q (g153), .QB (line148), .D(g8426), .CK(clk));
DFFX1 gate149(.Q (g962), .QB (line149), .D(g11404), .CK(clk));
DFFX1 gate150(.Q (g766), .QB (line150), .D(g6799), .CK(clk));
DFFX1 gate151(.Q (g588), .QB (line151), .D(g6296), .CK(clk));
DFFX1 gate152(.Q (g486), .QB (line152), .D(g11331), .CK(clk));
DFFX1 gate153(.Q (g471), .QB (line153), .D(g11469), .CK(clk));
DFFX1 gate154(.Q (g1397), .QB (line154), .D(g7322), .CK(clk));
DFFX1 gate155(.Q (g580), .QB (line155), .D(g6288), .CK(clk));
DFFX1 gate156(.Q (g1950), .QB (line156), .D(g8288), .CK(clk));
DFFX1 gate157(.Q (g756), .QB (line157), .D(g755), .CK(clk));
DFFX1 gate158(.Q (g635), .QB (line158), .D(g5656), .CK(clk));
DFFX1 gate159(.Q (g1101), .QB (line159), .D(g6814), .CK(clk));
DFFX1 gate160(.Q (g549), .QB (line160), .D(g11044), .CK(clk));
DFFX1 gate161(.Q (g1041), .QB (line161), .D(g7788), .CK(clk));
DFFX1 gate162(.Q (g105), .QB (line162), .D(g11180), .CK(clk));
DFFX1 gate163(.Q (g1669), .QB (line163), .D(g11036), .CK(clk));
DFFX1 gate164(.Q (g1368), .QB (line164), .D(g7308), .CK(clk));
DFFX1 gate165(.Q (g1531), .QB (line165), .D(g7340), .CK(clk));
DFFX1 gate166(.Q (g1458), .QB (line166), .D(g7327), .CK(clk));
DFFX1 gate167(.Q (g572), .QB (line167), .D(g10877), .CK(clk));
DFFX1 gate168(.Q (g1011), .QB (line168), .D(g7805), .CK(clk));
DFFX1 gate169(.Q (g33), .QB (line169), .D(g10867), .CK(clk));
DFFX1 gate170(.Q (g1411), .QB (line170), .D(g7331), .CK(clk));
DFFX1 gate171(.Q (g1074), .QB (line171), .D(g6813), .CK(clk));
DFFX1 gate172(.Q (g444), .QB (line172), .D(g11259), .CK(clk));
DFFX1 gate173(.Q (g1474), .QB (line173), .D(g8441), .CK(clk));
DFFX1 gate174(.Q (g1080), .QB (line174), .D(g6806), .CK(clk));
DFFX1 gate175(.Q (g1713), .QB (line175), .D(g6336), .CK(clk));
DFFX1 gate176(.Q (g333), .QB (line176), .D(g5651), .CK(clk));
DFFX1 gate177(.Q (g269), .QB (line177), .D(g7762), .CK(clk));
DFFX1 gate178(.Q (g401), .QB (line178), .D(g11266), .CK(clk));
DFFX1 gate179(.Q (g1857), .QB (line179), .D(g11409), .CK(clk));
DFFX1 gate180(.Q (g9), .QB (line180), .D(g7336), .CK(clk));
DFFX1 gate181(.Q (g664), .QB (line181), .D(g8782), .CK(clk));
DFFX1 gate182(.Q (g965), .QB (line182), .D(g11405), .CK(clk));
DFFX1 gate183(.Q (g1400), .QB (line183), .D(g7324), .CK(clk));
DFFX1 gate184(.Q (g309), .QB (line184), .D(g5652), .CK(clk));
DFFX1 gate185(.Q (g814), .QB (line185), .D(g8077), .CK(clk));
DFFX1 gate186(.Q (g231), .QB (line186), .D(g7319), .CK(clk));
DFFX1 gate187(.Q (g557), .QB (line187), .D(g11048), .CK(clk));
DFFX1 gate188(.Q (g586), .QB (line188), .D(g6294), .CK(clk));
DFFX1 gate189(.Q (g869), .QB (line189), .D(g875), .CK(clk));
DFFX1 gate190(.Q (g1383), .QB (line190), .D(g7316), .CK(clk));
DFFX1 gate191(.Q (g158), .QB (line191), .D(g8425), .CK(clk));
DFFX1 gate192(.Q (g627), .QB (line192), .D(g5657), .CK(clk));
DFFX1 gate193(.Q (g1023), .QB (line193), .D(g7799), .CK(clk));
DFFX1 gate194(.Q (g259), .QB (line194), .D(g7755), .CK(clk));
DFFX1 gate195(.Q (g1361), .QB (line195), .D(g1206), .CK(clk));
DFFX1 gate196(.Q (g1327), .QB (line196), .D(g11633), .CK(clk));
DFFX1 gate197(.Q (g654), .QB (line197), .D(g8067), .CK(clk));
DFFX1 gate198(.Q (g293), .QB (line198), .D(g7770), .CK(clk));
DFFX1 gate199(.Q (g1346), .QB (line199), .D(g11656), .CK(clk));
DFFX1 gate200(.Q (g1633), .QB (line200), .D(g8873), .CK(clk));
DFFX1 gate201(.Q (g1753), .QB (line201), .D(g5666), .CK(clk));
DFFX1 gate202(.Q (g1508), .QB (line202), .D(g7329), .CK(clk));
DFFX1 gate203(.Q (g1240), .QB (line203), .D(g7297), .CK(clk));
DFFX1 gate204(.Q (g538), .QB (line204), .D(g11326), .CK(clk));
DFFX1 gate205(.Q (g416), .QB (line205), .D(g11269), .CK(clk));
DFFX1 gate206(.Q (g542), .QB (line206), .D(g11325), .CK(clk));
DFFX1 gate207(.Q (g1681), .QB (line207), .D(g11040), .CK(clk));
DFFX1 gate208(.Q (g374), .QB (line208), .D(g11440), .CK(clk));
DFFX1 gate209(.Q (g563), .QB (line209), .D(g11050), .CK(clk));
DFFX1 gate210(.Q (g1914), .QB (line210), .D(g8284), .CK(clk));
DFFX1 gate211(.Q (g530), .QB (line211), .D(g11328), .CK(clk));
DFFX1 gate212(.Q (g575), .QB (line212), .D(g11052), .CK(clk));
DFFX1 gate213(.Q (g1936), .QB (line213), .D(g9355), .CK(clk));
DFFX1 gate214(.Q (g55), .QB (line214), .D(g7778), .CK(clk));
DFFX1 gate215(.Q (g1117), .QB (line215), .D(g6299), .CK(clk));
DFFX1 gate216(.Q (g1317), .QB (line216), .D(g1356), .CK(clk));
DFFX1 gate217(.Q (g357), .QB (line217), .D(g11509), .CK(clk));
DFFX1 gate218(.Q (g386), .QB (line218), .D(g11263), .CK(clk));
DFFX1 gate219(.Q (g1601), .QB (line219), .D(g7363), .CK(clk));
DFFX1 gate220(.Q (g553), .QB (line220), .D(g11046), .CK(clk));
DFFX1 gate221(.Q (g166), .QB (line221), .D(g7747), .CK(clk));
DFFX1 gate222(.Q (g501), .QB (line222), .D(g11334), .CK(clk));
DFFX1 gate223(.Q (g262), .QB (line223), .D(g7758), .CK(clk));
DFFX1 gate224(.Q (g1840), .QB (line224), .D(g8694), .CK(clk));
DFFX1 gate225(.Q (g70), .QB (line225), .D(g7783), .CK(clk));
DFFX1 gate226(.Q (g318), .QB (line226), .D(g5646), .CK(clk));
DFFX1 gate227(.Q (g1356), .QB (line227), .D(g6818), .CK(clk));
DFFX1 gate228(.Q (g794), .QB (line228), .D(g6800), .CK(clk));
DFFX1 gate229(.Q (g36), .QB (line229), .D(g10870), .CK(clk));
DFFX1 gate230(.Q (g302), .QB (line230), .D(g7773), .CK(clk));
DFFX1 gate231(.Q (g342), .QB (line231), .D(g11513), .CK(clk));
DFFX1 gate232(.Q (g1250), .QB (line232), .D(g7299), .CK(clk));
DFFX1 gate233(.Q (g1163), .QB (line233), .D(g6301), .CK(clk));
DFFX1 gate234(.Q (g1810), .QB (line234), .D(g2044), .CK(clk));
DFFX1 gate235(.Q (g1032), .QB (line235), .D(g7800), .CK(clk));
DFFX1 gate236(.Q (g1432), .QB (line236), .D(g8990), .CK(clk));
DFFX1 gate237(.Q (g1053), .QB (line237), .D(g7792), .CK(clk));
DFFX1 gate238(.Q (g1453), .QB (line238), .D(g7326), .CK(clk));
DFFX1 gate239(.Q (g363), .QB (line239), .D(g11511), .CK(clk));
DFFX1 gate240(.Q (g330), .QB (line240), .D(g5650), .CK(clk));
DFFX1 gate241(.Q (g1157), .QB (line241), .D(g6303), .CK(clk));
DFFX1 gate242(.Q (g1357), .QB (line242), .D(g6330), .CK(clk));
DFFX1 gate243(.Q (g35), .QB (line243), .D(g10869), .CK(clk));
DFFX1 gate244(.Q (g928), .QB (line244), .D(g8569), .CK(clk));
DFFX1 gate245(.Q (g261), .QB (line245), .D(g7757), .CK(clk));
DFFX1 gate246(.Q (g516), .QB (line246), .D(g11337), .CK(clk));
DFFX1 gate247(.Q (g254), .QB (line247), .D(g7759), .CK(clk));
DFFX1 gate248(.Q (g778), .QB (line248), .D(g8076), .CK(clk));
DFFX1 gate249(.Q (g861), .QB (line249), .D(g4190), .CK(clk));
DFFX1 gate250(.Q (g1627), .QB (line250), .D(g8871), .CK(clk));
DFFX1 gate251(.Q (g1292), .QB (line251), .D(g7293), .CK(clk));
DFFX1 gate252(.Q (g290), .QB (line252), .D(g7769), .CK(clk));
DFFX1 gate253(.Q (g1850), .QB (line253), .D(g5671), .CK(clk));
DFFX1 gate254(.Q (g770), .QB (line254), .D(g7288), .CK(clk));
DFFX1 gate255(.Q (g1583), .QB (line255), .D(g7357), .CK(clk));
DFFX1 gate256(.Q (g466), .QB (line256), .D(g11468), .CK(clk));
DFFX1 gate257(.Q (g1561), .QB (line257), .D(g7350), .CK(clk));
DFFX1 gate258(.Q (g1527), .QB (line258), .D(g4899), .CK(clk));
DFFX1 gate259(.Q (g1546), .QB (line259), .D(g7345), .CK(clk));
DFFX1 gate260(.Q (g287), .QB (line260), .D(g7768), .CK(clk));
DFFX1 gate261(.Q (g560), .QB (line261), .D(g11049), .CK(clk));
DFFX1 gate262(.Q (g617), .QB (line262), .D(g8780), .CK(clk));
DFFX1 gate263(.Q (g17), .QB (line263), .D(g4894), .CK(clk));
DFFX1 gate264(.Q (g336), .QB (line264), .D(g11653), .CK(clk));
DFFX1 gate265(.Q (g456), .QB (line265), .D(g11466), .CK(clk));
DFFX1 gate266(.Q (g305), .QB (line266), .D(g5643), .CK(clk));
DFFX1 gate267(.Q (g345), .QB (line267), .D(g11642), .CK(clk));
DFFX1 gate268(.Q (g8), .QB (line268), .D(g2613), .CK(clk));
DFFX1 gate269(.Q (g1771), .QB (line269), .D(g7811), .CK(clk));
DFFX1 gate270(.Q (g865), .QB (line270), .D(g8275), .CK(clk));
DFFX1 gate271(.Q (g255), .QB (line271), .D(g7751), .CK(clk));
DFFX1 gate272(.Q (g1945), .QB (line272), .D(g9356), .CK(clk));
DFFX1 gate273(.Q (g1738), .QB (line273), .D(g5661), .CK(clk));
DFFX1 gate274(.Q (g1478), .QB (line274), .D(g8442), .CK(clk));
DFFX1 gate275(.Q (g1035), .QB (line275), .D(g7787), .CK(clk));
DFFX1 gate276(.Q (g1959), .QB (line276), .D(g4217), .CK(clk));
DFFX1 gate277(.Q (g1690), .QB (line277), .D(g6844), .CK(clk));
DFFX1 gate278(.Q (g1482), .QB (line278), .D(g8443), .CK(clk));
DFFX1 gate279(.Q (g1110), .QB (line279), .D(g6817), .CK(clk));
DFFX1 gate280(.Q (g296), .QB (line280), .D(g7771), .CK(clk));
DFFX1 gate281(.Q (g1663), .QB (line281), .D(g11034), .CK(clk));
DFFX1 gate282(.Q (g700), .QB (line282), .D(g8431), .CK(clk));
DFFX1 gate283(.Q (g1762), .QB (line283), .D(g5669), .CK(clk));
DFFX1 gate284(.Q (g360), .QB (line284), .D(g11510), .CK(clk));
DFFX1 gate285(.Q (g192), .QB (line285), .D(g6837), .CK(clk));
DFFX1 gate286(.Q (g1657), .QB (line286), .D(g10875), .CK(clk));
DFFX1 gate287(.Q (g722), .QB (line287), .D(g9346), .CK(clk));
DFFX1 gate288(.Q (g61), .QB (line288), .D(g7780), .CK(clk));
DFFX1 gate289(.Q (g566), .QB (line289), .D(g11051), .CK(clk));
DFFX1 gate290(.Q (g1394), .QB (line290), .D(g7809), .CK(clk));
DFFX1 gate291(.Q (g1089), .QB (line291), .D(g6809), .CK(clk));
DFFX1 gate292(.Q (g883), .QB (line292), .D(g4897), .CK(clk));
DFFX1 gate293(.Q (g1071), .QB (line293), .D(g6804), .CK(clk));
DFFX1 gate294(.Q (g986), .QB (line294), .D(g11473), .CK(clk));
DFFX1 gate295(.Q (g971), .QB (line295), .D(g11470), .CK(clk));
DFFX1 gate296(.Q (g1955), .QB (line296), .D(g6338), .CK(clk));
DFFX1 gate297(.Q (g143), .QB (line297), .D(g7746), .CK(clk));
DFFX1 gate298(.Q (g1814), .QB (line298), .D(g9825), .CK(clk));
DFFX1 gate299(.Q (g1038), .QB (line299), .D(g7797), .CK(clk));
DFFX1 gate300(.Q (g1212), .QB (line300), .D(g1217), .CK(clk));
DFFX1 gate301(.Q (g1918), .QB (line301), .D(g9353), .CK(clk));
DFFX1 gate302(.Q (g782), .QB (line302), .D(g8273), .CK(clk));
DFFX1 gate303(.Q (g1822), .QB (line303), .D(g9826), .CK(clk));
DFFX1 gate304(.Q (g237), .QB (line304), .D(g7306), .CK(clk));
DFFX1 gate305(.Q (g746), .QB (line305), .D(g2638), .CK(clk));
DFFX1 gate306(.Q (g1062), .QB (line306), .D(g7795), .CK(clk));
DFFX1 gate307(.Q (g1462), .QB (line307), .D(g8438), .CK(clk));
DFFX1 gate308(.Q (g178), .QB (line308), .D(g7748), .CK(clk));
DFFX1 gate309(.Q (g366), .QB (line309), .D(g11512), .CK(clk));
DFFX1 gate310(.Q (g837), .QB (line310), .D(g4184), .CK(clk));
DFFX1 gate311(.Q (g599), .QB (line311), .D(g9819), .CK(clk));
DFFX1 gate312(.Q (g1854), .QB (line312), .D(g11408), .CK(clk));
DFFX1 gate313(.Q (g944), .QB (line313), .D(g11398), .CK(clk));
DFFX1 gate314(.Q (g1941), .QB (line314), .D(g8287), .CK(clk));
DFFX1 gate315(.Q (g170), .QB (line315), .D(g8422), .CK(clk));
DFFX1 gate316(.Q (g1520), .QB (line316), .D(g7334), .CK(clk));
DFFX1 gate317(.Q (g686), .QB (line317), .D(g9342), .CK(clk));
DFFX1 gate318(.Q (g953), .QB (line318), .D(g11401), .CK(clk));
DFFX1 gate319(.Q (g1958), .QB (line319), .D(g6339), .CK(clk));
DFFX1 gate320(.Q (g40), .QB (line320), .D(g10775), .CK(clk));
DFFX1 gate321(.Q (g1765), .QB (line321), .D(g3329), .CK(clk));
DFFX1 gate322(.Q (g1733), .QB (line322), .D(g10882), .CK(clk));
DFFX1 gate323(.Q (g1270), .QB (line323), .D(g7303), .CK(clk));
DFFX1 gate324(.Q (g1610), .QB (line324), .D(g6845), .CK(clk));
DFFX1 gate325(.Q (g1796), .QB (line325), .D(g8280), .CK(clk));
DFFX1 gate326(.Q (g1324), .QB (line326), .D(g11632), .CK(clk));
DFFX1 gate327(.Q (g1540), .QB (line327), .D(g7343), .CK(clk));
DFFX1 gate328(.Q (g1377), .QB (line328), .D(g7312), .CK(clk));
DFFX1 gate329(.Q (g1206), .QB (line329), .D(g4898), .CK(clk));
DFFX1 gate330(.Q (g491), .QB (line330), .D(g11332), .CK(clk));
DFFX1 gate331(.Q (g1849), .QB (line331), .D(g5670), .CK(clk));
DFFX1 gate332(.Q (g213), .QB (line332), .D(g7313), .CK(clk));
DFFX1 gate333(.Q (g1781), .QB (line333), .D(g7813), .CK(clk));
DFFX1 gate334(.Q (g1900), .QB (line334), .D(g9351), .CK(clk));
DFFX1 gate335(.Q (g1245), .QB (line335), .D(g7298), .CK(clk));
DFFX1 gate336(.Q (g108), .QB (line336), .D(g11593), .CK(clk));
DFFX1 gate337(.Q (g630), .QB (line337), .D(g7287), .CK(clk));
DFFX1 gate338(.Q (g148), .QB (line338), .D(g8427), .CK(clk));
DFFX1 gate339(.Q (g833), .QB (line339), .D(g4183), .CK(clk));
DFFX1 gate340(.Q (g1923), .QB (line340), .D(g8285), .CK(clk));
DFFX1 gate341(.Q (g936), .QB (line341), .D(g8571), .CK(clk));
DFFX1 gate342(.Q (g1215), .QB (line342), .D(g6315), .CK(clk));
DFFX1 gate343(.Q (g1314), .QB (line343), .D(g11629), .CK(clk));
DFFX1 gate344(.Q (g849), .QB (line344), .D(g4187), .CK(clk));
DFFX1 gate345(.Q (g1336), .QB (line345), .D(g11654), .CK(clk));
DFFX1 gate346(.Q (g272), .QB (line346), .D(g7763), .CK(clk));
DFFX1 gate347(.Q (g1806), .QB (line347), .D(g8573), .CK(clk));
DFFX1 gate348(.Q (g826), .QB (line348), .D(g8568), .CK(clk));
DFFX1 gate349(.Q (g1065), .QB (line349), .D(g7796), .CK(clk));
DFFX1 gate350(.Q (g1887), .QB (line350), .D(g8281), .CK(clk));
DFFX1 gate351(.Q (g37), .QB (line351), .D(g10871), .CK(clk));
DFFX1 gate352(.Q (g968), .QB (line352), .D(g11406), .CK(clk));
DFFX1 gate353(.Q (g1845), .QB (line353), .D(g5673), .CK(clk));
DFFX1 gate354(.Q (g1137), .QB (line354), .D(g6310), .CK(clk));
DFFX1 gate355(.Q (g1891), .QB (line355), .D(g9350), .CK(clk));
DFFX1 gate356(.Q (g1255), .QB (line356), .D(g7300), .CK(clk));
DFFX1 gate357(.Q (g257), .QB (line357), .D(g7753), .CK(clk));
DFFX1 gate358(.Q (g874), .QB (line358), .D(g9821), .CK(clk));
DFFX1 gate359(.Q (g591), .QB (line359), .D(g9818), .CK(clk));
DFFX1 gate360(.Q (g731), .QB (line360), .D(g9347), .CK(clk));
DFFX1 gate361(.Q (g636), .QB (line361), .D(g8781), .CK(clk));
DFFX1 gate362(.Q (g1218), .QB (line362), .D(g8276), .CK(clk));
DFFX1 gate363(.Q (g605), .QB (line363), .D(g9820), .CK(clk));
DFFX1 gate364(.Q (g79), .QB (line364), .D(g7776), .CK(clk));
DFFX1 gate365(.Q (g182), .QB (line365), .D(g7749), .CK(clk));
DFFX1 gate366(.Q (g950), .QB (line366), .D(g11400), .CK(clk));
DFFX1 gate367(.Q (g1129), .QB (line367), .D(g6308), .CK(clk));
DFFX1 gate368(.Q (g857), .QB (line368), .D(g4189), .CK(clk));
DFFX1 gate369(.Q (g448), .QB (line369), .D(g11258), .CK(clk));
DFFX1 gate370(.Q (g1828), .QB (line370), .D(g9827), .CK(clk));
DFFX1 gate371(.Q (g1727), .QB (line371), .D(g10880), .CK(clk));
DFFX1 gate372(.Q (g1592), .QB (line372), .D(g7360), .CK(clk));
DFFX1 gate373(.Q (g1703), .QB (line373), .D(g6843), .CK(clk));
DFFX1 gate374(.Q (g1932), .QB (line374), .D(g8286), .CK(clk));
DFFX1 gate375(.Q (g1624), .QB (line375), .D(g8870), .CK(clk));
DFFX1 gate376(.Q (g26), .QB (line376), .D(g4885), .CK(clk));
DFFX1 gate377(.Q (g1068), .QB (line377), .D(g6803), .CK(clk));
DFFX1 gate378(.Q (g578), .QB (line378), .D(g6286), .CK(clk));
DFFX1 gate379(.Q (g440), .QB (line379), .D(g11260), .CK(clk));
DFFX1 gate380(.Q (g476), .QB (line380), .D(g11338), .CK(clk));
DFFX1 gate381(.Q (g119), .QB (line381), .D(g7745), .CK(clk));
DFFX1 gate382(.Q (g668), .QB (line382), .D(g9340), .CK(clk));
DFFX1 gate383(.Q (g139), .QB (line383), .D(g8418), .CK(clk));
DFFX1 gate384(.Q (g1149), .QB (line384), .D(g6305), .CK(clk));
DFFX1 gate385(.Q (g34), .QB (line385), .D(g10868), .CK(clk));
DFFX1 gate386(.Q (g1848), .QB (line386), .D(g7366), .CK(clk));
DFFX1 gate387(.Q (g263), .QB (line387), .D(g7760), .CK(clk));
DFFX1 gate388(.Q (g818), .QB (line388), .D(g8274), .CK(clk));
DFFX1 gate389(.Q (g1747), .QB (line389), .D(g5664), .CK(clk));
DFFX1 gate390(.Q (g802), .QB (line390), .D(g6802), .CK(clk));
DFFX1 gate391(.Q (g275), .QB (line391), .D(g7764), .CK(clk));
DFFX1 gate392(.Q (g1524), .QB (line392), .D(g7338), .CK(clk));
DFFX1 gate393(.Q (g1577), .QB (line393), .D(g7355), .CK(clk));
DFFX1 gate394(.Q (g810), .QB (line394), .D(g7786), .CK(clk));
DFFX1 gate395(.Q (g391), .QB (line395), .D(g11264), .CK(clk));
DFFX1 gate396(.Q (g658), .QB (line396), .D(g9339), .CK(clk));
DFFX1 gate397(.Q (g1386), .QB (line397), .D(g7318), .CK(clk));
DFFX1 gate398(.Q (g253), .QB (line398), .D(g7750), .CK(clk));
DFFX1 gate399(.Q (g875), .QB (line399), .D(g9822), .CK(clk));
DFFX1 gate400(.Q (g1125), .QB (line400), .D(g6307), .CK(clk));
DFFX1 gate401(.Q (g201), .QB (line401), .D(g7304), .CK(clk));
DFFX1 gate402(.Q (g1280), .QB (line402), .D(g7295), .CK(clk));
DFFX1 gate403(.Q (g1083), .QB (line403), .D(g6807), .CK(clk));
DFFX1 gate404(.Q (g650), .QB (line404), .D(g8066), .CK(clk));
DFFX1 gate405(.Q (g1636), .QB (line405), .D(g8874), .CK(clk));
DFFX1 gate406(.Q (g853), .QB (line406), .D(g4188), .CK(clk));
DFFX1 gate407(.Q (g421), .QB (line407), .D(g11270), .CK(clk));
DFFX1 gate408(.Q (g762), .QB (line408), .D(g6798), .CK(clk));
DFFX1 gate409(.Q (g956), .QB (line409), .D(g11402), .CK(clk));
DFFX1 gate410(.Q (g378), .QB (line410), .D(g11441), .CK(clk));
DFFX1 gate411(.Q (g1756), .QB (line411), .D(g5667), .CK(clk));
DFFX1 gate412(.Q (g589), .QB (line412), .D(g6297), .CK(clk));
DFFX1 gate413(.Q (g841), .QB (line413), .D(g4185), .CK(clk));
DFFX1 gate414(.Q (g1027), .QB (line414), .D(g7798), .CK(clk));
DFFX1 gate415(.Q (g1003), .QB (line415), .D(g7803), .CK(clk));
DFFX1 gate416(.Q (g1403), .QB (line416), .D(g8991), .CK(clk));
DFFX1 gate417(.Q (g1145), .QB (line417), .D(g6312), .CK(clk));
DFFX1 gate418(.Q (g1107), .QB (line418), .D(g6816), .CK(clk));
DFFX1 gate419(.Q (g1223), .QB (line419), .D(g8277), .CK(clk));
DFFX1 gate420(.Q (g406), .QB (line420), .D(g11267), .CK(clk));
DFFX1 gate421(.Q (g1811), .QB (line421), .D(g11185), .CK(clk));
DFFX1 gate422(.Q (g1642), .QB (line422), .D(g11183), .CK(clk));
DFFX1 gate423(.Q (g1047), .QB (line423), .D(g7790), .CK(clk));
DFFX1 gate424(.Q (g1654), .QB (line424), .D(g10874), .CK(clk));
DFFX1 gate425(.Q (g197), .QB (line425), .D(g6835), .CK(clk));
DFFX1 gate426(.Q (g1595), .QB (line426), .D(g7361), .CK(clk));
DFFX1 gate427(.Q (g1537), .QB (line427), .D(g7342), .CK(clk));
DFFX1 gate428(.Q (g727), .QB (line428), .D(g8434), .CK(clk));
DFFX1 gate429(.Q (g999), .QB (line429), .D(g7804), .CK(clk));
DFFX1 gate430(.Q (g798), .QB (line430), .D(g6801), .CK(clk));
DFFX1 gate431(.Q (g481), .QB (line431), .D(g11324), .CK(clk));
DFFX1 gate432(.Q (g754), .QB (line432), .D(g4895), .CK(clk));
DFFX1 gate433(.Q (g1330), .QB (line433), .D(g11634), .CK(clk));
DFFX1 gate434(.Q (g845), .QB (line434), .D(g4186), .CK(clk));
DFFX1 gate435(.Q (g790), .QB (line435), .D(g8567), .CK(clk));
DFFX1 gate436(.Q (g1512), .QB (line436), .D(g8449), .CK(clk));
DFFX1 gate437(.Q (g114), .QB (line437), .D(g113), .CK(clk));
DFFX1 gate438(.Q (g1490), .QB (line438), .D(g8445), .CK(clk));
DFFX1 gate439(.Q (g1166), .QB (line439), .D(g6300), .CK(clk));
DFFX1 gate440(.Q (g1056), .QB (line440), .D(g7793), .CK(clk));
DFFX1 gate441(.Q (g348), .QB (line441), .D(g11506), .CK(clk));
DFFX1 gate442(.Q (g868), .QB (line442), .D(g874), .CK(clk));
DFFX1 gate443(.Q (g1260), .QB (line443), .D(g7301), .CK(clk));
DFFX1 gate444(.Q (g260), .QB (line444), .D(g7756), .CK(clk));
DFFX1 gate445(.Q (g131), .QB (line445), .D(g8420), .CK(clk));
DFFX1 gate446(.Q (g7), .QB (line446), .D(g2731), .CK(clk));
DFFX1 gate447(.Q (g258), .QB (line447), .D(g7754), .CK(clk));
DFFX1 gate448(.Q (g521), .QB (line448), .D(g11330), .CK(clk));
DFFX1 gate449(.Q (g1318), .QB (line449), .D(g11630), .CK(clk));
DFFX1 gate450(.Q (g1872), .QB (line450), .D(g9348), .CK(clk));
DFFX1 gate451(.Q (g677), .QB (line451), .D(g9341), .CK(clk));
DFFX1 gate452(.Q (g582), .QB (line452), .D(g6290), .CK(clk));
DFFX1 gate453(.Q (g1393), .QB (line453), .D(g7320), .CK(clk));
DFFX1 gate454(.Q (g1549), .QB (line454), .D(g7346), .CK(clk));
DFFX1 gate455(.Q (g947), .QB (line455), .D(g11399), .CK(clk));
DFFX1 gate456(.Q (g1834), .QB (line456), .D(g9895), .CK(clk));
DFFX1 gate457(.Q (g1598), .QB (line457), .D(g7362), .CK(clk));
DFFX1 gate458(.Q (g1121), .QB (line458), .D(g6306), .CK(clk));
DFFX1 gate459(.Q (g1321), .QB (line459), .D(g11631), .CK(clk));
DFFX1 gate460(.Q (g506), .QB (line460), .D(g11335), .CK(clk));
DFFX1 gate461(.Q (g546), .QB (line461), .D(g11043), .CK(clk));
DFFX1 gate462(.Q (g1909), .QB (line462), .D(g9352), .CK(clk));
DFFX1 gate463(.Q (g755), .QB (line463), .D(g6298), .CK(clk));
DFFX1 gate464(.Q (g1552), .QB (line464), .D(g7347), .CK(clk));
DFFX1 gate465(.Q (g584), .QB (line465), .D(g6292), .CK(clk));
DFFX1 gate466(.Q (g1687), .QB (line466), .D(g11042), .CK(clk));
DFFX1 gate467(.Q (g1586), .QB (line467), .D(g7358), .CK(clk));
DFFX1 gate468(.Q (g324), .QB (line468), .D(g5648), .CK(clk));
DFFX1 gate469(.Q (g1141), .QB (line469), .D(g6311), .CK(clk));
DFFX1 gate470(.Q (g1570), .QB (line470), .D(g4900), .CK(clk));
DFFX1 gate471(.Q (g1341), .QB (line471), .D(g11655), .CK(clk));
DFFX1 gate472(.Q (g1710), .QB (line472), .D(g4901), .CK(clk));
DFFX1 gate473(.Q (g1645), .QB (line473), .D(g11184), .CK(clk));
DFFX1 gate474(.Q (g115), .QB (line474), .D(g7321), .CK(clk));
DFFX1 gate475(.Q (g135), .QB (line475), .D(g8419), .CK(clk));
DFFX1 gate476(.Q (g525), .QB (line476), .D(g11329), .CK(clk));
DFFX1 gate477(.Q (g581), .QB (line477), .D(g6289), .CK(clk));
DFFX1 gate478(.Q (g1607), .QB (line478), .D(g7365), .CK(clk));
DFFX1 gate479(.Q (g321), .QB (line479), .D(g5647), .CK(clk));
DFFX1 gate480(.Q (g67), .QB (line480), .D(g7782), .CK(clk));
DFFX1 gate481(.Q (g1275), .QB (line481), .D(g11443), .CK(clk));
DFFX1 gate482(.Q (g1311), .QB (line482), .D(g11628), .CK(clk));
DFFX1 gate483(.Q (g1615), .QB (line483), .D(g8868), .CK(clk));
DFFX1 gate484(.Q (g382), .QB (line484), .D(g11442), .CK(clk));
DFFX1 gate485(.Q (g1374), .QB (line485), .D(g6825), .CK(clk));
DFFX1 gate486(.Q (g266), .QB (line486), .D(g7761), .CK(clk));
DFFX1 gate487(.Q (g1284), .QB (line487), .D(g7294), .CK(clk));
DFFX1 gate488(.Q (g1380), .QB (line488), .D(g7314), .CK(clk));
DFFX1 gate489(.Q (g673), .QB (line489), .D(g8428), .CK(clk));
DFFX1 gate490(.Q (g1853), .QB (line490), .D(g5672), .CK(clk));
DFFX1 gate491(.Q (g162), .QB (line491), .D(g8424), .CK(clk));
DFFX1 gate492(.Q (g411), .QB (line492), .D(g11268), .CK(clk));
DFFX1 gate493(.Q (g431), .QB (line493), .D(g11262), .CK(clk));
DFFX1 gate494(.Q (g1905), .QB (line494), .D(g8283), .CK(clk));
DFFX1 gate495(.Q (g1515), .QB (line495), .D(g7333), .CK(clk));
DFFX1 gate496(.Q (g1630), .QB (line496), .D(g8872), .CK(clk));
DFFX1 gate497(.Q (g49), .QB (line497), .D(g7774), .CK(clk));
DFFX1 gate498(.Q (g991), .QB (line498), .D(g7802), .CK(clk));
DFFX1 gate499(.Q (g1300), .QB (line499), .D(g7291), .CK(clk));
DFFX1 gate500(.Q (g339), .QB (line500), .D(g11505), .CK(clk));
DFFX1 gate501(.Q (g256), .QB (line501), .D(g7752), .CK(clk));
DFFX1 gate502(.Q (g1750), .QB (line502), .D(g5665), .CK(clk));
DFFX1 gate503(.Q (g585), .QB (line503), .D(g6293), .CK(clk));
DFFX1 gate504(.Q (g1440), .QB (line504), .D(g8988), .CK(clk));
DFFX1 gate505(.Q (g1666), .QB (line505), .D(g11035), .CK(clk));
DFFX1 gate506(.Q (g1528), .QB (line506), .D(g7339), .CK(clk));
DFFX1 gate507(.Q (g1351), .QB (line507), .D(g11657), .CK(clk));
DFFX1 gate508(.Q (g1648), .QB (line508), .D(g11181), .CK(clk));
DFFX1 gate509(.Q (g127), .QB (line509), .D(g8421), .CK(clk));
DFFX1 gate510(.Q (g1618), .QB (line510), .D(g11611), .CK(clk));
DFFX1 gate511(.Q (g1235), .QB (line511), .D(g7296), .CK(clk));
DFFX1 gate512(.Q (g299), .QB (line512), .D(g7772), .CK(clk));
DFFX1 gate513(.Q (g435), .QB (line513), .D(g11261), .CK(clk));
DFFX1 gate514(.Q (g64), .QB (line514), .D(g7781), .CK(clk));
DFFX1 gate515(.Q (g1555), .QB (line515), .D(g7348), .CK(clk));
DFFX1 gate516(.Q (g995), .QB (line516), .D(g7801), .CK(clk));
DFFX1 gate517(.Q (g1621), .QB (line517), .D(g8869), .CK(clk));
DFFX1 gate518(.Q (g1113), .QB (line518), .D(g6313), .CK(clk));
DFFX1 gate519(.Q (g643), .QB (line519), .D(g8064), .CK(clk));
DFFX1 gate520(.Q (g1494), .QB (line520), .D(g8446), .CK(clk));
DFFX1 gate521(.Q (g1567), .QB (line521), .D(g7352), .CK(clk));
DFFX1 gate522(.Q (g691), .QB (line522), .D(g8430), .CK(clk));
DFFX1 gate523(.Q (g534), .QB (line523), .D(g11327), .CK(clk));
DFFX1 gate524(.Q (g1776), .QB (line524), .D(g7812), .CK(clk));
DFFX1 gate525(.Q (g569), .QB (line525), .D(g10876), .CK(clk));
DFFX1 gate526(.Q (g1160), .QB (line526), .D(g6302), .CK(clk));
DFFX1 gate527(.Q (g1360), .QB (line527), .D(g9824), .CK(clk));
DFFX1 gate528(.Q (g1050), .QB (line528), .D(g7791), .CK(clk));
DFFX1 gate529(.Q (g1), .QB (line529), .D(g8078), .CK(clk));
DFFX1 gate530(.Q (g511), .QB (line530), .D(g11336), .CK(clk));
DFFX1 gate531(.Q (g1724), .QB (line531), .D(g10879), .CK(clk));
DFFX1 gate532(.Q (g12), .QB (line532), .D(g7337), .CK(clk));
DFFX1 gate533(.Q (g1878), .QB (line533), .D(g8695), .CK(clk));
DFFX1 gate534(.Q (g73), .QB (line534), .D(g7784), .CK(clk));
INVX1 gate535(.O (I8854), .I (g4500));
INVX1 gate536(.O (g5652), .I (I9117));
INVX1 gate537(.O (I12913), .I (g7845));
INVX1 gate538(.O (g11354), .I (I17179));
INVX1 gate539(.O (g6837), .I (I10891));
INVX1 gate540(.O (I10941), .I (g6555));
INVX1 gate541(.O (I6979), .I (g2888));
INVX1 gate542(.O (g5843), .I (I9458));
INVX1 gate543(.O (g2771), .I (I5854));
INVX1 gate544(.O (g3537), .I (g3164));
INVX1 gate545(.O (g6062), .I (I9699));
INVX1 gate546(.O (I9984), .I (g5529));
INVX1 gate547(.O (I14382), .I (g8886));
INVX1 gate548(.O (g7706), .I (I12335));
INVX1 gate549(.O (I13618), .I (g8345));
INVX1 gate550(.O (I15181), .I (g9968));
INVX1 gate551(.O (g6620), .I (I10573));
INVX1 gate552(.O (I12436), .I (g7659));
INVX1 gate553(.O (g5193), .I (g4682));
INVX1 gate554(.O (g6462), .I (I10394));
INVX1 gate555(.O (g8925), .I (I14252));
INVX1 gate556(.O (I14519), .I (g9106));
INVX1 gate557(.O (g10289), .I (I15691));
INVX1 gate558(.O (I14176), .I (g8784));
INVX1 gate559(.O (I14185), .I (g8790));
INVX1 gate560(.O (g11181), .I (I16944));
INVX1 gate561(.O (I14675), .I (g9263));
INVX1 gate562(.O (g2299), .I (g1707));
INVX1 gate563(.O (I12607), .I (g7633));
INVX1 gate564(.O (g3272), .I (g2450));
INVX1 gate565(.O (g2547), .I (g23));
INVX1 gate566(.O (g9291), .I (g8892));
INVX1 gate567(.O (I6001), .I (g2548));
INVX1 gate568(.O (I7048), .I (g2807));
INVX1 gate569(.O (g10309), .I (I15733));
INVX1 gate570(.O (g7029), .I (I11180));
INVX1 gate571(.O (g4440), .I (g4130));
INVX1 gate572(.O (I9544), .I (g5024));
INVX1 gate573(.O (g10288), .I (I15688));
INVX1 gate574(.O (I12274), .I (g7110));
INVX1 gate575(.O (I9483), .I (g5050));
INVX1 gate576(.O (g7787), .I (I12526));
INVX1 gate577(.O (I6676), .I (g2759));
INVX1 gate578(.O (I8520), .I (g4338));
INVX1 gate579(.O (g10571), .I (I16236));
INVX1 gate580(.O (I17692), .I (g11596));
INVX1 gate581(.O (I17761), .I (g11652));
INVX1 gate582(.O (I13469), .I (g8147));
INVX1 gate583(.O (g9344), .I (I14537));
INVX1 gate584(.O (g7956), .I (g7432));
INVX1 gate585(.O (g3417), .I (I6624));
INVX1 gate586(.O (g4323), .I (g4130));
INVX1 gate587(.O (I11286), .I (g6551));
INVX1 gate588(.O (I8031), .I (g3540));
INVX1 gate589(.O (g7675), .I (I12300));
INVX1 gate590(.O (g8320), .I (I13344));
INVX1 gate591(.O (I12565), .I (g7388));
INVX1 gate592(.O (I16644), .I (g10865));
INVX1 gate593(.O (I11306), .I (g6731));
INVX1 gate594(.O (g1981), .I (g650));
INVX1 gate595(.O (I7333), .I (g3729));
INVX1 gate596(.O (I13039), .I (g8054));
INVX1 gate597(.O (g3982), .I (g3052));
INVX1 gate598(.O (g6249), .I (I10006));
INVX1 gate599(.O (g9259), .I (g8892));
INVX1 gate600(.O (I15190), .I (g9974));
INVX1 gate601(.O (g11426), .I (I17331));
INVX1 gate602(.O (g9819), .I (I14958));
INVX1 gate603(.O (g8277), .I (I13203));
INVX1 gate604(.O (I5050), .I (g1216));
INVX1 gate605(.O (I5641), .I (g546));
INVX1 gate606(.O (g5121), .I (g4682));
INVX1 gate607(.O (g1997), .I (g798));
INVX1 gate608(.O (g3629), .I (g3228));
INVX1 gate609(.O (g3328), .I (I6501));
INVX1 gate610(.O (I12641), .I (g7709));
INVX1 gate611(.O (g5670), .I (I9171));
INVX1 gate612(.O (g6842), .I (I10898));
INVX1 gate613(.O (g8617), .I (g8465));
INVX1 gate614(.O (I15520), .I (g10035));
INVX1 gate615(.O (I7396), .I (g4102));
INVX1 gate616(.O (I7803), .I (g3820));
INVX1 gate617(.O (g3330), .I (I6507));
INVX1 gate618(.O (g2991), .I (I6233));
INVX1 gate619(.O (I9461), .I (g4940));
INVX1 gate620(.O (g2244), .I (I5251));
INVX1 gate621(.O (g6192), .I (I9923));
INVX1 gate622(.O (g6298), .I (I10153));
INVX1 gate623(.O (g6085), .I (I9734));
INVX1 gate624(.O (I12153), .I (g6874));
INVX1 gate625(.O (g4351), .I (I7630));
INVX1 gate626(.O (I11677), .I (g7056));
INVX1 gate627(.O (g10687), .I (I16356));
INVX1 gate628(.O (g4530), .I (I7935));
INVX1 gate629(.O (g8516), .I (I13717));
INVX1 gate630(.O (g5232), .I (g4640));
INVX1 gate631(.O (I13975), .I (g8588));
INVX1 gate632(.O (g2078), .I (g135));
INVX1 gate633(.O (I8911), .I (g4565));
INVX1 gate634(.O (g2340), .I (g1918));
INVX1 gate635(.O (g7684), .I (g7148));
INVX1 gate636(.O (I12409), .I (g7501));
INVX1 gate637(.O (g7745), .I (I12400));
INVX1 gate638(.O (g8987), .I (I14382));
INVX1 gate639(.O (g11546), .I (g11519));
INVX1 gate640(.O (I10729), .I (g5935));
INVX1 gate641(.O (g5253), .I (g4346));
INVX1 gate642(.O (g7338), .I (I11662));
INVX1 gate643(.O (I7509), .I (g3566));
INVX1 gate644(.O (I9427), .I (g4963));
INVX1 gate645(.O (g3800), .I (g3292));
INVX1 gate646(.O (I15088), .I (g9832));
INVX1 gate647(.O (g2907), .I (I6074));
INVX1 gate648(.O (g7791), .I (I12538));
INVX1 gate649(.O (I11143), .I (g6446));
INVX1 gate650(.O (g6854), .I (I10920));
INVX1 gate651(.O (g11088), .I (I16871));
INVX1 gate652(.O (g7309), .I (I11575));
INVX1 gate653(.O (g8299), .I (I13255));
INVX1 gate654(.O (I9046), .I (g4736));
INVX1 gate655(.O (g6941), .I (g6503));
INVX1 gate656(.O (g2435), .I (g201));
INVX1 gate657(.O (I14439), .I (g8969));
INVX1 gate658(.O (g4010), .I (g3144));
INVX1 gate659(.O (g2082), .I (g1371));
INVX1 gate660(.O (I6932), .I (g2850));
INVX1 gate661(.O (I7662), .I (g3336));
INVX1 gate662(.O (I9446), .I (g5052));
INVX1 gate663(.O (g5519), .I (g4811));
INVX1 gate664(.O (g5740), .I (I9302));
INVX1 gate665(.O (I5289), .I (g49));
INVX1 gate666(.O (I9514), .I (g5094));
INVX1 gate667(.O (g7808), .I (I12589));
INVX1 gate668(.O (g2482), .I (I5565));
INVX1 gate669(.O (I5658), .I (g560));
INVX1 gate670(.O (I15497), .I (g10119));
INVX1 gate671(.O (I6624), .I (g2629));
INVX1 gate672(.O (g8892), .I (I14242));
INVX1 gate673(.O (I11169), .I (g6481));
INVX1 gate674(.O (g3213), .I (I6388));
INVX1 gate675(.O (I6068), .I (g2227));
INVX1 gate676(.O (g11497), .I (I17510));
INVX1 gate677(.O (I13791), .I (g8518));
INVX1 gate678(.O (I16867), .I (g10913));
INVX1 gate679(.O (I10349), .I (g6215));
INVX1 gate680(.O (g10260), .I (g10125));
INVX1 gate681(.O (g7759), .I (I12442));
INVX1 gate682(.O (I8473), .I (g4577));
INVX1 gate683(.O (I14349), .I (g8958));
INVX1 gate684(.O (g6708), .I (I10689));
INVX1 gate685(.O (g10668), .I (g10563));
INVX1 gate686(.O (I5271), .I (g70));
INVX1 gate687(.O (I9191), .I (g5546));
INVX1 gate688(.O (I9391), .I (g5013));
INVX1 gate689(.O (g6219), .I (g5426));
INVX1 gate690(.O (I15250), .I (g9980));
INVX1 gate691(.O (I17100), .I (g11221));
INVX1 gate692(.O (I14906), .I (g9508));
INVX1 gate693(.O (g9825), .I (I14976));
INVX1 gate694(.O (g7201), .I (I11427));
INVX1 gate695(.O (I14083), .I (g8747));
INVX1 gate696(.O (g10195), .I (I15559));
INVX1 gate697(.O (I8324), .I (g4794));
INVX1 gate698(.O (g6031), .I (I9642));
INVX1 gate699(.O (g2915), .I (I6094));
INVX1 gate700(.O (I13666), .I (g8292));
INVX1 gate701(.O (I9695), .I (g5212));
INVX1 gate702(.O (I11363), .I (g6595));
INVX1 gate703(.O (I11217), .I (g6529));
INVX1 gate704(.O (g6431), .I (g6145));
INVX1 gate705(.O (g6252), .I (I10015));
INVX1 gate706(.O (g4172), .I (I7333));
INVX1 gate707(.O (g6812), .I (I10846));
INVX1 gate708(.O (g8991), .I (I14394));
INVX1 gate709(.O (g4372), .I (I7677));
INVX1 gate710(.O (g7049), .I (I11228));
INVX1 gate711(.O (I6576), .I (g2617));
INVX1 gate712(.O (g10525), .I (g10499));
INVX1 gate713(.O (g10488), .I (I16101));
INVX1 gate714(.O (I10566), .I (g5904));
INVX1 gate715(.O (I13478), .I (g8191));
INVX1 gate716(.O (g5586), .I (I8996));
INVX1 gate717(.O (g8709), .I (g8674));
INVX1 gate718(.O (g2214), .I (g115));
INVX1 gate719(.O (I9536), .I (g5008));
INVX1 gate720(.O (g6176), .I (I9905));
INVX1 gate721(.O (g4618), .I (g3829));
INVX1 gate722(.O (I15296), .I (g9995));
INVX1 gate723(.O (g4143), .I (I7291));
INVX1 gate724(.O (I7381), .I (g4078));
INVX1 gate725(.O (I9159), .I (g5033));
INVX1 gate726(.O (g11339), .I (I17142));
INVX1 gate727(.O (g8140), .I (I13017));
INVX1 gate728(.O (I16979), .I (g11088));
INVX1 gate729(.O (I16496), .I (g10707));
INVX1 gate730(.O (g8078), .I (I12936));
INVX1 gate731(.O (I7847), .I (g3435));
INVX1 gate732(.O (I9359), .I (g5576));
INVX1 gate733(.O (g8340), .I (I13400));
INVX1 gate734(.O (g2110), .I (I5002));
INVX1 gate735(.O (I15338), .I (g10013));
INVX1 gate736(.O (g6405), .I (g6133));
INVX1 gate737(.O (g8478), .I (I13678));
INVX1 gate738(.O (I16111), .I (g10385));
INVX1 gate739(.O (g4282), .I (g4013));
INVX1 gate740(.O (g11644), .I (I17736));
INVX1 gate741(.O (g7604), .I (I12162));
INVX1 gate742(.O (g9768), .I (g9432));
INVX1 gate743(.O (g4566), .I (g3753));
INVX1 gate744(.O (g7098), .I (I11333));
INVX1 gate745(.O (g10893), .I (I16641));
INVX1 gate746(.O (I4961), .I (g254));
INVX1 gate747(.O (g4988), .I (I8358));
INVX1 gate748(.O (g6286), .I (I10117));
INVX1 gate749(.O (g8959), .I (I14326));
INVX1 gate750(.O (I13580), .I (g8338));
INVX1 gate751(.O (I9016), .I (g4722));
INVX1 gate752(.O (I6398), .I (g2335));
INVX1 gate753(.O (g8517), .I (I13720));
INVX1 gate754(.O (g3348), .I (g2733));
INVX1 gate755(.O (I15060), .I (g9696));
INVX1 gate756(.O (I15968), .I (g10408));
INVX1 gate757(.O (I5332), .I (g756));
INVX1 gate758(.O (g8482), .I (g8329));
INVX1 gate759(.O (g2002), .I (g818));
INVX1 gate760(.O (I10138), .I (g5677));
INVX1 gate761(.O (g11060), .I (g10937));
INVX1 gate762(.O (I17407), .I (g11417));
INVX1 gate763(.O (I12303), .I (g7242));
INVX1 gate764(.O (g5645), .I (I9096));
INVX1 gate765(.O (I15855), .I (g10336));
INVX1 gate766(.O (g2824), .I (I5932));
INVX1 gate767(.O (g11197), .I (g11112));
INVX1 gate768(.O (g4555), .I (I7964));
INVX1 gate769(.O (g5691), .I (g5236));
INVX1 gate770(.O (I9642), .I (g5229));
INVX1 gate771(.O (g7539), .I (I11953));
INVX1 gate772(.O (g7896), .I (I12678));
INVX1 gate773(.O (g8656), .I (I13941));
INVX1 gate774(.O (g9887), .I (I15068));
INVX1 gate775(.O (I8199), .I (g4013));
INVX1 gate776(.O (g6974), .I (g6365));
INVX1 gate777(.O (g6270), .I (I10069));
INVX1 gate778(.O (I14415), .I (g8940));
INVX1 gate779(.O (g3260), .I (I6428));
INVX1 gate780(.O (g11411), .I (I17274));
INVX1 gate781(.O (I10852), .I (g6751));
INVX1 gate782(.O (g10042), .I (I15253));
INVX1 gate783(.O (g10255), .I (g10139));
INVX1 gate784(.O (g6073), .I (I9712));
INVX1 gate785(.O (g10189), .I (I15545));
INVX1 gate786(.O (I4903), .I (g259));
INVX1 gate787(.O (g2877), .I (I6025));
INVX1 gate788(.O (I11531), .I (g7126));
INVX1 gate789(.O (g10679), .I (g10584));
INVX1 gate790(.O (g6796), .I (g6252));
INVX1 gate791(.O (I8900), .I (g4560));
INVX1 gate792(.O (I16735), .I (g10855));
INVX1 gate793(.O (g1968), .I (g369));
INVX1 gate794(.O (g5879), .I (I9498));
INVX1 gate795(.O (I10963), .I (g6793));
INVX1 gate796(.O (g10270), .I (g10156));
INVX1 gate797(.O (g3463), .I (g3256));
INVX1 gate798(.O (g7268), .I (I11505));
INVX1 gate799(.O (g7362), .I (I11734));
INVX1 gate800(.O (I11740), .I (g7030));
INVX1 gate801(.O (g10188), .I (I15542));
INVX1 gate802(.O (I12174), .I (g6939));
INVX1 gate803(.O (I12796), .I (g7543));
INVX1 gate804(.O (g5659), .I (I9138));
INVX1 gate805(.O (g7419), .I (g7206));
INVX1 gate806(.O (I15503), .I (g10044));
INVX1 gate807(.O (I17441), .I (g11445));
INVX1 gate808(.O (g6980), .I (I11127));
INVX1 gate809(.O (I17206), .I (g11323));
INVX1 gate810(.O (g4113), .I (I7255));
INVX1 gate811(.O (g6069), .I (I9706));
INVX1 gate812(.O (g11503), .I (I17528));
INVX1 gate813(.O (g7052), .I (I11235));
INVX1 gate814(.O (g8110), .I (g7996));
INVX1 gate815(.O (g2556), .I (g186));
INVX1 gate816(.O (g4313), .I (g3586));
INVX1 gate817(.O (I16196), .I (g10496));
INVX1 gate818(.O (I7817), .I (g3399));
INVX1 gate819(.O (g8310), .I (I13314));
INVX1 gate820(.O (g10460), .I (I15971));
INVX1 gate821(.O (g2222), .I (g158));
INVX1 gate822(.O (I11953), .I (g6907));
INVX1 gate823(.O (I13373), .I (g8226));
INVX1 gate824(.O (I6818), .I (g2758));
INVX1 gate825(.O (g4202), .I (I7423));
INVX1 gate826(.O (I6867), .I (g2949));
INVX1 gate827(.O (I9880), .I (g5405));
INVX1 gate828(.O (g10093), .I (I15326));
INVX1 gate829(.O (I10484), .I (g6155));
INVX1 gate830(.O (g9845), .I (g9679));
INVX1 gate831(.O (g3720), .I (I6888));
INVX1 gate832(.O (g10267), .I (g10130));
INVX1 gate833(.O (g10294), .I (I15704));
INVX1 gate834(.O (I11800), .I (g7246));
INVX1 gate835(.O (g4908), .I (g4396));
INVX1 gate836(.O (g5111), .I (I8499));
INVX1 gate837(.O (g11450), .I (I17407));
INVX1 gate838(.O (I13800), .I (g8500));
INVX1 gate839(.O (g5275), .I (g4371));
INVX1 gate840(.O (I11417), .I (g6638));
INVX1 gate841(.O (I17758), .I (g11647));
INVX1 gate842(.O (g3318), .I (g2245));
INVX1 gate843(.O (g11315), .I (I17108));
INVX1 gate844(.O (g4094), .I (g2744));
INVX1 gate845(.O (I17435), .I (g11454));
INVX1 gate846(.O (g10065), .I (I15293));
INVX1 gate847(.O (I5092), .I (g32));
INVX1 gate848(.O (g8002), .I (I12832));
INVX1 gate849(.O (g5615), .I (I9043));
INVX1 gate850(.O (g4567), .I (g3374));
INVX1 gate851(.O (I8259), .I (g4590));
INVX1 gate852(.O (g11202), .I (g11112));
INVX1 gate853(.O (g7728), .I (I12369));
INVX1 gate854(.O (g6287), .I (I10120));
INVX1 gate855(.O (I14312), .I (g8814));
INVX1 gate856(.O (I9612), .I (g5149));
INVX1 gate857(.O (g10875), .I (I16595));
INVX1 gate858(.O (I9243), .I (g5245));
INVX1 gate859(.O (g11055), .I (g10950));
INVX1 gate860(.O (g3393), .I (g3144));
INVX1 gate861(.O (g9807), .I (g9490));
INVX1 gate862(.O (g11111), .I (g10974));
INVX1 gate863(.O (g4776), .I (g3586));
INVX1 gate864(.O (I9935), .I (g5477));
INVX1 gate865(.O (g4593), .I (I8004));
INVX1 gate866(.O (I11964), .I (g6910));
INVX1 gate867(.O (I7441), .I (g3473));
INVX1 gate868(.O (I15986), .I (g10417));
INVX1 gate869(.O (g3971), .I (I7104));
INVX1 gate870(.O (g7070), .I (I11289));
INVX1 gate871(.O (g2237), .I (g713));
INVX1 gate872(.O (g6399), .I (I10305));
INVX1 gate873(.O (g5284), .I (g4376));
INVX1 gate874(.O (I11423), .I (g6488));
INVX1 gate875(.O (g7470), .I (g6927));
INVX1 gate876(.O (I15741), .I (g10260));
INVX1 gate877(.O (g7897), .I (g7712));
INVX1 gate878(.O (g7025), .I (g6400));
INVX1 gate879(.O (I6370), .I (g2356));
INVX1 gate880(.O (g7425), .I (g7214));
INVX1 gate881(.O (I11587), .I (g6828));
INVX1 gate882(.O (g2844), .I (I5966));
INVX1 gate883(.O (I12553), .I (g7676));
INVX1 gate884(.O (I12862), .I (g7638));
INVX1 gate885(.O (I8215), .I (g3981));
INVX1 gate886(.O (I10813), .I (g6397));
INVX1 gate887(.O (g11384), .I (I17209));
INVX1 gate888(.O (I14799), .I (g9661));
INVX1 gate889(.O (I6821), .I (g3015));
INVX1 gate890(.O (g2194), .I (g47));
INVX1 gate891(.O (g10160), .I (I15476));
INVX1 gate892(.O (g6797), .I (I10801));
INVX1 gate893(.O (g11067), .I (g10974));
INVX1 gate894(.O (g9342), .I (I14531));
INVX1 gate895(.O (I12326), .I (g7246));
INVX1 gate896(.O (g8928), .I (I14257));
INVX1 gate897(.O (g3121), .I (g2462));
INVX1 gate898(.O (I16280), .I (g10537));
INVX1 gate899(.O (g4160), .I (I7303));
INVX1 gate900(.O (g3321), .I (I6484));
INVX1 gate901(.O (g2089), .I (I4917));
INVX1 gate902(.O (g4933), .I (I8298));
INVX1 gate903(.O (I14973), .I (g9733));
INVX1 gate904(.O (g2731), .I (I5789));
INVX1 gate905(.O (I16688), .I (g10800));
INVX1 gate906(.O (I11543), .I (g6881));
INVX1 gate907(.O (g5420), .I (g4300));
INVX1 gate908(.O (I15801), .I (g10282));
INVX1 gate909(.O (I12948), .I (g8019));
INVX1 gate910(.O (g10455), .I (I15956));
INVX1 gate911(.O (g8064), .I (I12910));
INVX1 gate912(.O (g4521), .I (g3586));
INVX1 gate913(.O (I14805), .I (g9360));
INVX1 gate914(.O (g6291), .I (I10132));
INVX1 gate915(.O (g2557), .I (g1840));
INVX1 gate916(.O (g4050), .I (I7163));
INVX1 gate917(.O (I13117), .I (g7904));
INVX1 gate918(.O (I12904), .I (g7985));
INVX1 gate919(.O (I4873), .I (g105));
INVX1 gate920(.O (g8785), .I (I14090));
INVX1 gate921(.O (g4450), .I (g3914));
INVX1 gate922(.O (g5794), .I (I9394));
INVX1 gate923(.O (g9097), .I (g8892));
INVX1 gate924(.O (g2071), .I (I4873));
INVX1 gate925(.O (g7678), .I (I12307));
INVX1 gate926(.O (g6144), .I (I9857));
INVX1 gate927(.O (I11569), .I (g6821));
INVX1 gate928(.O (g3253), .I (I6417));
INVX1 gate929(.O (I7743), .I (g3762));
INVX1 gate930(.O (g6344), .I (I10251));
INVX1 gate931(.O (g3938), .I (g2991));
INVX1 gate932(.O (g7331), .I (I11641));
INVX1 gate933(.O (I15196), .I (g9974));
INVX1 gate934(.O (g9354), .I (I14567));
INVX1 gate935(.O (g10201), .I (g10175));
INVX1 gate936(.O (g7406), .I (I11786));
INVX1 gate937(.O (g10277), .I (I15675));
INVX1 gate938(.O (g2242), .I (I5245));
INVX1 gate939(.O (I9213), .I (g4944));
INVX1 gate940(.O (g3909), .I (g2920));
INVX1 gate941(.O (I6106), .I (g2116));
INVX1 gate942(.O (g7635), .I (I12245));
INVX1 gate943(.O (I4869), .I (g253));
INVX1 gate944(.O (I13568), .I (g8343));
INVX1 gate945(.O (I13747), .I (g8299));
INVX1 gate946(.O (I15526), .I (g10051));
INVX1 gate947(.O (g8563), .I (I13782));
INVX1 gate948(.O (g10075), .I (I15302));
INVX1 gate949(.O (g4724), .I (g3586));
INVX1 gate950(.O (g6259), .I (I10036));
INVX1 gate951(.O (g4179), .I (I7354));
INVX1 gate952(.O (g7766), .I (I12463));
INVX1 gate953(.O (I5722), .I (g2075));
INVX1 gate954(.O (g7682), .I (g7148));
INVX1 gate955(.O (I13242), .I (g8267));
INVX1 gate956(.O (I17500), .I (g11478));
INVX1 gate957(.O (g6694), .I (I10663));
INVX1 gate958(.O (g4379), .I (g3698));
INVX1 gate959(.O (g3519), .I (g3164));
INVX1 gate960(.O (g7801), .I (I12568));
INVX1 gate961(.O (g7305), .I (I11563));
INVX1 gate962(.O (I7411), .I (g4140));
INVX1 gate963(.O (g8295), .I (I13239));
INVX1 gate964(.O (g2955), .I (I6156));
INVX1 gate965(.O (I8136), .I (g4144));
INVX1 gate966(.O (g5628), .I (I9062));
INVX1 gate967(.O (I6061), .I (g2246));
INVX1 gate968(.O (I12183), .I (g7007));
INVX1 gate969(.O (g6852), .I (I10914));
INVX1 gate970(.O (I11814), .I (g7196));
INVX1 gate971(.O (g5515), .I (g4429));
INVX1 gate972(.O (I6461), .I (g2261));
INVX1 gate973(.O (g5630), .I (I9068));
INVX1 gate974(.O (I12397), .I (g7284));
INVX1 gate975(.O (I4917), .I (g584));
INVX1 gate976(.O (g2254), .I (g131));
INVX1 gate977(.O (g2814), .I (I5916));
INVX1 gate978(.O (g11402), .I (I17249));
INVX1 gate979(.O (g4289), .I (g4013));
INVX1 gate980(.O (g7748), .I (I12409));
INVX1 gate981(.O (g4777), .I (g3992));
INVX1 gate982(.O (I11807), .I (g6854));
INVX1 gate983(.O (g11457), .I (I17424));
INVX1 gate984(.O (I9090), .I (g5567));
INVX1 gate985(.O (g4835), .I (I8192));
INVX1 gate986(.O (I14400), .I (g8891));
INVX1 gate987(.O (g2350), .I (I5424));
INVX1 gate988(.O (g7755), .I (I12430));
INVX1 gate989(.O (g9267), .I (g8892));
INVX1 gate990(.O (g9312), .I (I14509));
INVX1 gate991(.O (I13639), .I (g8321));
INVX1 gate992(.O (g2038), .I (g1776));
INVX1 gate993(.O (I8943), .I (g4585));
INVX1 gate994(.O (I16763), .I (g10890));
INVX1 gate995(.O (I12933), .I (g7899));
INVX1 gate996(.O (g7226), .I (I11464));
INVX1 gate997(.O (g8089), .I (g7934));
INVX1 gate998(.O (g10352), .I (I15820));
INVX1 gate999(.O (g2438), .I (g243));
INVX1 gate1000(.O (I11293), .I (g6516));
INVX1 gate1001(.O (I13230), .I (g8244));
INVX1 gate1002(.O (g2773), .I (I5858));
INVX1 gate1003(.O (g4271), .I (g3971));
INVX1 gate1004(.O (I6904), .I (g2820));
INVX1 gate1005(.O (I12508), .I (g7731));
INVX1 gate1006(.O (I11638), .I (g6948));
INVX1 gate1007(.O (I12634), .I (g7727));
INVX1 gate1008(.O (g10155), .I (I15461));
INVX1 gate1009(.O (I17613), .I (g11550));
INVX1 gate1010(.O (g10822), .I (I16534));
INVX1 gate1011(.O (I4786), .I (g109));
INVX1 gate1012(.O (I6046), .I (g2218));
INVX1 gate1013(.O (I9056), .I (g4753));
INVX1 gate1014(.O (g6951), .I (I11097));
INVX1 gate1015(.O (g10266), .I (g10129));
INVX1 gate1016(.O (I8228), .I (g4468));
INVX1 gate1017(.O (I14005), .I (g8631));
INVX1 gate1018(.O (g10170), .I (g10118));
INVX1 gate1019(.O (I8465), .I (g4807));
INVX1 gate1020(.O (I16660), .I (g10793));
INVX1 gate1021(.O (g7045), .I (g6435));
INVX1 gate1022(.O (I10538), .I (g5910));
INVX1 gate1023(.O (I8934), .I (g4271));
INVX1 gate1024(.O (I5424), .I (g910));
INVX1 gate1025(.O (I5795), .I (g2462));
INVX1 gate1026(.O (g7445), .I (I11845));
INVX1 gate1027(.O (g6114), .I (I9795));
INVX1 gate1028(.O (I5737), .I (g2100));
INVX1 gate1029(.O (I6403), .I (g2337));
INVX1 gate1030(.O (I5809), .I (g2356));
INVX1 gate1031(.O (g6314), .I (I10201));
INVX1 gate1032(.O (I7713), .I (g3750));
INVX1 gate1033(.O (g9761), .I (g9454));
INVX1 gate1034(.O (I11841), .I (g7226));
INVX1 gate1035(.O (I11992), .I (g7058));
INVX1 gate1036(.O (I11391), .I (g6387));
INVX1 gate1037(.O (I9851), .I (g5405));
INVX1 gate1038(.O (g2212), .I (g686));
INVX1 gate1039(.O (I13391), .I (g8178));
INVX1 gate1040(.O (g6870), .I (I10952));
INVX1 gate1041(.O (g4674), .I (I8050));
INVX1 gate1042(.O (g8948), .I (I14299));
INVX1 gate1043(.O (g3141), .I (g2563));
INVX1 gate1044(.O (I6391), .I (g2478));
INVX1 gate1045(.O (I5672), .I (g569));
INVX1 gate1046(.O (I15688), .I (g10207));
INVX1 gate1047(.O (g5040), .I (I8421));
INVX1 gate1048(.O (I5077), .I (g35));
INVX1 gate1049(.O (g1983), .I (g750));
INVX1 gate1050(.O (g6825), .I (I10873));
INVX1 gate1051(.O (g3710), .I (g3215));
INVX1 gate1052(.O (g7369), .I (g7273));
INVX1 gate1053(.O (g7602), .I (I12156));
INVX1 gate1054(.O (g10167), .I (I15497));
INVX1 gate1055(.O (g10194), .I (g10062));
INVX1 gate1056(.O (g10589), .I (I16252));
INVX1 gate1057(.O (I16550), .I (g10726));
INVX1 gate1058(.O (g4541), .I (I7946));
INVX1 gate1059(.O (g7007), .I (I11146));
INVX1 gate1060(.O (I17371), .I (g11410));
INVX1 gate1061(.O (I17234), .I (g11353));
INVX1 gate1062(.O (g7920), .I (g7516));
INVX1 gate1063(.O (I11578), .I (g6824));
INVX1 gate1064(.O (I12574), .I (g7522));
INVX1 gate1065(.O (g10524), .I (g10458));
INVX1 gate1066(.O (g2229), .I (g162));
INVX1 gate1067(.O (I15157), .I (g9931));
INVX1 gate1068(.O (I16307), .I (g10589));
INVX1 gate1069(.O (g4332), .I (g4130));
INVX1 gate1070(.O (I12205), .I (g6993));
INVX1 gate1071(.O (g7767), .I (I12466));
INVX1 gate1072(.O (I6159), .I (g2123));
INVX1 gate1073(.O (g11157), .I (g10950));
INVX1 gate1074(.O (g4680), .I (g3829));
INVX1 gate1075(.O (g6136), .I (I9845));
INVX1 gate1076(.O (g8150), .I (I13039));
INVX1 gate1077(.O (g4209), .I (I7444));
INVX1 gate1078(.O (g4353), .I (I7636));
INVX1 gate1079(.O (g5666), .I (I9159));
INVX1 gate1080(.O (g6336), .I (I10231));
INVX1 gate1081(.O (g8350), .I (I13430));
INVX1 gate1082(.O (I13586), .I (g8356));
INVX1 gate1083(.O (g10119), .I (I15365));
INVX1 gate1084(.O (I8337), .I (g4352));
INVX1 gate1085(.O (g8438), .I (I13612));
INVX1 gate1086(.O (g6594), .I (I10560));
INVX1 gate1087(.O (g11066), .I (g10974));
INVX1 gate1088(.O (g4802), .I (g3337));
INVX1 gate1089(.O (I13442), .I (g8182));
INVX1 gate1090(.O (g8009), .I (I12849));
INVX1 gate1091(.O (I5304), .I (g79));
INVX1 gate1092(.O (g10118), .I (I15362));
INVX1 gate1093(.O (I6016), .I (g2201));
INVX1 gate1094(.O (I6757), .I (g2732));
INVX1 gate1095(.O (g7793), .I (I12544));
INVX1 gate1096(.O (I9279), .I (g5314));
INVX1 gate1097(.O (g5648), .I (I9105));
INVX1 gate1098(.O (g6806), .I (I10828));
INVX1 gate1099(.O (g5875), .I (g5361));
INVX1 gate1100(.O (g6943), .I (I11079));
INVX1 gate1101(.O (I16269), .I (g10558));
INVX1 gate1102(.O (I9720), .I (g5248));
INVX1 gate1103(.O (I12592), .I (g7445));
INVX1 gate1104(.O (g10616), .I (I16289));
INVX1 gate1105(.O (g4558), .I (g3880));
INVX1 gate1106(.O (g5655), .I (I9126));
INVX1 gate1107(.O (I13615), .I (g8333));
INVX1 gate1108(.O (g7415), .I (I11797));
INVX1 gate1109(.O (g7227), .I (I11467));
INVX1 gate1110(.O (I9872), .I (g5557));
INVX1 gate1111(.O (g10313), .I (I15741));
INVX1 gate1112(.O (I5926), .I (g2172));
INVX1 gate1113(.O (I13720), .I (g8358));
INVX1 gate1114(.O (I9652), .I (g5426));
INVX1 gate1115(.O (I5754), .I (g2304));
INVX1 gate1116(.O (I10991), .I (g6759));
INVX1 gate1117(.O (I15763), .I (g10244));
INVX1 gate1118(.O (I11275), .I (g6502));
INVX1 gate1119(.O (g10276), .I (I15672));
INVX1 gate1120(.O (g11511), .I (I17552));
INVX1 gate1121(.O (g4901), .I (I8268));
INVX1 gate1122(.O (I7760), .I (g3768));
INVX1 gate1123(.O (I16670), .I (g10797));
INVX1 gate1124(.O (I11746), .I (g6857));
INVX1 gate1125(.O (I13430), .I (g8241));
INVX1 gate1126(.O (g10305), .I (I15725));
INVX1 gate1127(.O (g10254), .I (g10196));
INVX1 gate1128(.O (g4511), .I (g3586));
INVX1 gate1129(.O (g10900), .I (I16656));
INVX1 gate1130(.O (g9576), .I (I14713));
INVX1 gate1131(.O (g2837), .I (g2130));
INVX1 gate1132(.O (g10466), .I (I15989));
INVX1 gate1133(.O (g5884), .I (I9505));
INVX1 gate1134(.O (I5044), .I (g1182));
INVX1 gate1135(.O (g6433), .I (I10349));
INVX1 gate1136(.O (g5839), .I (I9452));
INVX1 gate1137(.O (g8229), .I (g7826));
INVX1 gate1138(.O (I6654), .I (g2952));
INVX1 gate1139(.O (g8993), .I (I14400));
INVX1 gate1140(.O (g2620), .I (g1998));
INVX1 gate1141(.O (I12846), .I (g7685));
INVX1 gate1142(.O (g2462), .I (I5555));
INVX1 gate1143(.O (g9349), .I (I14552));
INVX1 gate1144(.O (I8815), .I (g4471));
INVX1 gate1145(.O (g10101), .I (I15335));
INVX1 gate1146(.O (g10177), .I (I15523));
INVX1 gate1147(.O (I16667), .I (g10780));
INVX1 gate1148(.O (I13806), .I (g8478));
INVX1 gate1149(.O (I7220), .I (g3213));
INVX1 gate1150(.O (I5862), .I (g2537));
INVX1 gate1151(.O (I9598), .I (g5120));
INVX1 gate1152(.O (I7779), .I (g3774));
INVX1 gate1153(.O (I17724), .I (g11625));
INVX1 gate1154(.O (g6845), .I (I10907));
INVX1 gate1155(.O (g7502), .I (I11882));
INVX1 gate1156(.O (I8154), .I (g3636));
INVX1 gate1157(.O (I10584), .I (g5864));
INVX1 gate1158(.O (I17359), .I (g11372));
INVX1 gate1159(.O (g3545), .I (I6733));
INVX1 gate1160(.O (I15314), .I (g10007));
INVX1 gate1161(.O (g11550), .I (I17591));
INVX1 gate1162(.O (I15287), .I (g9980));
INVX1 gate1163(.O (g6195), .I (g5426));
INVX1 gate1164(.O (I7423), .I (g3331));
INVX1 gate1165(.O (g6137), .I (I9848));
INVX1 gate1166(.O (g5667), .I (I9162));
INVX1 gate1167(.O (g6395), .I (I10293));
INVX1 gate1168(.O (g3380), .I (I6576));
INVX1 gate1169(.O (g5143), .I (g4682));
INVX1 gate1170(.O (g6337), .I (I10234));
INVX1 gate1171(.O (I16487), .I (g10771));
INVX1 gate1172(.O (g6913), .I (I11021));
INVX1 gate1173(.O (g10064), .I (I15290));
INVX1 gate1174(.O (g11287), .I (g11207));
INVX1 gate1175(.O (I15085), .I (g9720));
INVX1 gate1176(.O (g2249), .I (g127));
INVX1 gate1177(.O (I9625), .I (g5405));
INVX1 gate1178(.O (g4580), .I (g3880));
INVX1 gate1179(.O (I10759), .I (g5803));
INVX1 gate1180(.O (g11307), .I (I17092));
INVX1 gate1181(.O (g11076), .I (I16843));
INVX1 gate1182(.O (I9232), .I (g4944));
INVX1 gate1183(.O (g7188), .I (I11408));
INVX1 gate1184(.O (g7689), .I (I12322));
INVX1 gate1185(.O (I17121), .I (g11231));
INVX1 gate1186(.O (g11596), .I (g11580));
INVX1 gate1187(.O (g7388), .I (I11773));
INVX1 gate1188(.O (I10114), .I (g5768));
INVX1 gate1189(.O (I9253), .I (g5052));
INVX1 gate1190(.O (I9938), .I (g5478));
INVX1 gate1191(.O (g10874), .I (I16592));
INVX1 gate1192(.O (g11054), .I (g10950));
INVX1 gate1193(.O (g6807), .I (I10831));
INVX1 gate1194(.O (I9813), .I (g5241));
INVX1 gate1195(.O (I6417), .I (g2344));
INVX1 gate1196(.O (g5693), .I (I9224));
INVX1 gate1197(.O (g11243), .I (g11112));
INVX1 gate1198(.O (I17344), .I (g11369));
INVX1 gate1199(.O (g3507), .I (g3307));
INVX1 gate1200(.O (g4262), .I (g4013));
INVX1 gate1201(.O (g2298), .I (I5336));
INVX1 gate1202(.O (g2085), .I (I4903));
INVX1 gate1203(.O (I7665), .I (g3732));
INVX1 gate1204(.O (g10630), .I (I16311));
INVX1 gate1205(.O (g11431), .I (I17344));
INVX1 gate1206(.O (g6859), .I (I10937));
INVX1 gate1207(.O (g7028), .I (g6407));
INVX1 gate1208(.O (I6982), .I (g2889));
INVX1 gate1209(.O (g6266), .I (I10057));
INVX1 gate1210(.O (I15269), .I (g9993));
INVX1 gate1211(.O (g10166), .I (I15494));
INVX1 gate1212(.O (g7030), .I (I11183));
INVX1 gate1213(.O (I12583), .I (g7546));
INVX1 gate1214(.O (I9519), .I (g4998));
INVX1 gate1215(.O (g8062), .I (I12904));
INVX1 gate1216(.O (g7430), .I (g7221));
INVX1 gate1217(.O (I15341), .I (g10019));
INVX1 gate1218(.O (I5414), .I (g904));
INVX1 gate1219(.O (I16286), .I (g10540));
INVX1 gate1220(.O (I7999), .I (g4114));
INVX1 gate1221(.O (g2854), .I (I5986));
INVX1 gate1222(.O (I17173), .I (g11293));
INVX1 gate1223(.O (I5946), .I (g2176));
INVX1 gate1224(.O (I10849), .I (g6734));
INVX1 gate1225(.O (g11341), .I (I17146));
INVX1 gate1226(.O (I7633), .I (g3474));
INVX1 gate1227(.O (g4889), .I (I8240));
INVX1 gate1228(.O (g2941), .I (I6118));
INVX1 gate1229(.O (g6248), .I (I10003));
INVX1 gate1230(.O (g11655), .I (I17767));
INVX1 gate1231(.O (g9258), .I (g8892));
INVX1 gate1232(.O (g3905), .I (g2920));
INVX1 gate1233(.O (g10892), .I (I16638));
INVX1 gate1234(.O (g9818), .I (I14955));
INVX1 gate1235(.O (g9352), .I (I14561));
INVX1 gate1236(.O (I7303), .I (g3262));
INVX1 gate1237(.O (I8293), .I (g4779));
INVX1 gate1238(.O (I10398), .I (g5820));
INVX1 gate1239(.O (I13475), .I (g8173));
INVX1 gate1240(.O (g11180), .I (I16941));
INVX1 gate1241(.O (g7826), .I (I12627));
INVX1 gate1242(.O (g3628), .I (g3111));
INVX1 gate1243(.O (g6255), .I (I10024));
INVX1 gate1244(.O (g4175), .I (I7342));
INVX1 gate1245(.O (g6081), .I (g4977));
INVX1 gate1246(.O (g6815), .I (I10855));
INVX1 gate1247(.O (I10141), .I (g5683));
INVX1 gate1248(.O (g4375), .I (g3638));
INVX1 gate1249(.O (I10804), .I (g6388));
INVX1 gate1250(.O (I5513), .I (g255));
INVX1 gate1251(.O (g3630), .I (I6789));
INVX1 gate1252(.O (g8788), .I (I14097));
INVX1 gate1253(.O (I11222), .I (g6533));
INVX1 gate1254(.O (I12282), .I (g7113));
INVX1 gate1255(.O (I15335), .I (g10007));
INVX1 gate1256(.O (I16601), .I (g10806));
INVX1 gate1257(.O (g5113), .I (I8503));
INVX1 gate1258(.O (g6692), .I (I10659));
INVX1 gate1259(.O (I16187), .I (g10492));
INVX1 gate1260(.O (g6097), .I (I9754));
INVX1 gate1261(.O (I7732), .I (g3758));
INVX1 gate1262(.O (g7910), .I (g7460));
INVX1 gate1263(.O (I12357), .I (g7147));
INVX1 gate1264(.O (g2219), .I (g94));
INVX1 gate1265(.O (g9893), .I (I15082));
INVX1 gate1266(.O (g2640), .I (g1984));
INVX1 gate1267(.O (g6154), .I (I9875));
INVX1 gate1268(.O (g4285), .I (g3688));
INVX1 gate1269(.O (g6354), .I (g5867));
INVX1 gate1270(.O (g2031), .I (g1690));
INVX1 gate1271(.O (g10907), .I (I16673));
INVX1 gate1272(.O (g5202), .I (g4640));
INVX1 gate1273(.O (g6960), .I (I11112));
INVX1 gate1274(.O (I15694), .I (g10234));
INVX1 gate1275(.O (I5378), .I (g1857));
INVX1 gate1276(.O (g2431), .I (I5510));
INVX1 gate1277(.O (I15965), .I (g10405));
INVX1 gate1278(.O (g2252), .I (I5271));
INVX1 gate1279(.O (g2812), .I (g2158));
INVX1 gate1280(.O (I7240), .I (g2824));
INVX1 gate1281(.O (g7609), .I (I12177));
INVX1 gate1282(.O (I10135), .I (g6249));
INVX1 gate1283(.O (g7308), .I (I11572));
INVX1 gate1284(.O (g8192), .I (I13117));
INVX1 gate1285(.O (g2958), .I (I6163));
INVX1 gate1286(.O (g8085), .I (g7932));
INVX1 gate1287(.O (g10074), .I (I15299));
INVX1 gate1288(.O (g5094), .I (I8462));
INVX1 gate1289(.O (I13347), .I (g8122));
INVX1 gate1290(.O (g2176), .I (g82));
INVX1 gate1291(.O (g9026), .I (I14415));
INVX1 gate1292(.O (g8485), .I (g8341));
INVX1 gate1293(.O (g4184), .I (I7369));
INVX1 gate1294(.O (g5494), .I (g4412));
INVX1 gate1295(.O (g3750), .I (I6941));
INVX1 gate1296(.O (g2005), .I (g928));
INVX1 gate1297(.O (g7883), .I (g7689));
INVX1 gate1298(.O (I7043), .I (g2908));
INVX1 gate1299(.O (g4384), .I (I7707));
INVX1 gate1300(.O (I9141), .I (g5402));
INVX1 gate1301(.O (I9860), .I (g5405));
INVX1 gate1302(.O (g5567), .I (I8982));
INVX1 gate1303(.O (g4339), .I (g4144));
INVX1 gate1304(.O (I9341), .I (g5013));
INVX1 gate1305(.O (g10238), .I (g10191));
INVX1 gate1306(.O (I16169), .I (g10448));
INVX1 gate1307(.O (I9525), .I (g5001));
INVX1 gate1308(.O (I14361), .I (g8951));
INVX1 gate1309(.O (g2829), .I (I5943));
INVX1 gate1310(.O (g11619), .I (I17675));
INVX1 gate1311(.O (g2765), .I (g2184));
INVX1 gate1312(.O (g9821), .I (I14964));
INVX1 gate1313(.O (g11502), .I (I17525));
INVX1 gate1314(.O (g7758), .I (I12439));
INVX1 gate1315(.O (I5916), .I (g2217));
INVX1 gate1316(.O (I13236), .I (g8245));
INVX1 gate1317(.O (g7066), .I (I11275));
INVX1 gate1318(.O (g7589), .I (I12099));
INVX1 gate1319(.O (g4424), .I (g3688));
INVX1 gate1320(.O (g3040), .I (g2135));
INVX1 gate1321(.O (g4737), .I (g3440));
INVX1 gate1322(.O (I11351), .I (g6698));
INVX1 gate1323(.O (I13952), .I (g8451));
INVX1 gate1324(.O (g5593), .I (I9013));
INVX1 gate1325(.O (g6112), .I (I9789));
INVX1 gate1326(.O (I13351), .I (g8214));
INVX1 gate1327(.O (g6218), .I (I9965));
INVX1 gate1328(.O (g6267), .I (I10060));
INVX1 gate1329(.O (g3440), .I (g3041));
INVX1 gate1330(.O (g6312), .I (I10195));
INVX1 gate1331(.O (g11618), .I (I17672));
INVX1 gate1332(.O (g9984), .I (I15184));
INVX1 gate1333(.O (I11821), .I (g7205));
INVX1 gate1334(.O (g10176), .I (I15520));
INVX1 gate1335(.O (g10185), .I (g10040));
INVX1 gate1336(.O (g10675), .I (g10574));
INVX1 gate1337(.O (I16479), .I (g10767));
INVX1 gate1338(.O (g10092), .I (I15323));
INVX1 gate1339(.O (I10048), .I (g5734));
INVX1 gate1340(.O (I16363), .I (g10599));
INVX1 gate1341(.O (I16217), .I (g10501));
INVX1 gate1342(.O (g3323), .I (g2157));
INVX1 gate1343(.O (I15278), .I (g10033));
INVX1 gate1344(.O (g7571), .I (I12035));
INVX1 gate1345(.O (g7365), .I (I11743));
INVX1 gate1346(.O (g2733), .I (I5795));
INVX1 gate1347(.O (g4077), .I (I7202));
INVX1 gate1348(.O (g6001), .I (I9625));
INVX1 gate1349(.O (g7048), .I (I11225));
INVX1 gate1350(.O (g10154), .I (I15458));
INVX1 gate1351(.O (g2270), .I (I5311));
INVX1 gate1352(.O (I5798), .I (g2085));
INVX1 gate1353(.O (I17240), .I (g11395));
INVX1 gate1354(.O (g7711), .I (I12344));
INVX1 gate1355(.O (g4523), .I (g3546));
INVX1 gate1356(.O (I10221), .I (g6117));
INVX1 gate1357(.O (I11790), .I (g7246));
INVX1 gate1358(.O (g8520), .I (I13729));
INVX1 gate1359(.O (g6293), .I (I10138));
INVX1 gate1360(.O (g11469), .I (I17444));
INVX1 gate1361(.O (g8219), .I (g7826));
INVX1 gate1362(.O (g2225), .I (I5210));
INVX1 gate1363(.O (g8640), .I (g8512));
INVX1 gate1364(.O (g10935), .I (g10827));
INVX1 gate1365(.O (g2610), .I (I5731));
INVX1 gate1366(.O (g2073), .I (I4879));
INVX1 gate1367(.O (g2796), .I (g2276));
INVX1 gate1368(.O (g11468), .I (I17441));
INVX1 gate1369(.O (g11039), .I (I16778));
INVX1 gate1370(.O (I6851), .I (g2937));
INVX1 gate1371(.O (g4205), .I (I7432));
INVX1 gate1372(.O (I7697), .I (g3743));
INVX1 gate1373(.O (I10613), .I (g6000));
INVX1 gate1374(.O (I11873), .I (g6863));
INVX1 gate1375(.O (g10883), .I (g10809));
INVX1 gate1376(.O (I17755), .I (g11646));
INVX1 gate1377(.O (g7333), .I (I11647));
INVX1 gate1378(.O (g9106), .I (I14439));
INVX1 gate1379(.O (I7210), .I (g2798));
INVX1 gate1380(.O (g7774), .I (I12487));
INVX1 gate1381(.O (g5521), .I (g4530));
INVX1 gate1382(.O (g3528), .I (g3164));
INVX1 gate1383(.O (g8958), .I (I14323));
INVX1 gate1384(.O (I16580), .I (g10826));
INVX1 gate1385(.O (I17770), .I (g11649));
INVX1 gate1386(.O (g11038), .I (I16775));
INVX1 gate1387(.O (g5050), .I (I8429));
INVX1 gate1388(.O (g2124), .I (I5050));
INVX1 gate1389(.O (g3351), .I (I6535));
INVX1 gate1390(.O (g5641), .I (I9084));
INVX1 gate1391(.O (I17563), .I (g11492));
INVX1 gate1392(.O (g2980), .I (g1983));
INVX1 gate1393(.O (g6727), .I (g5997));
INVX1 gate1394(.O (g8376), .I (I13478));
INVX1 gate1395(.O (I5632), .I (g932));
INVX1 gate1396(.O (I5095), .I (g37));
INVX1 gate1397(.O (I6260), .I (g2025));
INVX1 gate1398(.O (g2069), .I (I4869));
INVX1 gate1399(.O (I9111), .I (g5596));
INVX1 gate1400(.O (g7196), .I (I11420));
INVX1 gate1401(.O (g4551), .I (g3946));
INVX1 gate1402(.O (I15601), .I (g10173));
INVX1 gate1403(.O (I9311), .I (g4915));
INVX1 gate1404(.O (I15187), .I (g9968));
INVX1 gate1405(.O (g7803), .I (I12574));
INVX1 gate1406(.O (I12248), .I (g7098));
INVX1 gate1407(.O (I13209), .I (g8198));
INVX1 gate1408(.O (g4499), .I (g3546));
INVX1 gate1409(.O (I8848), .I (g4490));
INVX1 gate1410(.O (g2540), .I (I5655));
INVX1 gate1411(.O (g7538), .I (I11950));
INVX1 gate1412(.O (I13834), .I (g8488));
INVX1 gate1413(.O (I5579), .I (g1197));
INVX1 gate1414(.O (g7780), .I (I12505));
INVX1 gate1415(.O (g5724), .I (I9268));
INVX1 gate1416(.O (g9027), .I (I14418));
INVX1 gate1417(.O (g2206), .I (I5171));
INVX1 gate1418(.O (I12779), .I (g7608));
INVX1 gate1419(.O (g10729), .I (g10630));
INVX1 gate1420(.O (g6703), .I (I10678));
INVX1 gate1421(.O (I9174), .I (g4903));
INVX1 gate1422(.O (I5719), .I (g2072));
INVX1 gate1423(.O (g10577), .I (g10526));
INVX1 gate1424(.O (I17767), .I (g11648));
INVX1 gate1425(.O (g7509), .I (I11889));
INVX1 gate1426(.O (g9427), .I (g9079));
INVX1 gate1427(.O (I10033), .I (g5693));
INVX1 gate1428(.O (I7820), .I (g3811));
INVX1 gate1429(.O (I10234), .I (g6114));
INVX1 gate1430(.O (g4754), .I (g3440));
INVX1 gate1431(.O (I16531), .I (g10720));
INVX1 gate1432(.O (g10439), .I (g10334));
INVX1 gate1433(.O (I11021), .I (g6398));
INVX1 gate1434(.O (I12081), .I (g6934));
INVX1 gate1435(.O (g5878), .I (g5309));
INVX1 gate1436(.O (g6932), .I (I11058));
INVX1 gate1437(.O (g7662), .I (I12279));
INVX1 gate1438(.O (g4273), .I (g4013));
INVX1 gate1439(.O (I16178), .I (g10490));
INVX1 gate1440(.O (I12786), .I (g7622));
INVX1 gate1441(.O (I17633), .I (g11578));
INVX1 gate1442(.O (g5658), .I (I9135));
INVX1 gate1443(.O (g5777), .I (I9365));
INVX1 gate1444(.O (I10795), .I (g6123));
INVX1 gate1445(.O (I13726), .I (g8375));
INVX1 gate1446(.O (g7467), .I (g7148));
INVX1 gate1447(.O (g1990), .I (g774));
INVX1 gate1448(.O (I6118), .I (g2248));
INVX1 gate1449(.O (g8225), .I (g7826));
INVX1 gate1450(.O (I17191), .I (g11315));
INVX1 gate1451(.O (I17719), .I (g11623));
INVX1 gate1452(.O (I11614), .I (g6838));
INVX1 gate1453(.O (g8610), .I (g8483));
INVX1 gate1454(.O (I6367), .I (g2045));
INVX1 gate1455(.O (I9180), .I (g4905));
INVX1 gate1456(.O (I12647), .I (g7711));
INVX1 gate1457(.O (I16676), .I (g10798));
INVX1 gate1458(.O (I16685), .I (g10785));
INVX1 gate1459(.O (I11436), .I (g6488));
INVX1 gate1460(.O (I9380), .I (g5013));
INVX1 gate1461(.O (g10349), .I (I15811));
INVX1 gate1462(.O (g9345), .I (I14540));
INVX1 gate1463(.O (I16953), .I (g11082));
INVX1 gate1464(.O (I13436), .I (g8187));
INVX1 gate1465(.O (I9591), .I (g5095));
INVX1 gate1466(.O (I16373), .I (g10593));
INVX1 gate1467(.O (g4444), .I (I7800));
INVX1 gate1468(.O (g8473), .I (I13669));
INVX1 gate1469(.O (g2199), .I (g48));
INVX1 gate1470(.O (g11410), .I (I17271));
INVX1 gate1471(.O (g2399), .I (g605));
INVX1 gate1472(.O (g9763), .I (I14906));
INVX1 gate1473(.O (g7093), .I (I11326));
INVX1 gate1474(.O (I12999), .I (g7844));
INVX1 gate1475(.O (g3372), .I (g3121));
INVX1 gate1476(.O (I10514), .I (g6154));
INVX1 gate1477(.O (I12380), .I (g7204));
INVX1 gate1478(.O (g10906), .I (I16670));
INVX1 gate1479(.O (I15479), .I (g10091));
INVX1 gate1480(.O (I13320), .I (g8096));
INVX1 gate1481(.O (g10083), .I (I15311));
INVX1 gate1482(.O (I9020), .I (g4773));
INVX1 gate1483(.O (g8124), .I (g8011));
INVX1 gate1484(.O (g10284), .I (g10167));
INVX1 gate1485(.O (g7256), .I (I11489));
INVX1 gate1486(.O (g8980), .I (I14361));
INVX1 gate1487(.O (g7816), .I (I12613));
INVX1 gate1488(.O (g8324), .I (I13354));
INVX1 gate1489(.O (g11479), .I (I17470));
INVX1 gate1490(.O (I6193), .I (g2155));
INVX1 gate1491(.O (I11593), .I (g6830));
INVX1 gate1492(.O (g3143), .I (I6363));
INVX1 gate1493(.O (g11363), .I (I17188));
INVX1 gate1494(.O (g3343), .I (g2779));
INVX1 gate1495(.O (I11122), .I (g6450));
INVX1 gate1496(.O (g2797), .I (g2524));
INVX1 gate1497(.O (I13122), .I (g7966));
INVX1 gate1498(.O (I6549), .I (g2838));
INVX1 gate1499(.O (g4543), .I (g3946));
INVX1 gate1500(.O (I10421), .I (g5826));
INVX1 gate1501(.O (I11464), .I (g6443));
INVX1 gate1502(.O (g3566), .I (I6738));
INVX1 gate1503(.O (I6971), .I (g2882));
INVX1 gate1504(.O (g6716), .I (g5949));
INVX1 gate1505(.O (I14421), .I (g8944));
INVX1 gate1506(.O (g2245), .I (I5254));
INVX1 gate1507(.O (g6149), .I (I9866));
INVX1 gate1508(.O (g3988), .I (g3121));
INVX1 gate1509(.O (I6686), .I (g3015));
INVX1 gate1510(.O (g6349), .I (I10258));
INVX1 gate1511(.O (g7847), .I (I12638));
INVX1 gate1512(.O (g3693), .I (g2920));
INVX1 gate1513(.O (I11034), .I (g6629));
INVX1 gate1514(.O (I10012), .I (g5543));
INVX1 gate1515(.O (g3334), .I (I6517));
INVX1 gate1516(.O (I5725), .I (g2079));
INVX1 gate1517(.O (g7685), .I (g7148));
INVX1 gate1518(.O (g7197), .I (I11423));
INVX1 gate1519(.O (I11641), .I (g6960));
INVX1 gate1520(.O (I11797), .I (g6852));
INVX1 gate1521(.O (g5997), .I (I9617));
INVX1 gate1522(.O (I15580), .I (g10155));
INVX1 gate1523(.O (I13797), .I (g8473));
INVX1 gate1524(.O (I6598), .I (g2623));
INVX1 gate1525(.O (g7021), .I (I11162));
INVX1 gate1526(.O (g4729), .I (g3586));
INVX1 gate1527(.O (g4961), .I (I8333));
INVX1 gate1528(.O (g7421), .I (I11807));
INVX1 gate1529(.O (g10139), .I (I15415));
INVX1 gate1530(.O (g2344), .I (I5410));
INVX1 gate1531(.O (I8211), .I (g3566));
INVX1 gate1532(.O (I9905), .I (g5300));
INVX1 gate1533(.O (g6398), .I (I10302));
INVX1 gate1534(.O (I10541), .I (g6176));
INVX1 gate1535(.O (I6121), .I (g2121));
INVX1 gate1536(.O (g1963), .I (g110));
INVX1 gate1537(.O (I17324), .I (g11347));
INVX1 gate1538(.O (g7263), .I (I11498));
INVX1 gate1539(.O (I14473), .I (g8921));
INVX1 gate1540(.O (g2207), .I (I5174));
INVX1 gate1541(.O (g10138), .I (I15412));
INVX1 gate1542(.O (I17701), .I (g11617));
INVX1 gate1543(.O (I10789), .I (g5867));
INVX1 gate1544(.O (I12448), .I (g7530));
INVX1 gate1545(.O (I13409), .I (g8141));
INVX1 gate1546(.O (I17534), .I (g11495));
INVX1 gate1547(.O (g3792), .I (I7017));
INVX1 gate1548(.O (g5353), .I (I8820));
INVX1 gate1549(.O (g8849), .I (g8745));
INVX1 gate1550(.O (g2259), .I (I5292));
INVX1 gate1551(.O (g6241), .I (I9992));
INVX1 gate1552(.O (g2819), .I (g2159));
INVX1 gate1553(.O (I11408), .I (g6405));
INVX1 gate1554(.O (I12505), .I (g7728));
INVX1 gate1555(.O (I11635), .I (g6947));
INVX1 gate1556(.O (I10724), .I (g6096));
INVX1 gate1557(.O (g11084), .I (I16863));
INVX1 gate1558(.O (g4885), .I (I8228));
INVX1 gate1559(.O (g4414), .I (I7752));
INVX1 gate1560(.O (I10325), .I (g6003));
INVX1 gate1561(.O (g11110), .I (g10974));
INVX1 gate1562(.O (g3621), .I (I6754));
INVX1 gate1563(.O (I6938), .I (g2854));
INVX1 gate1564(.O (I7668), .I (g3733));
INVX1 gate1565(.O (g2852), .I (I5982));
INVX1 gate1566(.O (I7840), .I (g3431));
INVX1 gate1567(.O (I16543), .I (g10747));
INVX1 gate1568(.O (g10852), .I (g10740));
INVX1 gate1569(.O (g8781), .I (I14080));
INVX1 gate1570(.O (I8614), .I (g4414));
INVX1 gate1571(.O (I10920), .I (g6733));
INVX1 gate1572(.O (I10535), .I (g5867));
INVX1 gate1573(.O (I12026), .I (g7119));
INVX1 gate1574(.O (I10434), .I (g5843));
INVX1 gate1575(.O (g11179), .I (I16938));
INVX1 gate1576(.O (g2701), .I (g2040));
INVX1 gate1577(.O (g3113), .I (I6343));
INVX1 gate1578(.O (g7562), .I (g6984));
INVX1 gate1579(.O (I14358), .I (g8950));
INVX1 gate1580(.O (I7390), .I (g4087));
INVX1 gate1581(.O (I10828), .I (g6708));
INVX1 gate1582(.O (I10946), .I (g6548));
INVX1 gate1583(.O (g8797), .I (I14116));
INVX1 gate1584(.O (g6644), .I (I10601));
INVX1 gate1585(.O (g4513), .I (g3546));
INVX1 gate1586(.O (g7631), .I (I12235));
INVX1 gate1587(.O (I5171), .I (g1419));
INVX1 gate1588(.O (g7723), .I (I12354));
INVX1 gate1589(.O (g6119), .I (I9810));
INVX1 gate1590(.O (I9973), .I (g5502));
INVX1 gate1591(.O (g7817), .I (I12616));
INVX1 gate1592(.O (g5901), .I (g5361));
INVX1 gate1593(.O (I4920), .I (g260));
INVX1 gate1594(.O (g8291), .I (I13227));
INVX1 gate1595(.O (g11373), .I (I17198));
INVX1 gate1596(.O (g3094), .I (I6302));
INVX1 gate1597(.O (g6258), .I (I10033));
INVX1 gate1598(.O (g4178), .I (I7351));
INVX1 gate1599(.O (g4436), .I (g3638));
INVX1 gate1600(.O (g6818), .I (I10864));
INVX1 gate1601(.O (g4679), .I (g4013));
INVX1 gate1602(.O (g11654), .I (I17764));
INVX1 gate1603(.O (g4378), .I (I7697));
INVX1 gate1604(.O (g7605), .I (I12165));
INVX1 gate1605(.O (g5511), .I (I8934));
INVX1 gate1606(.O (I11575), .I (g6823));
INVX1 gate1607(.O (g3518), .I (g3164));
INVX1 gate1608(.O (I10682), .I (g6051));
INVX1 gate1609(.O (g10576), .I (g10524));
INVX1 gate1610(.O (I9040), .I (g4794));
INVX1 gate1611(.O (g8144), .I (I13027));
INVX1 gate1612(.O (g8344), .I (I13412));
INVX1 gate1613(.O (g6717), .I (I10706));
INVX1 gate1614(.O (I9440), .I (g5078));
INVX1 gate1615(.O (g11417), .I (I17302));
INVX1 gate1616(.O (I13711), .I (g8342));
INVX1 gate1617(.O (I16814), .I (g10910));
INVX1 gate1618(.O (I12433), .I (g7657));
INVX1 gate1619(.O (g4335), .I (I7612));
INVX1 gate1620(.O (I9123), .I (g4890));
INVX1 gate1621(.O (I11109), .I (g6464));
INVX1 gate1622(.O (g7751), .I (I12418));
INVX1 gate1623(.O (g4182), .I (I7363));
INVX1 gate1624(.O (I9323), .I (g5620));
INVX1 gate1625(.O (I13109), .I (g7981));
INVX1 gate1626(.O (g4288), .I (g4130));
INVX1 gate1627(.O (I11537), .I (g7144));
INVX1 gate1628(.O (g4382), .I (g3638));
INVX1 gate1629(.O (I16772), .I (g10887));
INVX1 gate1630(.O (g3776), .I (g2579));
INVX1 gate1631(.O (g6893), .I (I10991));
INVX1 gate1632(.O (g5574), .I (g4300));
INVX1 gate1633(.O (g5864), .I (I9483));
INVX1 gate1634(.O (g10200), .I (g10169));
INVX1 gate1635(.O (g8694), .I (I13975));
INVX1 gate1636(.O (g2825), .I (I5935));
INVX1 gate1637(.O (g2650), .I (g2006));
INVX1 gate1638(.O (g10608), .I (I16283));
INVX1 gate1639(.O (g10115), .I (I15353));
INVX1 gate1640(.O (g6386), .I (I10282));
INVX1 gate1641(.O (g7585), .I (I12081));
INVX1 gate1642(.O (I17447), .I (g11457));
INVX1 gate1643(.O (I5684), .I (g572));
INVX1 gate1644(.O (I8061), .I (g3381));
INVX1 gate1645(.O (g4805), .I (g3337));
INVX1 gate1646(.O (I7163), .I (g2643));
INVX1 gate1647(.O (I5963), .I (g2179));
INVX1 gate1648(.O (I7810), .I (g3799));
INVX1 gate1649(.O (g7041), .I (g6427));
INVX1 gate1650(.O (I7363), .I (g4005));
INVX1 gate1651(.O (I16638), .I (g10863));
INVX1 gate1652(.O (g2008), .I (g971));
INVX1 gate1653(.O (I13606), .I (g8311));
INVX1 gate1654(.O (I12971), .I (g8039));
INVX1 gate1655(.O (I11303), .I (g6526));
INVX1 gate1656(.O (g6274), .I (I10081));
INVX1 gate1657(.O (I7432), .I (g3663));
INVX1 gate1658(.O (g6426), .I (I10340));
INVX1 gate1659(.O (g11423), .I (I17324));
INVX1 gate1660(.O (g2336), .I (g1900));
INVX1 gate1661(.O (I16416), .I (g10664));
INVX1 gate1662(.O (I12369), .I (g7189));
INVX1 gate1663(.O (I9875), .I (g5278));
INVX1 gate1664(.O (I7453), .I (g3708));
INVX1 gate1665(.O (g6170), .I (g5426));
INVX1 gate1666(.O (I14506), .I (g8923));
INVX1 gate1667(.O (g7673), .I (I12296));
INVX1 gate1668(.O (I9655), .I (g5173));
INVX1 gate1669(.O (g6125), .I (I9822));
INVX1 gate1670(.O (I5707), .I (g2418));
INVX1 gate1671(.O (g8886), .I (I14228));
INVX1 gate1672(.O (g3521), .I (g3164));
INVX1 gate1673(.O (g8951), .I (I14306));
INVX1 gate1674(.O (I16510), .I (g10712));
INVX1 gate1675(.O (g5262), .I (g4353));
INVX1 gate1676(.O (g3050), .I (I6260));
INVX1 gate1677(.O (I11091), .I (g6657));
INVX1 gate1678(.O (g10973), .I (I16720));
INVX1 gate1679(.O (g5736), .I (I9296));
INVX1 gate1680(.O (g6984), .I (g6382));
INVX1 gate1681(.O (g6280), .I (I10099));
INVX1 gate1682(.O (g6939), .I (I11071));
INVX1 gate1683(.O (g7669), .I (I12286));
INVX1 gate1684(.O (I17246), .I (g11341));
INVX1 gate1685(.O (g11543), .I (g11519));
INVX1 gate1686(.O (g3996), .I (g3144));
INVX1 gate1687(.O (g10184), .I (g10039));
INVX1 gate1688(.O (I12412), .I (g7520));
INVX1 gate1689(.O (I8403), .I (g4264));
INVX1 gate1690(.O (g10674), .I (g10584));
INVX1 gate1691(.O (g8314), .I (I13326));
INVX1 gate1692(.O (g5623), .I (I9053));
INVX1 gate1693(.O (g7772), .I (I12481));
INVX1 gate1694(.O (I7157), .I (g3015));
INVX1 gate1695(.O (g7058), .I (I11255));
INVX1 gate1696(.O (I12133), .I (g6870));
INVX1 gate1697(.O (I5957), .I (g2178));
INVX1 gate1698(.O (I7357), .I (g4077));
INVX1 gate1699(.O (g2122), .I (I5044));
INVX1 gate1700(.O (g2228), .I (g28));
INVX1 gate1701(.O (g7531), .I (I11929));
INVX1 gate1702(.O (g4095), .I (I7233));
INVX1 gate1703(.O (g9554), .I (I14697));
INVX1 gate1704(.O (g8870), .I (I14182));
INVX1 gate1705(.O (g2322), .I (I5378));
INVX1 gate1706(.O (I10927), .I (g6755));
INVX1 gate1707(.O (g7458), .I (g7123));
INVX1 gate1708(.O (g5889), .I (I9514));
INVX1 gate1709(.O (I12229), .I (g7070));
INVX1 gate1710(.O (I6962), .I (g2791));
INVX1 gate1711(.O (g4495), .I (I7886));
INVX1 gate1712(.O (I9839), .I (g5226));
INVX1 gate1713(.O (g2230), .I (g704));
INVX1 gate1714(.O (g4437), .I (g3345));
INVX1 gate1715(.O (g4102), .I (I7244));
INVX1 gate1716(.O (I17591), .I (g11514));
INVX1 gate1717(.O (g4208), .I (I7441));
INVX1 gate1718(.O (g7890), .I (g7479));
INVX1 gate1719(.O (g8650), .I (I13933));
INVX1 gate1720(.O (I13840), .I (g8488));
INVX1 gate1721(.O (I16586), .I (g10850));
INVX1 gate1722(.O (g3379), .I (g3121));
INVX1 gate1723(.O (I15568), .I (g10094));
INVX1 gate1724(.O (g10934), .I (g10827));
INVX1 gate1725(.O (g6106), .I (I9773));
INVX1 gate1726(.O (g5175), .I (g4682));
INVX1 gate1727(.O (g6306), .I (I10177));
INVX1 gate1728(.O (g7505), .I (g7148));
INVX1 gate1729(.O (g3878), .I (g2920));
INVX1 gate1730(.O (g11242), .I (g11112));
INVX1 gate1731(.O (I5098), .I (g38));
INVX1 gate1732(.O (g8008), .I (I12846));
INVX1 gate1733(.O (I10240), .I (g5937));
INVX1 gate1734(.O (g7011), .I (g6503));
INVX1 gate1735(.O (g4719), .I (g3586));
INVX1 gate1736(.O (g10692), .I (I16363));
INVX1 gate1737(.O (g5651), .I (I9114));
INVX1 gate1738(.O (I6587), .I (g2620));
INVX1 gate1739(.O (I10648), .I (g6030));
INVX1 gate1740(.O (I15814), .I (g10202));
INVX1 gate1741(.O (g8336), .I (I13388));
INVX1 gate1742(.O (I14903), .I (g9507));
INVX1 gate1743(.O (I5833), .I (g2103));
INVX1 gate1744(.O (g6387), .I (g6121));
INVX1 gate1745(.O (g5285), .I (g4355));
INVX1 gate1746(.O (g6461), .I (I10391));
INVX1 gate1747(.O (I15807), .I (g10284));
INVX1 gate1748(.O (I15974), .I (g10411));
INVX1 gate1749(.O (I8858), .I (g4506));
INVX1 gate1750(.O (g2550), .I (g1834));
INVX1 gate1751(.O (g7074), .I (I11299));
INVX1 gate1752(.O (I16720), .I (g10854));
INVX1 gate1753(.O (g3271), .I (I6443));
INVX1 gate1754(.O (g10400), .I (g10348));
INVX1 gate1755(.O (g2845), .I (g2168));
INVX1 gate1756(.O (I9282), .I (g5633));
INVX1 gate1757(.O (I15639), .I (g10179));
INVX1 gate1758(.O (I10563), .I (g6043));
INVX1 gate1759(.O (I5584), .I (g1200));
INVX1 gate1760(.O (g10214), .I (I15586));
INVX1 gate1761(.O (g9490), .I (g9324));
INVX1 gate1762(.O (g9823), .I (I14970));
INVX1 gate1763(.O (g2195), .I (g83));
INVX1 gate1764(.O (g4265), .I (g3664));
INVX1 gate1765(.O (I15293), .I (g10001));
INVX1 gate1766(.O (I9988), .I (g5526));
INVX1 gate1767(.O (g6427), .I (I10343));
INVX1 gate1768(.O (I12627), .I (g7697));
INVX1 gate1769(.O (g2395), .I (g231));
INVX1 gate1770(.O (g2891), .I (I6055));
INVX1 gate1771(.O (g5184), .I (g4682));
INVX1 gate1772(.O (g2337), .I (I5395));
INVX1 gate1773(.O (I11483), .I (g6567));
INVX1 gate1774(.O (g2913), .I (I6088));
INVX1 gate1775(.O (g10329), .I (I15775));
INVX1 gate1776(.O (g10207), .I (g10186));
INVX1 gate1777(.O (g4442), .I (g3638));
INVX1 gate1778(.O (I6985), .I (g2890));
INVX1 gate1779(.O (g6904), .I (I11008));
INVX1 gate1780(.O (g6200), .I (I9935));
INVX1 gate1781(.O (g11638), .I (I17724));
INVX1 gate1782(.O (g10539), .I (I16184));
INVX1 gate1783(.O (g4786), .I (I8154));
INVX1 gate1784(.O (g6046), .I (I9669));
INVX1 gate1785(.O (g8065), .I (I12913));
INVX1 gate1786(.O (g3799), .I (I7022));
INVX1 gate1787(.O (I8315), .I (g4788));
INVX1 gate1788(.O (I8811), .I (g4465));
INVX1 gate1789(.O (g6446), .I (I10370));
INVX1 gate1790(.O (g8122), .I (I12981));
INVX1 gate1791(.O (g3981), .I (I7118));
INVX1 gate1792(.O (g8465), .I (g8289));
INVX1 gate1793(.O (g9529), .I (I14672));
INVX1 gate1794(.O (g4164), .I (I7311));
INVX1 gate1795(.O (g10538), .I (I16181));
INVX1 gate1796(.O (g4233), .I (g3698));
INVX1 gate1797(.O (g5424), .I (I8865));
INVX1 gate1798(.O (g9348), .I (I14549));
INVX1 gate1799(.O (I11326), .I (g6660));
INVX1 gate1800(.O (I13949), .I (g8451));
INVX1 gate1801(.O (g6403), .I (g6128));
INVX1 gate1802(.O (I13326), .I (g8203));
INVX1 gate1803(.O (I9804), .I (g5417));
INVX1 gate1804(.O (g6145), .I (I9860));
INVX1 gate1805(.O (g2859), .I (I5995));
INVX1 gate1806(.O (g3997), .I (I7131));
INVX1 gate1807(.O (I15510), .I (g10035));
INVX1 gate1808(.O (g9355), .I (I14570));
INVX1 gate1809(.O (I9792), .I (g5403));
INVX1 gate1810(.O (I6832), .I (g2909));
INVX1 gate1811(.O (g4454), .I (g3914));
INVX1 gate1812(.O (g8033), .I (I12875));
INVX1 gate1813(.O (g11510), .I (I17549));
INVX1 gate1814(.O (g6191), .I (g5446));
INVX1 gate1815(.O (g7569), .I (I12029));
INVX1 gate1816(.O (g5672), .I (I9177));
INVX1 gate1817(.O (g4296), .I (I7559));
INVX1 gate1818(.O (I11904), .I (g6902));
INVX1 gate1819(.O (I10633), .I (g6015));
INVX1 gate1820(.O (I10898), .I (g6735));
INVX1 gate1821(.O (g5231), .I (g4640));
INVX1 gate1822(.O (I17318), .I (g11340));
INVX1 gate1823(.O (g3332), .I (I6513));
INVX1 gate1824(.O (I11252), .I (g6542));
INVX1 gate1825(.O (g10241), .I (g10192));
INVX1 gate1826(.O (g9260), .I (g8892));
INVX1 gate1827(.O (g6695), .I (I10666));
INVX1 gate1828(.O (I10719), .I (g6003));
INVX1 gate1829(.O (I13621), .I (g8315));
INVX1 gate1830(.O (g5643), .I (I9090));
INVX1 gate1831(.O (g3353), .I (g3121));
INVX1 gate1832(.O (I7735), .I (g3759));
INVX1 gate1833(.O (I6507), .I (g2808));
INVX1 gate1834(.O (I14191), .I (g8795));
INVX1 gate1835(.O (g8096), .I (I12953));
INVX1 gate1836(.O (g2248), .I (g99));
INVX1 gate1837(.O (g11578), .I (I17616));
INVX1 gate1838(.O (g2342), .I (I5406));
INVX1 gate1839(.O (I7782), .I (g3775));
INVX1 gate1840(.O (g6107), .I (I9776));
INVX1 gate1841(.O (I17540), .I (g11498));
INVX1 gate1842(.O (I12857), .I (g7638));
INVX1 gate1843(.O (g11014), .I (I16735));
INVX1 gate1844(.O (g6307), .I (I10180));
INVX1 gate1845(.O (g3744), .I (g3307));
INVX1 gate1846(.O (g6536), .I (I10456));
INVX1 gate1847(.O (I4883), .I (g581));
INVX1 gate1848(.O (g5205), .I (g4366));
INVX1 gate1849(.O (I15586), .I (g10159));
INVX1 gate1850(.O (I8880), .I (g4537));
INVX1 gate1851(.O (g2255), .I (I5276));
INVX1 gate1852(.O (I5728), .I (g2084));
INVX1 gate1853(.O (g7688), .I (g7148));
INVX1 gate1854(.O (I12793), .I (g7619));
INVX1 gate1855(.O (g2481), .I (g882));
INVX1 gate1856(.O (I9202), .I (g4915));
INVX1 gate1857(.O (g8195), .I (I13122));
INVX1 gate1858(.O (g7976), .I (I12776));
INVX1 gate1859(.O (g8137), .I (I13010));
INVX1 gate1860(.O (g8891), .I (I14239));
INVX1 gate1861(.O (g8337), .I (I13391));
INVX1 gate1862(.O (g10235), .I (g10189));
INVX1 gate1863(.O (g4012), .I (I7154));
INVX1 gate1864(.O (I11183), .I (g6507));
INVX1 gate1865(.O (I16193), .I (g10485));
INVX1 gate1866(.O (g11442), .I (I17377));
INVX1 gate1867(.O (g2097), .I (I4935));
INVX1 gate1868(.O (I12765), .I (g7638));
INVX1 gate1869(.O (g10683), .I (g10612));
INVX1 gate1870(.O (g5742), .I (I9308));
INVX1 gate1871(.O (g2726), .I (g2021));
INVX1 gate1872(.O (g4412), .I (I7746));
INVX1 gate1873(.O (I11397), .I (g6713));
INVX1 gate1874(.O (I13397), .I (g8138));
INVX1 gate1875(.O (g2154), .I (I5067));
INVX1 gate1876(.O (g6016), .I (I9632));
INVX1 gate1877(.O (I12690), .I (g7555));
INVX1 gate1878(.O (g4189), .I (I7384));
INVX1 gate1879(.O (I5070), .I (g1194));
INVX1 gate1880(.O (g2960), .I (I6173));
INVX1 gate1881(.O (I10861), .I (g6694));
INVX1 gate1882(.O (I10573), .I (g5980));
INVX1 gate1883(.O (I9567), .I (g5556));
INVX1 gate1884(.O (g8807), .I (I14140));
INVX1 gate1885(.O (I14573), .I (g9029));
INVX1 gate1886(.O (g4888), .I (I8237));
INVX1 gate1887(.O (g7126), .I (I11367));
INVX1 gate1888(.O (I13933), .I (g8505));
INVX1 gate1889(.O (I17377), .I (g11412));
INVX1 gate1890(.O (g7326), .I (I11626));
INVX1 gate1891(.O (I10045), .I (g5727));
INVX1 gate1892(.O (g6115), .I (I9798));
INVX1 gate1893(.O (g6251), .I (I10012));
INVX1 gate1894(.O (g4171), .I (I7330));
INVX1 gate1895(.O (g6315), .I (I10204));
INVX1 gate1896(.O (g6811), .I (I10843));
INVX1 gate1897(.O (I15275), .I (g9994));
INVX1 gate1898(.O (g4371), .I (I7674));
INVX1 gate1899(.O (I14045), .I (g8603));
INVX1 gate1900(.O (I17739), .I (g11641));
INVX1 gate1901(.O (g4429), .I (I7779));
INVX1 gate1902(.O (g4787), .I (g3423));
INVX1 gate1903(.O (I8982), .I (g4728));
INVX1 gate1904(.O (g11041), .I (I16784));
INVX1 gate1905(.O (g10882), .I (I16616));
INVX1 gate1906(.O (g5754), .I (I9332));
INVX1 gate1907(.O (I9776), .I (g5353));
INVX1 gate1908(.O (I10099), .I (g5800));
INVX1 gate1909(.O (I16475), .I (g10765));
INVX1 gate1910(.O (g6447), .I (g6166));
INVX1 gate1911(.O (I10388), .I (g5830));
INVX1 gate1912(.O (I8234), .I (g4232));
INVX1 gate1913(.O (g7760), .I (I12445));
INVX1 gate1914(.O (I14388), .I (g8924));
INVX1 gate1915(.O (I8328), .I (g4801));
INVX1 gate1916(.O (I17146), .I (g11305));
INVX1 gate1917(.O (I16863), .I (g10972));
INVX1 gate1918(.O (g3092), .I (g2181));
INVX1 gate1919(.O (I14701), .I (g9291));
INVX1 gate1920(.O (I10251), .I (g6126));
INVX1 gate1921(.O (I14534), .I (g9290));
INVX1 gate1922(.O (g4281), .I (g3586));
INVX1 gate1923(.O (I9965), .I (g5493));
INVX1 gate1924(.O (g5613), .I (g4840));
INVX1 gate1925(.O (g6874), .I (I10958));
INVX1 gate1926(.O (g8142), .I (I13023));
INVX1 gate1927(.O (g2112), .I (g639));
INVX1 gate1928(.O (g8342), .I (I13406));
INVX1 gate1929(.O (g2218), .I (g85));
INVX1 gate1930(.O (I15983), .I (g10414));
INVX1 gate1931(.O (g2267), .I (I5304));
INVX1 gate1932(.O (I17698), .I (g11616));
INVX1 gate1933(.O (g11035), .I (I16766));
INVX1 gate1934(.O (g8255), .I (g7986));
INVX1 gate1935(.O (g8081), .I (g8000));
INVX1 gate1936(.O (g8481), .I (g8324));
INVX1 gate1937(.O (g2001), .I (g814));
INVX1 gate1938(.O (g7608), .I (I12174));
INVX1 gate1939(.O (g7924), .I (g7470));
INVX1 gate1940(.O (I5406), .I (g898));
INVX1 gate1941(.O (g7220), .I (I11456));
INVX1 gate1942(.O (g5572), .I (I8989));
INVX1 gate1943(.O (g5862), .I (I9479));
INVX1 gate1944(.O (I12245), .I (g7093));
INVX1 gate1945(.O (g7779), .I (I12502));
INVX1 gate1946(.O (I4780), .I (g872));
INVX1 gate1947(.O (I6040), .I (g2216));
INVX1 gate1948(.O (g6595), .I (I10563));
INVX1 gate1949(.O (g10584), .I (g10522));
INVX1 gate1950(.O (I15517), .I (g10051));
INVX1 gate1951(.O (I13574), .I (g8360));
INVX1 gate1952(.O (g2329), .I (I5383));
INVX1 gate1953(.O (g8354), .I (I13442));
INVX1 gate1954(.O (I14140), .I (g8717));
INVX1 gate1955(.O (g7023), .I (I11166));
INVX1 gate1956(.O (I7952), .I (g3664));
INVX1 gate1957(.O (g4963), .I (I8337));
INVX1 gate1958(.O (g10206), .I (g10178));
INVX1 gate1959(.O (I5801), .I (g1984));
INVX1 gate1960(.O (I7276), .I (g2861));
INVX1 gate1961(.O (g9670), .I (I14799));
INVX1 gate1962(.O (I16781), .I (g10893));
INVX1 gate1963(.O (g4791), .I (I8161));
INVX1 gate1964(.O (g7977), .I (I12779));
INVX1 gate1965(.O (g2828), .I (I5940));
INVX1 gate1966(.O (g6272), .I (I10075));
INVX1 gate1967(.O (I16236), .I (g10535));
INVX1 gate1968(.O (g3262), .I (I6432));
INVX1 gate1969(.O (g2727), .I (g2022));
INVX1 gate1970(.O (g3736), .I (I6924));
INVX1 gate1971(.O (g5534), .I (g4545));
INVX1 gate1972(.O (g5729), .I (I9279));
INVX1 gate1973(.O (g7361), .I (I11731));
INVX1 gate1974(.O (g10114), .I (I15350));
INVX1 gate1975(.O (I16175), .I (g10488));
INVX1 gate1976(.O (g9813), .I (I14948));
INVX1 gate1977(.O (I15193), .I (g9968));
INVX1 gate1978(.O (g6417), .I (g6136));
INVX1 gate1979(.O (I13051), .I (g8060));
INVX1 gate1980(.O (I15362), .I (g9987));
INVX1 gate1981(.O (g6935), .I (I11065));
INVX1 gate1982(.O (g11193), .I (g11112));
INVX1 gate1983(.O (g7051), .I (I11232));
INVX1 gate1984(.O (g10107), .I (I15341));
INVX1 gate1985(.O (I11756), .I (g7191));
INVX1 gate1986(.O (g2221), .I (I5198));
INVX1 gate1987(.O (g3076), .I (I6282));
INVX1 gate1988(.O (I13592), .I (g8362));
INVX1 gate1989(.O (g8783), .I (g8746));
INVX1 gate1990(.O (I15523), .I (g10058));
INVX1 gate1991(.O (g7327), .I (I11629));
INVX1 gate1992(.O (I12232), .I (g7072));
INVX1 gate1993(.O (I6528), .I (g3274));
INVX1 gate1994(.O (I16264), .I (g10557));
INVX1 gate1995(.O (g8979), .I (I14358));
INVX1 gate1996(.O (I16790), .I (g10900));
INVX1 gate1997(.O (I8490), .I (g4526));
INVX1 gate1998(.O (g4201), .I (I7420));
INVX1 gate1999(.O (I6648), .I (g2635));
INVX1 gate2000(.O (g8218), .I (g7826));
INVX1 gate2001(.O (I9658), .I (g5150));
INVX1 gate2002(.O (g8312), .I (I13320));
INVX1 gate2003(.O (I7546), .I (g4105));
INVX1 gate2004(.O (g6128), .I (I9829));
INVX1 gate2005(.O (g6629), .I (I10584));
INVX1 gate2006(.O (g5885), .I (g5361));
INVX1 gate2007(.O (g10345), .I (I15801));
INVX1 gate2008(.O (g7999), .I (I12825));
INVX1 gate2009(.O (g7146), .I (I11391));
INVX1 gate2010(.O (g5660), .I (I9141));
INVX1 gate2011(.O (I5445), .I (g922));
INVX1 gate2012(.O (g6330), .I (I10221));
INVX1 gate2013(.O (g7346), .I (I11686));
INVX1 gate2014(.O (I10162), .I (g5943));
INVX1 gate2015(.O (g7633), .I (I12239));
INVX1 gate2016(.O (g4049), .I (g3144));
INVX1 gate2017(.O (g3375), .I (I6569));
INVX1 gate2018(.O (g8001), .I (I12829));
INVX1 gate2019(.O (I12261), .I (g7078));
INVX1 gate2020(.O (g4449), .I (g4144));
INVX1 gate2021(.O (g3722), .I (I6894));
INVX1 gate2022(.O (I8456), .I (g4472));
INVX1 gate2023(.O (g7103), .I (I11338));
INVX1 gate2024(.O (g5903), .I (I9536));
INVX1 gate2025(.O (g4575), .I (g3880));
INVX1 gate2026(.O (g10848), .I (I16546));
INVX1 gate2027(.O (g11475), .I (I17466));
INVX1 gate2028(.O (g8293), .I (I13233));
INVX1 gate2029(.O (g8129), .I (g8015));
INVX1 gate2030(.O (I6010), .I (g2256));
INVX1 gate2031(.O (g2068), .I (I4866));
INVX1 gate2032(.O (I11152), .I (g6469));
INVX1 gate2033(.O (g8329), .I (I13367));
INVX1 gate2034(.O (g10141), .I (I15421));
INVX1 gate2035(.O (g7696), .I (g7148));
INVX1 gate2036(.O (g10804), .I (I16514));
INVX1 gate2037(.O (g6800), .I (I10810));
INVX1 gate2038(.O (g4098), .I (I7240));
INVX1 gate2039(.O (g3500), .I (I6690));
INVX1 gate2040(.O (I15437), .I (g10050));
INVX1 gate2041(.O (I16209), .I (g10452));
INVX1 gate2042(.O (I8851), .I (g4498));
INVX1 gate2043(.O (I11731), .I (g7021));
INVX1 gate2044(.O (g8828), .I (g8744));
INVX1 gate2045(.O (g11437), .I (I17362));
INVX1 gate2046(.O (g2677), .I (g2034));
INVX1 gate2047(.O (g10263), .I (g10127));
INVX1 gate2048(.O (g7753), .I (I12424));
INVX1 gate2049(.O (I9981), .I (g5514));
INVX1 gate2050(.O (g8727), .I (g8592));
INVX1 gate2051(.O (g5679), .I (I9194));
INVX1 gate2052(.O (g7508), .I (g6950));
INVX1 gate2053(.O (g3384), .I (g3143));
INVX1 gate2054(.O (g10332), .I (I15782));
INVX1 gate2055(.O (g6213), .I (g5426));
INVX1 gate2056(.O (g8592), .I (I13837));
INVX1 gate2057(.O (g7944), .I (g7410));
INVX1 gate2058(.O (I15347), .I (g9995));
INVX1 gate2059(.O (g7072), .I (I11293));
INVX1 gate2060(.O (I15253), .I (g9987));
INVX1 gate2061(.O (g10135), .I (I15403));
INVX1 gate2062(.O (I12445), .I (g7521));
INVX1 gate2063(.O (g11347), .I (I17164));
INVX1 gate2064(.O (g4896), .I (I8253));
INVX1 gate2065(.O (I7906), .I (g3907));
INVX1 gate2066(.O (g2349), .I (I5421));
INVX1 gate2067(.O (g7043), .I (I11214));
INVX1 gate2068(.O (I12499), .I (g7725));
INVX1 gate2069(.O (I11405), .I (g6627));
INVX1 gate2070(.O (g5288), .I (g4438));
INVX1 gate2071(.O (g9341), .I (I14528));
INVX1 gate2072(.O (g3424), .I (g2896));
INVX1 gate2073(.O (I9132), .I (g4893));
INVX1 gate2074(.O (g10361), .I (g10268));
INVX1 gate2075(.O (g3737), .I (g2834));
INVX1 gate2076(.O (g7443), .I (I11841));
INVX1 gate2077(.O (I9332), .I (g4935));
INVX1 gate2078(.O (g9525), .I (g9257));
INVX1 gate2079(.O (I9153), .I (g5027));
INVX1 gate2080(.O (I9680), .I (g5194));
INVX1 gate2081(.O (I10147), .I (g5697));
INVX1 gate2082(.O (I6343), .I (g1963));
INVX1 gate2083(.O (I10355), .I (g6003));
INVX1 gate2084(.O (g7116), .I (I11351));
INVX1 gate2085(.O (g5805), .I (I9409));
INVX1 gate2086(.O (g5916), .I (I9550));
INVX1 gate2087(.O (g7316), .I (I11596));
INVX1 gate2088(.O (g2198), .I (g668));
INVX1 gate2089(.O (I6282), .I (g2231));
INVX1 gate2090(.O (g4268), .I (I7523));
INVX1 gate2091(.O (I7771), .I (g3418));
INVX1 gate2092(.O (I16607), .I (g10787));
INVX1 gate2093(.O (g2855), .I (I5989));
INVX1 gate2094(.O (g4362), .I (I7651));
INVX1 gate2095(.O (I11929), .I (g6901));
INVX1 gate2096(.O (I14355), .I (g8948));
INVX1 gate2097(.O (I12989), .I (g8043));
INVX1 gate2098(.O (g11351), .I (I17170));
INVX1 gate2099(.O (g3077), .I (g2213));
INVX1 gate2100(.O (g5422), .I (g4470));
INVX1 gate2101(.O (g7034), .I (I11191));
INVX1 gate2102(.O (I10825), .I (g6588));
INVX1 gate2103(.O (g4419), .I (I7763));
INVX1 gate2104(.O (I9744), .I (g5263));
INVX1 gate2105(.O (I12056), .I (g6929));
INVX1 gate2106(.O (I10370), .I (g5857));
INVX1 gate2107(.O (g6166), .I (I9893));
INVX1 gate2108(.O (g8624), .I (g8486));
INVX1 gate2109(.O (g3523), .I (g2971));
INVX1 gate2110(.O (I14370), .I (g8954));
INVX1 gate2111(.O (g8953), .I (I14312));
INVX1 gate2112(.O (I10858), .I (g6688));
INVX1 gate2113(.O (I13020), .I (g8049));
INVX1 gate2114(.O (I13583), .I (g8344));
INVX1 gate2115(.O (g4452), .I (g3365));
INVX1 gate2116(.O (I8872), .I (g4529));
INVX1 gate2117(.O (I15063), .I (g9699));
INVX1 gate2118(.O (g2241), .I (g722));
INVX1 gate2119(.O (g7147), .I (I11394));
INVX1 gate2120(.O (g6056), .I (g5426));
INVX1 gate2121(.O (g5947), .I (I9585));
INVX1 gate2122(.O (g7347), .I (I11689));
INVX1 gate2123(.O (g11063), .I (g10974));
INVX1 gate2124(.O (I11046), .I (g6635));
INVX1 gate2125(.O (I10996), .I (g6786));
INVX1 gate2126(.O (I12271), .I (g7218));
INVX1 gate2127(.O (g7681), .I (g7148));
INVX1 gate2128(.O (g6649), .I (I10610));
INVX1 gate2129(.O (I8989), .I (g4746));
INVX1 gate2130(.O (g8677), .I (I13962));
INVX1 gate2131(.O (g110), .I (I4786));
INVX1 gate2132(.O (I10367), .I (g6234));
INVX1 gate2133(.O (I10394), .I (g5824));
INVX1 gate2134(.O (I9901), .I (g5557));
INVX1 gate2135(.O (g7697), .I (g7101));
INVX1 gate2136(.O (I14367), .I (g8953));
INVX1 gate2137(.O (I14394), .I (g8884));
INVX1 gate2138(.O (I16641), .I (g10864));
INVX1 gate2139(.O (g3742), .I (I6929));
INVX1 gate2140(.O (g7914), .I (g7651));
INVX1 gate2141(.O (g8576), .I (I13819));
INVX1 gate2142(.O (g2524), .I (g986));
INVX1 gate2143(.O (g7210), .I (I11440));
INVX1 gate2144(.O (g4728), .I (I8080));
INVX1 gate2145(.O (I16292), .I (g10551));
INVX1 gate2146(.O (g2644), .I (g1990));
INVX1 gate2147(.O (g6698), .I (I10671));
INVX1 gate2148(.O (g4730), .I (g3546));
INVX1 gate2149(.O (g8716), .I (g8576));
INVX1 gate2150(.O (I17546), .I (g11500));
INVX1 gate2151(.O (g8149), .I (I13036));
INVX1 gate2152(.O (g10947), .I (I16708));
INVX1 gate2153(.O (g4504), .I (I7899));
INVX1 gate2154(.O (I11357), .I (g6594));
INVX1 gate2155(.O (g6964), .I (g6509));
INVX1 gate2156(.O (g8349), .I (I13427));
INVX1 gate2157(.O (g2119), .I (I5031));
INVX1 gate2158(.O (g5095), .I (I8465));
INVX1 gate2159(.O (g6260), .I (I10039));
INVX1 gate2160(.O (g5037), .I (I8414));
INVX1 gate2161(.O (I13357), .I (g8125));
INVX1 gate2162(.O (I12199), .I (g7278));
INVX1 gate2163(.O (g4185), .I (I7372));
INVX1 gate2164(.O (I7244), .I (g3226));
INVX1 gate2165(.O (g9311), .I (I14506));
INVX1 gate2166(.O (g11422), .I (I17321));
INVX1 gate2167(.O (I11743), .I (g7035));
INVX1 gate2168(.O (I13105), .I (g7929));
INVX1 gate2169(.O (g5653), .I (I9120));
INVX1 gate2170(.O (g4385), .I (I7710));
INVX1 gate2171(.O (g7413), .I (g7197));
INVX1 gate2172(.O (g5102), .I (I8476));
INVX1 gate2173(.O (g2258), .I (I5289));
INVX1 gate2174(.O (I14319), .I (g8816));
INVX1 gate2175(.O (g2352), .I (I5430));
INVX1 gate2176(.O (g2818), .I (I5922));
INVX1 gate2177(.O (I7140), .I (g2641));
INVX1 gate2178(.O (g6063), .I (g5446));
INVX1 gate2179(.O (I12529), .I (g7589));
INVX1 gate2180(.O (I5940), .I (g2175));
INVX1 gate2181(.O (g2867), .I (I6007));
INVX1 gate2182(.O (I16635), .I (g10862));
INVX1 gate2183(.O (g10463), .I (I15980));
INVX1 gate2184(.O (g11208), .I (g11077));
INVX1 gate2185(.O (g4470), .I (I7843));
INVX1 gate2186(.O (g8198), .I (I13131));
INVX1 gate2187(.O (g4897), .I (I8256));
INVX1 gate2188(.O (g8747), .I (I14040));
INVX1 gate2189(.O (I7478), .I (g3566));
INVX1 gate2190(.O (g5719), .I (I9259));
INVX1 gate2191(.O (g4425), .I (I7771));
INVX1 gate2192(.O (I12843), .I (g7683));
INVX1 gate2193(.O (I15542), .I (g10065));
INVX1 gate2194(.O (g10972), .I (I16717));
INVX1 gate2195(.O (g10033), .I (I15235));
INVX1 gate2196(.O (I5388), .I (g889));
INVX1 gate2197(.O (g10234), .I (g10188));
INVX1 gate2198(.O (I7435), .I (g3459));
INVX1 gate2199(.O (g7936), .I (g7712));
INVX1 gate2200(.O (g11542), .I (g11519));
INVX1 gate2201(.O (g11453), .I (I17416));
INVX1 gate2202(.O (g5752), .I (I9326));
INVX1 gate2203(.O (I6094), .I (g2110));
INVX1 gate2204(.O (I13803), .I (g8476));
INVX1 gate2205(.O (g3044), .I (I6256));
INVX1 gate2206(.O (g2211), .I (g153));
INVX1 gate2207(.O (I14540), .I (g9310));
INVX1 gate2208(.O (g6279), .I (I10096));
INVX1 gate2209(.O (g2186), .I (g90));
INVX1 gate2210(.O (g7317), .I (I11599));
INVX1 gate2211(.O (g6720), .I (I10713));
INVX1 gate2212(.O (I8253), .I (g4637));
INVX1 gate2213(.O (g6118), .I (I9807));
INVX1 gate2214(.O (g3983), .I (g3222));
INVX1 gate2215(.O (g11614), .I (I17662));
INVX1 gate2216(.O (g7601), .I (I12153));
INVX1 gate2217(.O (I5430), .I (g916));
INVX1 gate2218(.O (g5265), .I (g4362));
INVX1 gate2219(.O (g11436), .I (I17359));
INVX1 gate2220(.O (g3862), .I (g2920));
INVX1 gate2221(.O (g5042), .I (g4840));
INVX1 gate2222(.O (I15320), .I (g10013));
INVX1 gate2223(.O (g9832), .I (I14989));
INVX1 gate2224(.O (g6652), .I (I10613));
INVX1 gate2225(.O (g4678), .I (g3546));
INVX1 gate2226(.O (g6057), .I (g5446));
INVX1 gate2227(.O (g6843), .I (I10901));
INVX1 gate2228(.O (I15530), .I (g10107));
INVX1 gate2229(.O (g11073), .I (g10913));
INVX1 gate2230(.O (g4331), .I (I7606));
INVX1 gate2231(.O (g3543), .I (g3101));
INVX1 gate2232(.O (g2170), .I (g30));
INVX1 gate2233(.O (g2614), .I (g1994));
INVX1 gate2234(.O (g7775), .I (I12490));
INVX1 gate2235(.O (g11593), .I (I17633));
INVX1 gate2236(.O (g7922), .I (I12712));
INVX1 gate2237(.O (g2125), .I (I5053));
INVX1 gate2238(.O (g8319), .I (I13341));
INVX1 gate2239(.O (g11346), .I (I17161));
INVX1 gate2240(.O (I15565), .I (g10101));
INVX1 gate2241(.O (g2821), .I (I5929));
INVX1 gate2242(.O (g9507), .I (g9268));
INVX1 gate2243(.O (I15464), .I (g10094));
INVX1 gate2244(.O (I6965), .I (g2880));
INVX1 gate2245(.O (I10120), .I (g6248));
INVX1 gate2246(.O (g4766), .I (g3440));
INVX1 gate2247(.O (I11662), .I (g7033));
INVX1 gate2248(.O (I10739), .I (g5942));
INVX1 gate2249(.O (g4087), .I (I7220));
INVX1 gate2250(.O (g4105), .I (I7249));
INVX1 gate2251(.O (g8152), .I (I13043));
INVX1 gate2252(.O (g10421), .I (g10331));
INVX1 gate2253(.O (I16537), .I (g10721));
INVX1 gate2254(.O (g8352), .I (I13436));
INVX1 gate2255(.O (g4305), .I (g4013));
INVX1 gate2256(.O (g6971), .I (g6517));
INVX1 gate2257(.O (I13027), .I (g8051));
INVX1 gate2258(.O (I12258), .I (g7103));
INVX1 gate2259(.O (g3729), .I (I6907));
INVX1 gate2260(.O (I6264), .I (g2118));
INVX1 gate2261(.O (I16108), .I (g10383));
INVX1 gate2262(.O (g6686), .I (I10651));
INVX1 gate2263(.O (g10163), .I (I15485));
INVX1 gate2264(.O (g8717), .I (I14010));
INVX1 gate2265(.O (g11034), .I (I16763));
INVX1 gate2266(.O (g7460), .I (g7148));
INVX1 gate2267(.O (g7597), .I (I12133));
INVX1 gate2268(.O (g5296), .I (g4444));
INVX1 gate2269(.O (I11249), .I (g6541));
INVX1 gate2270(.O (I5638), .I (g936));
INVX1 gate2271(.O (I14645), .I (g9088));
INVX1 gate2272(.O (I16283), .I (g10538));
INVX1 gate2273(.O (g2083), .I (g139));
INVX1 gate2274(.O (I6360), .I (g2261));
INVX1 gate2275(.O (g4748), .I (g3546));
INVX1 gate2276(.O (I16492), .I (g10773));
INVX1 gate2277(.O (I13482), .I (g8193));
INVX1 gate2278(.O (I5308), .I (g97));
INVX1 gate2279(.O (I11710), .I (g7020));
INVX1 gate2280(.O (g7784), .I (I12517));
INVX1 gate2281(.O (I4992), .I (g1170));
INVX1 gate2282(.O (g4755), .I (g3440));
INVX1 gate2283(.O (g10541), .I (I16190));
INVX1 gate2284(.O (I10698), .I (g5856));
INVX1 gate2285(.O (g6121), .I (I9816));
INVX1 gate2286(.O (I15409), .I (g10065));
INVX1 gate2287(.O (I7002), .I (g2907));
INVX1 gate2288(.O (g8186), .I (I13109));
INVX1 gate2289(.O (g10473), .I (g10380));
INVX1 gate2290(.O (g4226), .I (g3698));
INVX1 gate2291(.O (I11204), .I (g6523));
INVX1 gate2292(.O (g6670), .I (I10633));
INVX1 gate2293(.O (I7402), .I (g4121));
INVX1 gate2294(.O (g11409), .I (I17268));
INVX1 gate2295(.O (I6996), .I (g2904));
INVX1 gate2296(.O (g3946), .I (I7099));
INVX1 gate2297(.O (I13779), .I (g8514));
INVX1 gate2298(.O (I7236), .I (g3219));
INVX1 gate2299(.O (I15635), .I (g10185));
INVX1 gate2300(.O (I16982), .I (g11088));
INVX1 gate2301(.O (g8599), .I (g8546));
INVX1 gate2302(.O (g7995), .I (I12817));
INVX1 gate2303(.O (g2790), .I (g2276));
INVX1 gate2304(.O (g11408), .I (I17265));
INVX1 gate2305(.O (g7079), .I (I11312));
INVX1 gate2306(.O (g11635), .I (I17719));
INVX1 gate2307(.O (I11778), .I (g7210));
INVX1 gate2308(.O (g3903), .I (I7070));
INVX1 gate2309(.O (g5012), .I (I8388));
INVX1 gate2310(.O (g9100), .I (g8892));
INVX1 gate2311(.O (g8274), .I (I13194));
INVX1 gate2312(.O (I10427), .I (g5839));
INVX1 gate2313(.O (g7479), .I (I11873));
INVX1 gate2314(.O (g8426), .I (I13592));
INVX1 gate2315(.O (g1994), .I (g794));
INVX1 gate2316(.O (g4445), .I (I7803));
INVX1 gate2317(.O (g6253), .I (I10018));
INVX1 gate2318(.O (g2061), .I (g1828));
INVX1 gate2319(.O (g2187), .I (g746));
INVX1 gate2320(.O (g6938), .I (I11068));
INVX1 gate2321(.O (g4173), .I (I7336));
INVX1 gate2322(.O (g6813), .I (I10849));
INVX1 gate2323(.O (g4373), .I (I7680));
INVX1 gate2324(.O (I11786), .I (g7246));
INVX1 gate2325(.O (I16796), .I (g11016));
INVX1 gate2326(.O (g10535), .I (I16172));
INVX1 gate2327(.O (g4491), .I (g3546));
INVX1 gate2328(.O (g8125), .I (I12986));
INVX1 gate2329(.O (g7190), .I (I11412));
INVX1 gate2330(.O (g8325), .I (I13357));
INVX1 gate2331(.O (I11647), .I (g6925));
INVX1 gate2332(.O (g7390), .I (g6847));
INVX1 gate2333(.O (I12878), .I (g7638));
INVX1 gate2334(.O (g5888), .I (g5102));
INVX1 gate2335(.O (I13945), .I (g8488));
INVX1 gate2336(.O (I12171), .I (g6885));
INVX1 gate2337(.O (g10121), .I (I15371));
INVX1 gate2338(.O (g8984), .I (I14373));
INVX1 gate2339(.O (g3436), .I (g3144));
INVX1 gate2340(.O (g4369), .I (I7668));
INVX1 gate2341(.O (g8280), .I (I13212));
INVX1 gate2342(.O (I7556), .I (g4080));
INVX1 gate2343(.O (g4602), .I (I8011));
INVX1 gate2344(.O (g7501), .I (I11879));
INVX1 gate2345(.O (I17450), .I (g11450));
INVX1 gate2346(.O (g3378), .I (I6572));
INVX1 gate2347(.O (g5787), .I (I9383));
INVX1 gate2348(.O (I9424), .I (g4963));
INVX1 gate2349(.O (I9795), .I (g5404));
INVX1 gate2350(.O (I17315), .I (g11393));
INVX1 gate2351(.O (g10344), .I (I15798));
INVX1 gate2352(.O (I9737), .I (g5258));
INVX1 gate2353(.O (g2904), .I (I6065));
INVX1 gate2354(.O (g2200), .I (g92));
INVX1 gate2355(.O (g6552), .I (g5733));
INVX1 gate2356(.O (g7356), .I (I11716));
INVX1 gate2357(.O (g2046), .I (g1845));
INVX1 gate2358(.O (I17707), .I (g11619));
INVX1 gate2359(.O (g4920), .I (I8293));
INVX1 gate2360(.O (I5827), .I (g2271));
INVX1 gate2361(.O (g2446), .I (g1400));
INVX1 gate2362(.O (g4459), .I (I7820));
INVX1 gate2363(.O (I17202), .I (g11322));
INVX1 gate2364(.O (g3335), .I (I6520));
INVX1 gate2365(.O (I13233), .I (g8265));
INVX1 gate2366(.O (g8483), .I (g8332));
INVX1 gate2367(.O (g4767), .I (I8123));
INVX1 gate2368(.O (I7064), .I (g2984));
INVX1 gate2369(.O (g11575), .I (g11561));
INVX1 gate2370(.O (g2003), .I (g822));
INVX1 gate2371(.O (g5281), .I (g4428));
INVX1 gate2372(.O (g3382), .I (I6580));
INVX1 gate2373(.O (I9077), .I (g4765));
INVX1 gate2374(.O (I7899), .I (g3380));
INVX1 gate2375(.O (g4535), .I (g3946));
INVX1 gate2376(.O (I8358), .I (g4794));
INVX1 gate2377(.O (I6611), .I (g2626));
INVX1 gate2378(.O (I8506), .I (g4334));
INVX1 gate2379(.O (g2345), .I (g1936));
INVX1 gate2380(.O (g10173), .I (g10120));
INVX1 gate2381(.O (I17070), .I (g11233));
INVX1 gate2382(.O (g8106), .I (g7950));
INVX1 gate2383(.O (g11109), .I (g10974));
INVX1 gate2384(.O (g8306), .I (I13290));
INVX1 gate2385(.O (g2763), .I (I5847));
INVX1 gate2386(.O (g2191), .I (g1696));
INVX1 gate2387(.O (g2391), .I (I5478));
INVX1 gate2388(.O (g6586), .I (g5949));
INVX1 gate2389(.O (I12919), .I (g8003));
INVX1 gate2390(.O (I6799), .I (g2750));
INVX1 gate2391(.O (I11932), .I (g6908));
INVX1 gate2392(.O (g3749), .I (I6938));
INVX1 gate2393(.O (g8790), .I (I14101));
INVX1 gate2394(.O (I9205), .I (g5309));
INVX1 gate2395(.O (g11108), .I (g10974));
INVX1 gate2396(.O (g2695), .I (g2039));
INVX1 gate2397(.O (g9666), .I (I14793));
INVX1 gate2398(.O (g8061), .I (I12901));
INVX1 gate2399(.O (g5684), .I (I9205));
INVX1 gate2400(.O (I8275), .I (g4351));
INVX1 gate2401(.O (I8311), .I (g4794));
INVX1 gate2402(.O (g4415), .I (g3914));
INVX1 gate2403(.O (g5639), .I (I9080));
INVX1 gate2404(.O (I14127), .I (g8768));
INVX1 gate2405(.O (I17384), .I (g11437));
INVX1 gate2406(.O (g7810), .I (I12595));
INVX1 gate2407(.O (g7363), .I (I11737));
INVX1 gate2408(.O (g10134), .I (I15400));
INVX1 gate2409(.O (I7295), .I (g3260));
INVX1 gate2410(.O (I11961), .I (g7053));
INVX1 gate2411(.O (I16553), .I (g10754));
INVX1 gate2412(.O (g5109), .I (I8495));
INVX1 gate2413(.O (g5791), .I (I9391));
INVX1 gate2414(.O (g3798), .I (g3228));
INVX1 gate2415(.O (I13448), .I (g8150));
INVX1 gate2416(.O (I9099), .I (g5572));
INVX1 gate2417(.O (g2159), .I (I5080));
INVX1 gate2418(.O (g7432), .I (I11824));
INVX1 gate2419(.O (I14490), .I (g8885));
INVX1 gate2420(.O (g6141), .I (I9854));
INVX1 gate2421(.O (g8622), .I (g8485));
INVX1 gate2422(.O (g6570), .I (g5949));
INVX1 gate2423(.O (g6860), .I (g6475));
INVX1 gate2424(.O (g7053), .I (I11238));
INVX1 gate2425(.O (I11505), .I (g6585));
INVX1 gate2426(.O (g9351), .I (I14558));
INVX1 gate2427(.O (I5662), .I (g563));
INVX1 gate2428(.O (g9875), .I (I15036));
INVX1 gate2429(.O (g8427), .I (I13595));
INVX1 gate2430(.O (I5067), .I (g33));
INVX1 gate2431(.O (g9530), .I (I14675));
INVX1 gate2432(.O (g6710), .I (I10693));
INVX1 gate2433(.O (g5808), .I (g5320));
INVX1 gate2434(.O (I5418), .I (g907));
INVX1 gate2435(.O (g2858), .I (I5992));
INVX1 gate2436(.O (I12598), .I (g7628));
INVX1 gate2437(.O (I7194), .I (g2629));
INVX1 gate2438(.O (I14376), .I (g8959));
INVX1 gate2439(.O (I14385), .I (g8890));
INVX1 gate2440(.O (g4203), .I (I7426));
INVX1 gate2441(.O (I8985), .I (g4733));
INVX1 gate2442(.O (I13717), .I (g8354));
INVX1 gate2443(.O (g11381), .I (I17206));
INVX1 gate2444(.O (g4721), .I (g3546));
INVX1 gate2445(.O (g2016), .I (g1361));
INVX1 gate2446(.O (I13212), .I (g8195));
INVX1 gate2447(.O (g2757), .I (I5837));
INVX1 gate2448(.O (g8446), .I (I13636));
INVX1 gate2449(.O (g7568), .I (I12026));
INVX1 gate2450(.O (g5759), .I (I9341));
INVX1 gate2451(.O (I9754), .I (g5271));
INVX1 gate2452(.O (I10888), .I (g6333));
INVX1 gate2453(.O (g8514), .I (I13711));
INVX1 gate2454(.O (I6802), .I (g2751));
INVX1 gate2455(.O (g3632), .I (I6799));
INVX1 gate2456(.O (g3095), .I (g2482));
INVX1 gate2457(.O (g3037), .I (g2135));
INVX1 gate2458(.O (g8003), .I (I12835));
INVX1 gate2459(.O (I14888), .I (g9454));
INVX1 gate2460(.O (I16252), .I (g10515));
INVX1 gate2461(.O (g3437), .I (I6654));
INVX1 gate2462(.O (I12817), .I (g7692));
INVX1 gate2463(.O (I9273), .I (g5091));
INVX1 gate2464(.O (I10671), .I (g6045));
INVX1 gate2465(.O (I17695), .I (g11614));
INVX1 gate2466(.O (g3102), .I (g2482));
INVX1 gate2467(.O (I4924), .I (g123));
INVX1 gate2468(.O (g3208), .I (I6381));
INVX1 gate2469(.O (I12322), .I (g7246));
INVX1 gate2470(.O (g7912), .I (g7651));
INVX1 gate2471(.O (g8145), .I (I13030));
INVX1 gate2472(.O (g8345), .I (I13415));
INVX1 gate2473(.O (g2251), .I (g731));
INVX1 gate2474(.O (g2642), .I (g1988));
INVX1 gate2475(.O (I12159), .I (g7243));
INVX1 gate2476(.O (g7357), .I (I11719));
INVX1 gate2477(.O (g2047), .I (g1857));
INVX1 gate2478(.O (I12532), .I (g7594));
INVX1 gate2479(.O (I12901), .I (g7984));
INVX1 gate2480(.O (g8191), .I (I13114));
INVX1 gate2481(.O (g10927), .I (g10827));
INVX1 gate2482(.O (g9884), .I (I15063));
INVX1 gate2483(.O (g6158), .I (I9883));
INVX1 gate2484(.O (g3719), .I (g2920));
INVX1 gate2485(.O (I12783), .I (g7590));
INVX1 gate2486(.O (g11390), .I (I17219));
INVX1 gate2487(.O (I13723), .I (g8359));
INVX1 gate2488(.O (g5865), .I (I9486));
INVX1 gate2489(.O (g8695), .I (I13978));
INVX1 gate2490(.O (I5847), .I (g2275));
INVX1 gate2491(.O (I6901), .I (g2818));
INVX1 gate2492(.O (I11149), .I (g6468));
INVX1 gate2493(.O (g2874), .I (I6022));
INVX1 gate2494(.O (g7929), .I (g7519));
INVX1 gate2495(.O (g3752), .I (I6947));
INVX1 gate2496(.O (I16673), .I (g10782));
INVX1 gate2497(.O (I11433), .I (g6424));
INVX1 gate2498(.O (I16847), .I (g10886));
INVX1 gate2499(.O (I11387), .I (g6672));
INVX1 gate2500(.O (g5604), .I (I9032));
INVX1 gate2501(.O (I13433), .I (g8181));
INVX1 gate2502(.O (g5098), .I (g4840));
INVX1 gate2503(.O (g2654), .I (g2012));
INVX1 gate2504(.O (I11620), .I (g6840));
INVX1 gate2505(.O (g4188), .I (I7381));
INVX1 gate2506(.O (g5498), .I (I8919));
INVX1 gate2507(.O (I9712), .I (g5230));
INVX1 gate2508(.O (g6587), .I (g5827));
INVX1 gate2509(.O (g4388), .I (I7719));
INVX1 gate2510(.O (g10491), .I (I16108));
INVX1 gate2511(.O (g10903), .I (g10809));
INVX1 gate2512(.O (I11097), .I (g6748));
INVX1 gate2513(.O (I5421), .I (g549));
INVX1 gate2514(.O (g8359), .I (I13457));
INVX1 gate2515(.O (g6111), .I (I9786));
INVX1 gate2516(.O (g6275), .I (I10084));
INVX1 gate2517(.O (g6311), .I (I10192));
INVX1 gate2518(.O (g4216), .I (I7465));
INVX1 gate2519(.O (g10604), .I (I16280));
INVX1 gate2520(.O (g9343), .I (I14534));
INVX1 gate2521(.O (g8858), .I (g8743));
INVX1 gate2522(.O (g4671), .I (g3354));
INVX1 gate2523(.O (g2880), .I (I6028));
INVX1 gate2524(.O (g4428), .I (I7776));
INVX1 gate2525(.O (g2537), .I (I5646));
INVX1 gate2526(.O (I10546), .I (g5914));
INVX1 gate2527(.O (g5896), .I (I9525));
INVX1 gate2528(.O (g4430), .I (I7782));
INVX1 gate2529(.O (I14546), .I (g9312));
INVX1 gate2530(.O (I7438), .I (g3461));
INVX1 gate2531(.O (g3164), .I (I6370));
INVX1 gate2532(.O (g3364), .I (g3121));
INVX1 gate2533(.O (I7009), .I (g2913));
INVX1 gate2534(.O (I10024), .I (g5700));
INVX1 gate2535(.O (I8204), .I (g3976));
INVX1 gate2536(.O (I12631), .I (g7705));
INVX1 gate2537(.O (g8115), .I (g7953));
INVX1 gate2538(.O (g4564), .I (g3880));
INVX1 gate2539(.O (g8251), .I (I13166));
INVX1 gate2540(.O (g8315), .I (I13329));
INVX1 gate2541(.O (g2612), .I (I5737));
INVX1 gate2542(.O (I15326), .I (g10025));
INVX1 gate2543(.O (g2017), .I (g1218));
INVX1 gate2544(.O (g6284), .I (I10111));
INVX1 gate2545(.O (g2243), .I (I5248));
INVX1 gate2546(.O (g8447), .I (I13639));
INVX1 gate2547(.O (I6580), .I (g3186));
INVX1 gate2548(.O (g3770), .I (I6985));
INVX1 gate2549(.O (g6239), .I (I9988));
INVX1 gate2550(.O (g10794), .I (I16496));
INVX1 gate2551(.O (I15536), .I (g10111));
INVX1 gate2552(.O (g10395), .I (g10320));
INVX1 gate2553(.O (g5419), .I (I8858));
INVX1 gate2554(.O (g9804), .I (I14939));
INVX1 gate2555(.O (g10262), .I (g10142));
INVX1 gate2556(.O (g7683), .I (g7148));
INVX1 gate2557(.O (g11040), .I (I16781));
INVX1 gate2558(.O (g10899), .I (g10803));
INVX1 gate2559(.O (g6591), .I (I10553));
INVX1 gate2560(.O (I11412), .I (g6411));
INVX1 gate2561(.O (g5052), .I (g4394));
INVX1 gate2562(.O (I13412), .I (g8142));
INVX1 gate2563(.O (I5101), .I (g1960));
INVX1 gate2564(.O (g8874), .I (I14194));
INVX1 gate2565(.O (g3532), .I (g3164));
INVX1 gate2566(.O (g7778), .I (I12499));
INVX1 gate2567(.O (g2234), .I (g87));
INVX1 gate2568(.O (g6853), .I (I10917));
INVX1 gate2569(.O (I10126), .I (g5682));
INVX1 gate2570(.O (I10659), .I (g6038));
INVX1 gate2571(.O (I16574), .I (g10821));
INVX1 gate2572(.O (g2629), .I (g2001));
INVX1 gate2573(.O (g4638), .I (g3354));
INVX1 gate2574(.O (g2328), .I (g1882));
INVX1 gate2575(.O (I12289), .I (g7142));
INVX1 gate2576(.O (I6968), .I (g2881));
INVX1 gate2577(.O (g6420), .I (I10334));
INVX1 gate2578(.O (g11621), .I (I17681));
INVX1 gate2579(.O (g2130), .I (I5057));
INVX1 gate2580(.O (g10191), .I (I15551));
INVX1 gate2581(.O (g2542), .I (g1868));
INVX1 gate2582(.O (I8973), .I (g4488));
INVX1 gate2583(.O (g2330), .I (g1891));
INVX1 gate2584(.O (g7735), .I (I12384));
INVX1 gate2585(.O (I16311), .I (g10584));
INVX1 gate2586(.O (g4308), .I (g3863));
INVX1 gate2587(.O (I11228), .I (g6471));
INVX1 gate2588(.O (I17231), .I (g11303));
INVX1 gate2589(.O (g7782), .I (I12511));
INVX1 gate2590(.O (g6559), .I (g5758));
INVX1 gate2591(.O (I12571), .I (g7509));
INVX1 gate2592(.O (g3012), .I (I6247));
INVX1 gate2593(.O (I11011), .I (g6340));
INVX1 gate2594(.O (I5751), .I (g2296));
INVX1 gate2595(.O (g8595), .I (I13840));
INVX1 gate2596(.O (g6931), .I (I11055));
INVX1 gate2597(.O (g5728), .I (I9276));
INVX1 gate2598(.O (g5486), .I (g4395));
INVX1 gate2599(.O (I10296), .I (g6242));
INVX1 gate2600(.O (I11716), .I (g7026));
INVX1 gate2601(.O (g5730), .I (I9282));
INVX1 gate2602(.O (g5504), .I (g4419));
INVX1 gate2603(.O (g7949), .I (g7422));
INVX1 gate2604(.O (g4217), .I (I7468));
INVX1 gate2605(.O (g11183), .I (I16950));
INVX1 gate2606(.O (I8123), .I (g3630));
INVX1 gate2607(.O (g3990), .I (g3121));
INVX1 gate2608(.O (g2554), .I (I5672));
INVX1 gate2609(.O (g4758), .I (g3586));
INVX1 gate2610(.O (g4066), .I (I7191));
INVX1 gate2611(.O (g8272), .I (I13188));
INVX1 gate2612(.O (I16592), .I (g10781));
INVX1 gate2613(.O (g4589), .I (I7996));
INVX1 gate2614(.O (g5185), .I (g4682));
INVX1 gate2615(.O (g11397), .I (I17234));
INVX1 gate2616(.O (g5881), .I (g5361));
INVX1 gate2617(.O (g7627), .I (I12223));
INVX1 gate2618(.O (g9094), .I (g8892));
INVX1 gate2619(.O (I5041), .I (g1179));
INVX1 gate2620(.O (I9135), .I (g5198));
INVX1 gate2621(.O (g4466), .I (I7833));
INVX1 gate2622(.O (g1992), .I (g782));
INVX1 gate2623(.O (g6905), .I (I11011));
INVX1 gate2624(.O (g8978), .I (I14355));
INVX1 gate2625(.O (I5441), .I (g919));
INVX1 gate2626(.O (g3371), .I (g2837));
INVX1 gate2627(.O (g11062), .I (g10937));
INVX1 gate2628(.O (I10060), .I (g5752));
INVX1 gate2629(.O (g2213), .I (g1110));
INVX1 gate2630(.O (g11509), .I (I17546));
INVX1 gate2631(.O (g7998), .I (I12822));
INVX1 gate2632(.O (g10247), .I (I15639));
INVX1 gate2633(.O (g4165), .I (g3164));
INVX1 gate2634(.O (g4365), .I (g3880));
INVX1 gate2635(.O (I13627), .I (g8326));
INVX1 gate2636(.O (g5425), .I (g4300));
INVX1 gate2637(.O (g10389), .I (g10307));
INVX1 gate2638(.O (g10926), .I (g10827));
INVX1 gate2639(.O (I10855), .I (g6685));
INVX1 gate2640(.O (I13959), .I (g8451));
INVX1 gate2641(.O (I13379), .I (g8133));
INVX1 gate2642(.O (g11508), .I (I17543));
INVX1 gate2643(.O (g4711), .I (I8061));
INVX1 gate2644(.O (g6100), .I (I9759));
INVX1 gate2645(.O (I11112), .I (g6445));
INVX1 gate2646(.O (g8982), .I (I14367));
INVX1 gate2647(.O (g11634), .I (I17716));
INVX1 gate2648(.O (g10612), .I (I16286));
INVX1 gate2649(.O (g6300), .I (I10159));
INVX1 gate2650(.O (g7603), .I (I12159));
INVX1 gate2651(.O (g4055), .I (g3144));
INVX1 gate2652(.O (g7039), .I (I11204));
INVX1 gate2653(.O (I9749), .I (g5266));
INVX1 gate2654(.O (g10388), .I (g10305));
INVX1 gate2655(.O (I8351), .I (g4794));
INVX1 gate2656(.O (g8234), .I (g7826));
INVX1 gate2657(.O (g2902), .I (I6061));
INVX1 gate2658(.O (g7439), .I (I11833));
INVX1 gate2659(.O (g8128), .I (I12993));
INVX1 gate2660(.O (g8328), .I (I13364));
INVX1 gate2661(.O (g7850), .I (I12647));
INVX1 gate2662(.O (g10534), .I (I16169));
INVX1 gate2663(.O (g10098), .I (I15332));
INVX1 gate2664(.O (I17456), .I (g11453));
INVX1 gate2665(.O (g4333), .I (g4144));
INVX1 gate2666(.O (I7837), .I (g4158));
INVX1 gate2667(.O (g8330), .I (I13370));
INVX1 gate2668(.O (g10251), .I (g10195));
INVX1 gate2669(.O (g10272), .I (g10168));
INVX1 gate2670(.O (g2090), .I (I4920));
INVX1 gate2671(.O (g4774), .I (I8136));
INVX1 gate2672(.O (I7462), .I (g3721));
INVX1 gate2673(.O (I9798), .I (g5415));
INVX1 gate2674(.O (I13096), .I (g7925));
INVX1 gate2675(.O (g2166), .I (I5101));
INVX1 gate2676(.O (g6750), .I (I10759));
INVX1 gate2677(.O (g9264), .I (I14477));
INVX1 gate2678(.O (I6424), .I (g2462));
INVX1 gate2679(.O (g7702), .I (g7079));
INVX1 gate2680(.O (g4196), .I (I7405));
INVX1 gate2681(.O (g5678), .I (I9191));
INVX1 gate2682(.O (I10503), .I (g5858));
INVX1 gate2683(.O (I16413), .I (g10663));
INVX1 gate2684(.O (g10462), .I (I15977));
INVX1 gate2685(.O (g4396), .I (I7735));
INVX1 gate2686(.O (g3138), .I (I6356));
INVX1 gate2687(.O (g8800), .I (I14123));
INVX1 gate2688(.O (I14503), .I (g8920));
INVX1 gate2689(.O (I8410), .I (g4283));
INVX1 gate2690(.O (g2056), .I (I4859));
INVX1 gate2691(.O (I16691), .I (g10788));
INVX1 gate2692(.O (g9360), .I (I14579));
INVX1 gate2693(.O (g3109), .I (g2482));
INVX1 gate2694(.O (g3791), .I (I7014));
INVX1 gate2695(.O (g2456), .I (g1397));
INVX1 gate2696(.O (g7919), .I (g7512));
INVX1 gate2697(.O (g10032), .I (I15232));
INVX1 gate2698(.O (g2529), .I (I5638));
INVX1 gate2699(.O (g2649), .I (g2005));
INVX1 gate2700(.O (g10140), .I (I15418));
INVX1 gate2701(.O (g4780), .I (g3440));
INVX1 gate2702(.O (I8839), .I (g4484));
INVX1 gate2703(.O (g6040), .I (I9655));
INVX1 gate2704(.O (g2348), .I (I5418));
INVX1 gate2705(.O (I6077), .I (g2349));
INVX1 gate2706(.O (g11574), .I (g11561));
INVX1 gate2707(.O (g11452), .I (I17413));
INVX1 gate2708(.O (g11047), .I (I16802));
INVX1 gate2709(.O (g5682), .I (I9199));
INVX1 gate2710(.O (g5766), .I (I9346));
INVX1 gate2711(.O (g5105), .I (I8487));
INVX1 gate2712(.O (g4509), .I (I7906));
INVX1 gate2713(.O (g6440), .I (g6150));
INVX1 gate2714(.O (g1976), .I (g643));
INVX1 gate2715(.O (g11205), .I (g11112));
INVX1 gate2716(.O (I6477), .I (g2069));
INVX1 gate2717(.O (I9632), .I (g5557));
INVX1 gate2718(.O (g7952), .I (g7427));
INVX1 gate2719(.O (I15311), .I (g10013));
INVX1 gate2720(.O (g9450), .I (g9097));
INVX1 gate2721(.O (g5305), .I (g4378));
INVX1 gate2722(.O (g5801), .I (g5320));
INVX1 gate2723(.O (I5734), .I (g2097));
INVX1 gate2724(.O (I6523), .I (g2819));
INVX1 gate2725(.O (g2155), .I (I5070));
INVX1 gate2726(.O (I4820), .I (g865));
INVX1 gate2727(.O (I17243), .I (g11396));
INVX1 gate2728(.O (g2355), .I (I5435));
INVX1 gate2729(.O (g2851), .I (I5979));
INVX1 gate2730(.O (I7249), .I (g2833));
INVX1 gate2731(.O (I12559), .I (g7477));
INVX1 gate2732(.O (I14315), .I (g8815));
INVX1 gate2733(.O (I6643), .I (g3008));
INVX1 gate2734(.O (g8213), .I (g7826));
INVX1 gate2735(.O (I10819), .I (g6706));
INVX1 gate2736(.O (g11311), .I (I17100));
INVX1 gate2737(.O (I10910), .I (g6703));
INVX1 gate2738(.O (I12424), .I (g7635));
INVX1 gate2739(.O (I9102), .I (g5586));
INVX1 gate2740(.O (I9208), .I (g5047));
INVX1 gate2741(.O (g3707), .I (g2920));
INVX1 gate2742(.O (I9302), .I (g5576));
INVX1 gate2743(.O (I14910), .I (g9532));
INVX1 gate2744(.O (g7616), .I (I12196));
INVX1 gate2745(.O (g7561), .I (I12015));
INVX1 gate2746(.O (g4067), .I (I7194));
INVX1 gate2747(.O (g3759), .I (I6958));
INVX1 gate2748(.O (I8278), .I (g4495));
INVX1 gate2749(.O (I14257), .I (g8805));
INVX1 gate2750(.O (g5748), .I (I9320));
INVX1 gate2751(.O (I10979), .I (g6565));
INVX1 gate2752(.O (g2964), .I (I6193));
INVX1 gate2753(.O (g4418), .I (I7760));
INVX1 gate2754(.O (I9869), .I (g5405));
INVX1 gate2755(.O (g4467), .I (g3829));
INVX1 gate2756(.O (I15072), .I (g9713));
INVX1 gate2757(.O (I14979), .I (g9671));
INVX1 gate2758(.O (g4290), .I (g3586));
INVX1 gate2759(.O (I10111), .I (g5754));
INVX1 gate2760(.O (I14055), .I (g8650));
INVX1 gate2761(.O (g10871), .I (I16583));
INVX1 gate2762(.O (g11051), .I (I16814));
INVX1 gate2763(.O (I5992), .I (g2195));
INVX1 gate2764(.O (g7004), .I (I11143));
INVX1 gate2765(.O (I16583), .I (g10848));
INVX1 gate2766(.O (g11072), .I (g10913));
INVX1 gate2767(.O (I17773), .I (g11650));
INVX1 gate2768(.O (I15592), .I (g10163));
INVX1 gate2769(.O (I15756), .I (g10266));
INVX1 gate2770(.O (g7527), .I (g7148));
INVX1 gate2771(.O (I17268), .I (g11351));
INVX1 gate2772(.O (I6742), .I (g3326));
INVX1 gate2773(.O (I12544), .I (g7669));
INVX1 gate2774(.O (g4093), .I (g2965));
INVX1 gate2775(.O (I8282), .I (g4770));
INVX1 gate2776(.O (g6151), .I (I9872));
INVX1 gate2777(.O (g7764), .I (I12457));
INVX1 gate2778(.O (g4256), .I (g3664));
INVX1 gate2779(.O (g6648), .I (I10607));
INVX1 gate2780(.O (g9777), .I (g9474));
INVX1 gate2781(.O (g7546), .I (I11970));
INVX1 gate2782(.O (I5080), .I (g36));
INVX1 gate2783(.O (I15350), .I (g10001));
INVX1 gate2784(.O (I10384), .I (g5842));
INVX1 gate2785(.O (g10162), .I (I15482));
INVX1 gate2786(.O (g3715), .I (g2920));
INVX1 gate2787(.O (I9265), .I (g5085));
INVX1 gate2788(.O (I16787), .I (g10896));
INVX1 gate2789(.O (g11350), .I (g11287));
INVX1 gate2790(.O (I5713), .I (g2436));
INVX1 gate2791(.O (I15820), .I (g10204));
INVX1 gate2792(.O (g5091), .I (g4385));
INVX1 gate2793(.O (g8056), .I (g7671));
INVX1 gate2794(.O (I13317), .I (g8093));
INVX1 gate2795(.O (I12610), .I (g7627));
INVX1 gate2796(.O (g4181), .I (I7360));
INVX1 gate2797(.O (I6754), .I (g2906));
INVX1 gate2798(.O (g8529), .I (I13738));
INVX1 gate2799(.O (I14094), .I (g8700));
INVX1 gate2800(.O (g4381), .I (g3914));
INVX1 gate2801(.O (g7925), .I (g7476));
INVX1 gate2802(.O (I9786), .I (g5396));
INVX1 gate2803(.O (g2118), .I (g1854));
INVX1 gate2804(.O (g8348), .I (I13424));
INVX1 gate2805(.O (I12255), .I (g7203));
INVX1 gate2806(.O (I6273), .I (g2482));
INVX1 gate2807(.O (g2872), .I (I6016));
INVX1 gate2808(.O (I16105), .I (g10382));
INVX1 gate2809(.O (g10629), .I (g10583));
INVX1 gate2810(.O (I10150), .I (g5705));
INVX1 gate2811(.O (g5169), .I (g4596));
INVX1 gate2812(.O (g4197), .I (I7408));
INVX1 gate2813(.O (I10801), .I (g6536));
INVX1 gate2814(.O (g8155), .I (I13048));
INVX1 gate2815(.O (g11396), .I (I17231));
INVX1 gate2816(.O (I13002), .I (g8045));
INVX1 gate2817(.O (g8355), .I (I13445));
INVX1 gate2818(.O (g10220), .I (I15592));
INVX1 gate2819(.O (g5007), .I (I8379));
INVX1 gate2820(.O (I13057), .I (g7843));
INVX1 gate2821(.O (g2652), .I (g2008));
INVX1 gate2822(.O (g2057), .I (g754));
INVX1 gate2823(.O (g10628), .I (I16307));
INVX1 gate2824(.O (I12678), .I (g7376));
INVX1 gate2825(.O (I13128), .I (g7976));
INVX1 gate2826(.O (g2843), .I (I5963));
INVX1 gate2827(.O (g10911), .I (I16685));
INVX1 gate2828(.O (g7320), .I (I11608));
INVX1 gate2829(.O (g2989), .I (g2135));
INVX1 gate2830(.O (g3539), .I (g3015));
INVX1 gate2831(.O (g4263), .I (g3586));
INVX1 gate2832(.O (I13245), .I (g8269));
INVX1 gate2833(.O (I11626), .I (g7042));
INVX1 gate2834(.O (I16769), .I (g10894));
INVX1 gate2835(.O (g5718), .I (I9256));
INVX1 gate2836(.O (I12460), .I (g7569));
INVX1 gate2837(.O (I12939), .I (g7977));
INVX1 gate2838(.O (g5767), .I (I9349));
INVX1 gate2839(.O (I15691), .I (g10233));
INVX1 gate2840(.O (I9296), .I (g4908));
INVX1 gate2841(.O (I10018), .I (g5862));
INVX1 gate2842(.O (I11299), .I (g6727));
INVX1 gate2843(.O (I13323), .I (g8203));
INVX1 gate2844(.O (I7176), .I (g2623));
INVX1 gate2845(.O (I5976), .I (g2186));
INVX1 gate2846(.O (g2549), .I (g1386));
INVX1 gate2847(.O (I6572), .I (g2853));
INVX1 gate2848(.O (I10526), .I (g6161));
INVX1 gate2849(.O (g8063), .I (I12907));
INVX1 gate2850(.O (g2834), .I (I5952));
INVX1 gate2851(.O (g2971), .I (g2046));
INVX1 gate2852(.O (g6172), .I (I9901));
INVX1 gate2853(.O (g6278), .I (I10093));
INVX1 gate2854(.O (g7617), .I (I12199));
INVX1 gate2855(.O (I7405), .I (g3861));
INVX1 gate2856(.O (g7906), .I (I12694));
INVX1 gate2857(.O (g7789), .I (I12532));
INVX1 gate2858(.O (g11405), .I (I17258));
INVX1 gate2859(.O (g5261), .I (g4640));
INVX1 gate2860(.O (g10591), .I (I16258));
INVX1 gate2861(.O (I6543), .I (g3186));
INVX1 gate2862(.O (g3362), .I (I6546));
INVX1 gate2863(.O (g3419), .I (g3104));
INVX1 gate2864(.O (I7829), .I (g3425));
INVX1 gate2865(.O (g6667), .I (I10630));
INVX1 gate2866(.O (g7516), .I (g7148));
INVX1 gate2867(.O (g4562), .I (I7973));
INVX1 gate2868(.O (g6343), .I (I10248));
INVX1 gate2869(.O (g10754), .I (I16439));
INVX1 gate2870(.O (g9353), .I (I14564));
INVX1 gate2871(.O (g3052), .I (I6264));
INVX1 gate2872(.O (g10355), .I (I15829));
INVX1 gate2873(.O (g5415), .I (I8848));
INVX1 gate2874(.O (g6282), .I (I10105));
INVX1 gate2875(.O (g7771), .I (I12478));
INVX1 gate2876(.O (g6566), .I (g5791));
INVX1 gate2877(.O (I11737), .I (g7027));
INVX1 gate2878(.O (g8279), .I (I13209));
INVX1 gate2879(.O (g2121), .I (I5041));
INVX1 gate2880(.O (g4631), .I (g3820));
INVX1 gate2881(.O (I12875), .I (g7638));
INVX1 gate2882(.O (g10825), .I (I16537));
INVX1 gate2883(.O (I10917), .I (g6732));
INVX1 gate2884(.O (I15583), .I (g10157));
INVX1 gate2885(.O (g9802), .I (g9490));
INVX1 gate2886(.O (g1999), .I (g806));
INVX1 gate2887(.O (I11232), .I (g6537));
INVX1 gate2888(.O (g4257), .I (g3664));
INVX1 gate2889(.O (g6134), .I (I9839));
INVX1 gate2890(.O (g5664), .I (I9153));
INVX1 gate2891(.O (g8318), .I (I13338));
INVX1 gate2892(.O (g8872), .I (I14188));
INVX1 gate2893(.O (I9706), .I (g5221));
INVX1 gate2894(.O (g2232), .I (I5221));
INVX1 gate2895(.O (g10172), .I (I15510));
INVX1 gate2896(.O (g11046), .I (I16799));
INVX1 gate2897(.O (g3086), .I (g2276));
INVX1 gate2898(.O (g5203), .I (g4640));
INVX1 gate2899(.O (g2253), .I (g100));
INVX1 gate2900(.O (g3728), .I (I6904));
INVX1 gate2901(.O (g2813), .I (I5913));
INVX1 gate2902(.O (I9029), .I (g4781));
INVX1 gate2903(.O (g8989), .I (I14388));
INVX1 gate2904(.O (I14077), .I (g8758));
INVX1 gate2905(.O (I9171), .I (g4902));
INVX1 gate2906(.O (g6555), .I (g5740));
INVX1 gate2907(.O (I10706), .I (g6080));
INVX1 gate2908(.O (I9371), .I (g5075));
INVX1 gate2909(.O (g6804), .I (I10822));
INVX1 gate2910(.O (I15787), .I (g10269));
INVX1 gate2911(.O (I6414), .I (g2342));
INVX1 gate2912(.O (g3730), .I (g3015));
INVX1 gate2913(.O (g2909), .I (I6080));
INVX1 gate2914(.O (I9956), .I (g5485));
INVX1 gate2915(.O (I10689), .I (g6059));
INVX1 gate2916(.O (g3385), .I (g3121));
INVX1 gate2917(.O (I5383), .I (g886));
INVX1 gate2918(.O (I15302), .I (g10007));
INVX1 gate2919(.O (g11357), .I (I17182));
INVX1 gate2920(.O (g7991), .I (I12809));
INVX1 gate2921(.O (I6513), .I (g2812));
INVX1 gate2922(.O (g2606), .I (I5719));
INVX1 gate2923(.O (g10319), .I (g10270));
INVX1 gate2924(.O (g4441), .I (g3914));
INVX1 gate2925(.O (g6113), .I (I9792));
INVX1 gate2926(.O (g6313), .I (I10198));
INVX1 gate2927(.O (g7078), .I (I11309));
INVX1 gate2928(.O (g7340), .I (I11668));
INVX1 gate2929(.O (I10102), .I (g5730));
INVX1 gate2930(.O (I16778), .I (g10891));
INVX1 gate2931(.O (I13831), .I (g8560));
INVX1 gate2932(.O (g10318), .I (I15752));
INVX1 gate2933(.O (I8050), .I (g4089));
INVX1 gate2934(.O (I13445), .I (g8149));
INVX1 gate2935(.O (I5588), .I (g1203));
INVX1 gate2936(.O (g8121), .I (I12978));
INVX1 gate2937(.O (g10227), .I (I15601));
INVX1 gate2938(.O (g7907), .I (g7664));
INVX1 gate2939(.O (I6436), .I (g2351));
INVX1 gate2940(.O (I6679), .I (g2902));
INVX1 gate2941(.O (g8321), .I (I13347));
INVX1 gate2942(.O (g4673), .I (g4013));
INVX1 gate2943(.O (g6202), .I (g5426));
INVX1 gate2944(.O (g8670), .I (g8551));
INVX1 gate2945(.O (g5689), .I (I9216));
INVX1 gate2946(.O (I8996), .I (g4757));
INVX1 gate2947(.O (I9684), .I (g5426));
INVX1 gate2948(.O (g7035), .I (I11194));
INVX1 gate2949(.O (I15768), .I (g10249));
INVX1 gate2950(.O (I9138), .I (g5210));
INVX1 gate2951(.O (I9639), .I (g5126));
INVX1 gate2952(.O (g7959), .I (I12751));
INVX1 gate2953(.O (I10066), .I (g5778));
INVX1 gate2954(.O (I9338), .I (g5576));
INVX1 gate2955(.O (I10231), .I (g6111));
INVX1 gate2956(.O (g8625), .I (g8487));
INVX1 gate2957(.O (g7082), .I (I11315));
INVX1 gate2958(.O (g2586), .I (g1972));
INVX1 gate2959(.O (g5216), .I (g4445));
INVX1 gate2960(.O (g10540), .I (I16187));
INVX1 gate2961(.O (I17410), .I (g11419));
INVX1 gate2962(.O (g6094), .I (I9749));
INVX1 gate2963(.O (I11498), .I (g6578));
INVX1 gate2964(.O (I12595), .I (g7706));
INVX1 gate2965(.O (I16647), .I (g10866));
INVX1 gate2966(.O (g10058), .I (I15281));
INVX1 gate2967(.O (I16356), .I (g10597));
INVX1 gate2968(.O (g4669), .I (g4013));
INVX1 gate2969(.O (I8724), .I (g4791));
INVX1 gate2970(.O (g6567), .I (I10495));
INVX1 gate2971(.O (g5671), .I (I9174));
INVX1 gate2972(.O (g4368), .I (I7665));
INVX1 gate2973(.O (I11989), .I (g6919));
INVX1 gate2974(.O (I17666), .I (g11603));
INVX1 gate2975(.O (I10885), .I (g6332));
INVX1 gate2976(.O (I8379), .I (g4231));
INVX1 gate2977(.O (g3331), .I (I6510));
INVX1 gate2978(.O (g10203), .I (g10177));
INVX1 gate2979(.O (I14876), .I (g9526));
INVX1 gate2980(.O (I11611), .I (g6913));
INVX1 gate2981(.O (g7656), .I (I12265));
INVX1 gate2982(.O (g4772), .I (g3440));
INVX1 gate2983(.O (g3406), .I (I6611));
INVX1 gate2984(.O (I11722), .I (g7034));
INVX1 gate2985(.O (I7399), .I (g4113));
INVX1 gate2986(.O (g10044), .I (I15263));
INVX1 gate2987(.O (g3635), .I (I6812));
INVX1 gate2988(.O (I6022), .I (g2258));
INVX1 gate2989(.O (g4458), .I (I7817));
INVX1 gate2990(.O (g2570), .I (g207));
INVX1 gate2991(.O (g2860), .I (I5998));
INVX1 gate2992(.O (g2341), .I (I5403));
INVX1 gate2993(.O (g9262), .I (I14473));
INVX1 gate2994(.O (g3682), .I (g2920));
INVX1 gate2995(.O (g6593), .I (I10557));
INVX1 gate2996(.O (I9759), .I (g5344));
INVX1 gate2997(.O (g8519), .I (I13726));
INVX1 gate2998(.O (g3105), .I (g2482));
INVX1 gate2999(.O (g7915), .I (g7473));
INVX1 gate3000(.O (g3305), .I (I6474));
INVX1 gate3001(.O (g10281), .I (g10162));
INVX1 gate3002(.O (g98), .I (I4783));
INVX1 gate3003(.O (g2645), .I (g1991));
INVX1 gate3004(.O (I8835), .I (g4791));
INVX1 gate3005(.O (g5826), .I (I9440));
INVX1 gate3006(.O (I12418), .I (g7568));
INVX1 gate3007(.O (I12822), .I (g7677));
INVX1 gate3008(.O (g10902), .I (I16660));
INVX1 gate3009(.O (g10377), .I (I15855));
INVX1 gate3010(.O (g8606), .I (g8481));
INVX1 gate3011(.O (g7214), .I (I11450));
INVX1 gate3012(.O (I6947), .I (g2860));
INVX1 gate3013(.O (g10120), .I (I15368));
INVX1 gate3014(.O (g4011), .I (I7151));
INVX1 gate3015(.O (g9076), .I (g8892));
INVX1 gate3016(.O (g5741), .I (I9305));
INVX1 gate3017(.O (g3748), .I (g2971));
INVX1 gate3018(.O (g4411), .I (I7743));
INVX1 gate3019(.O (g4734), .I (g3586));
INVX1 gate3020(.O (I11342), .I (g6686));
INVX1 gate3021(.O (g9889), .I (I15072));
INVX1 gate3022(.O (g7110), .I (I11345));
INVX1 gate3023(.O (g6264), .I (I10051));
INVX1 gate3024(.O (g7310), .I (I11578));
INVX1 gate3025(.O (I6560), .I (g2845));
INVX1 gate3026(.O (I7291), .I (g3212));
INVX1 gate3027(.O (I8611), .I (g4562));
INVX1 gate3028(.O (I10456), .I (g5844));
INVX1 gate3029(.O (I15482), .I (g10115));
INVX1 gate3030(.O (g5638), .I (I9077));
INVX1 gate3031(.O (g3226), .I (I6403));
INVX1 gate3032(.O (g6933), .I (I11061));
INVX1 gate3033(.O (g7663), .I (I12282));
INVX1 gate3034(.O (I11650), .I (g6938));
INVX1 gate3035(.O (g10699), .I (I16376));
INVX1 gate3036(.O (g2607), .I (I5722));
INVX1 gate3037(.O (I12853), .I (g7638));
INVX1 gate3038(.O (I16897), .I (g10947));
INVX1 gate3039(.O (I5240), .I (g64));
INVX1 gate3040(.O (g2962), .I (I6183));
INVX1 gate3041(.O (g6521), .I (I10437));
INVX1 gate3042(.O (I17084), .I (g11249));
INVX1 gate3043(.O (g4474), .I (g3820));
INVX1 gate3044(.O (g10290), .I (I15694));
INVX1 gate3045(.O (g2158), .I (I5077));
INVX1 gate3046(.O (g6050), .I (I9677));
INVX1 gate3047(.O (g6641), .I (I10598));
INVX1 gate3048(.O (I11198), .I (g6521));
INVX1 gate3049(.O (I9498), .I (g5081));
INVX1 gate3050(.O (I12589), .I (g7571));
INVX1 gate3051(.O (g10698), .I (I16373));
INVX1 gate3052(.O (g2506), .I (g636));
INVX1 gate3053(.O (g6450), .I (I10378));
INVX1 gate3054(.O (I6037), .I (g2560));
INVX1 gate3055(.O (I17321), .I (g11348));
INVX1 gate3056(.O (g5883), .I (g5309));
INVX1 gate3057(.O (I10314), .I (g6251));
INVX1 gate3058(.O (g7402), .I (g6860));
INVX1 gate3059(.O (I6495), .I (g2076));
INVX1 gate3060(.O (I9833), .I (g5197));
INVX1 gate3061(.O (I17179), .I (g11307));
INVX1 gate3062(.O (I11528), .I (g6796));
INVX1 gate3063(.O (I6102), .I (g2240));
INVX1 gate3064(.O (I16717), .I (g10779));
INVX1 gate3065(.O (I17531), .I (g11488));
INVX1 gate3066(.O (I7694), .I (g3742));
INVX1 gate3067(.O (I11330), .I (g6571));
INVX1 gate3068(.O (I6302), .I (g2243));
INVX1 gate3069(.O (g3373), .I (I6565));
INVX1 gate3070(.O (I15778), .I (g10255));
INVX1 gate3071(.O (g7762), .I (I12451));
INVX1 gate3072(.O (g3491), .I (g2669));
INVX1 gate3073(.O (g4080), .I (g2903));
INVX1 gate3074(.O (I5116), .I (g40));
INVX1 gate3075(.O (g11081), .I (I16856));
INVX1 gate3076(.O (I7852), .I (g3438));
INVX1 gate3077(.O (I7923), .I (g3394));
INVX1 gate3078(.O (g5758), .I (I9338));
INVX1 gate3079(.O (g8141), .I (I13020));
INVX1 gate3080(.O (g8570), .I (I13803));
INVX1 gate3081(.O (g5066), .I (I8436));
INVX1 gate3082(.O (g5589), .I (I9001));
INVX1 gate3083(.O (g6724), .I (I10719));
INVX1 gate3084(.O (g8341), .I (I13403));
INVX1 gate3085(.O (I10054), .I (g5728));
INVX1 gate3086(.O (g2275), .I (g757));
INVX1 gate3087(.O (I9539), .I (g5354));
INVX1 gate3088(.O (I9896), .I (g5295));
INVX1 gate3089(.O (g4713), .I (g3546));
INVX1 gate3090(.O (I10243), .I (g5918));
INVX1 gate3091(.O (I11132), .I (g6451));
INVX1 gate3092(.O (I11869), .I (g6894));
INVX1 gate3093(.O (g7877), .I (g7479));
INVX1 gate3094(.O (I7701), .I (g3513));
INVX1 gate3095(.O (g3369), .I (I6557));
INVX1 gate3096(.O (I5565), .I (g1713));
INVX1 gate3097(.O (g3007), .I (I6240));
INVX1 gate3098(.O (g9339), .I (I14522));
INVX1 gate3099(.O (I15356), .I (g10013));
INVX1 gate3100(.O (g7657), .I (I12268));
INVX1 gate3101(.O (g6878), .I (I10966));
INVX1 gate3102(.O (I15826), .I (g10205));
INVX1 gate3103(.O (I6917), .I (g2832));
INVX1 gate3104(.O (I15380), .I (g10098));
INVX1 gate3105(.O (I4894), .I (g258));
INVX1 gate3106(.O (g2174), .I (g31));
INVX1 gate3107(.O (g3459), .I (I6661));
INVX1 gate3108(.O (g6289), .I (I10126));
INVX1 gate3109(.O (g9024), .I (I14409));
INVX1 gate3110(.O (g2374), .I (g591));
INVX1 gate3111(.O (I12616), .I (g7534));
INVX1 gate3112(.O (I9162), .I (g5035));
INVX1 gate3113(.O (g7556), .I (I11992));
INVX1 gate3114(.O (I9268), .I (g5305));
INVX1 gate3115(.O (I16723), .I (g10851));
INVX1 gate3116(.O (g3767), .I (I6976));
INVX1 gate3117(.O (g10547), .I (I16206));
INVX1 gate3118(.O (g9424), .I (g9076));
INVX1 gate3119(.O (g10895), .I (I16647));
INVX1 gate3120(.O (I7886), .I (g4076));
INVX1 gate3121(.O (I9362), .I (g5013));
INVX1 gate3122(.O (g6835), .I (I10885));
INVX1 gate3123(.O (g2985), .I (I6217));
INVX1 gate3124(.O (g9809), .I (I14944));
INVX1 gate3125(.O (g5827), .I (I9443));
INVX1 gate3126(.O (g6882), .I (I10974));
INVX1 gate3127(.O (g7928), .I (g7508));
INVX1 gate3128(.O (I10156), .I (g6100));
INVX1 gate3129(.O (I10655), .I (g6036));
INVX1 gate3130(.O (I15672), .I (g10132));
INVX1 gate3131(.O (g3582), .I (g3164));
INVX1 gate3132(.O (I16387), .I (g10629));
INVX1 gate3133(.O (I17334), .I (g11360));
INVX1 gate3134(.O (g6271), .I (I10072));
INVX1 gate3135(.O (I11225), .I (g6534));
INVX1 gate3136(.O (g10226), .I (I15598));
INVX1 gate3137(.O (I9452), .I (g5085));
INVX1 gate3138(.O (g11182), .I (I16947));
INVX1 gate3139(.O (g11651), .I (I17755));
INVX1 gate3140(.O (g7064), .I (I11269));
INVX1 gate3141(.O (I5210), .I (g58));
INVX1 gate3142(.O (g2239), .I (I5240));
INVX1 gate3143(.O (I10180), .I (g6107));
INVX1 gate3144(.O (g9672), .I (I14805));
INVX1 gate3145(.O (I13708), .I (g8337));
INVX1 gate3146(.O (g5774), .I (I9362));
INVX1 gate3147(.O (g7899), .I (I12683));
INVX1 gate3148(.O (g3793), .I (g2593));
INVX1 gate3149(.O (g7464), .I (I11858));
INVX1 gate3150(.O (I12053), .I (g6928));
INVX1 gate3151(.O (g8358), .I (I13454));
INVX1 gate3152(.O (I12809), .I (g7686));
INVX1 gate3153(.O (g7785), .I (I12520));
INVX1 gate3154(.O (I16811), .I (g10908));
INVX1 gate3155(.O (g10551), .I (I16214));
INVX1 gate3156(.O (I6233), .I (g2299));
INVX1 gate3157(.O (g2832), .I (I5946));
INVX1 gate3158(.O (I12466), .I (g7585));
INVX1 gate3159(.O (g3415), .I (g3121));
INVX1 gate3160(.O (g3227), .I (I6406));
INVX1 gate3161(.O (I7825), .I (g3414));
INVX1 gate3162(.O (g6799), .I (I10807));
INVX1 gate3163(.O (g2853), .I (g2171));
INVX1 gate3164(.O (I11043), .I (g6412));
INVX1 gate3165(.O (I6454), .I (g2368));
INVX1 gate3166(.O (I13043), .I (g8055));
INVX1 gate3167(.O (I17216), .I (g11291));
INVX1 gate3168(.O (g2420), .I (g237));
INVX1 gate3169(.O (g6674), .I (I10639));
INVX1 gate3170(.O (I9486), .I (g5066));
INVX1 gate3171(.O (g11513), .I (I17558));
INVX1 gate3172(.O (I12177), .I (g7259));
INVX1 gate3173(.O (g10127), .I (I15383));
INVX1 gate3174(.O (g3664), .I (g3209));
INVX1 gate3175(.O (g8275), .I (I13197));
INVX1 gate3176(.O (g2507), .I (I5584));
INVX1 gate3177(.O (g8311), .I (I13317));
INVX1 gate3178(.O (g3246), .I (g2482));
INVX1 gate3179(.O (I15448), .I (g10056));
INVX1 gate3180(.O (g5509), .I (g4739));
INVX1 gate3181(.O (g4326), .I (g3863));
INVX1 gate3182(.O (I14694), .I (g9259));
INVX1 gate3183(.O (I7408), .I (g4125));
INVX1 gate3184(.O (g7237), .I (I11477));
INVX1 gate3185(.O (g10490), .I (I16105));
INVX1 gate3186(.O (I9185), .I (g4915));
INVX1 gate3187(.O (I7336), .I (g3997));
INVX1 gate3188(.O (g3721), .I (I6891));
INVX1 gate3189(.O (g11505), .I (I17534));
INVX1 gate3190(.O (I11602), .I (g6833));
INVX1 gate3191(.O (I11810), .I (g7246));
INVX1 gate3192(.O (g11404), .I (I17255));
INVX1 gate3193(.O (g6132), .I (I9833));
INVX1 gate3194(.O (g5662), .I (I9147));
INVX1 gate3195(.O (I6553), .I (g3186));
INVX1 gate3196(.O (I4850), .I (g1958));
INVX1 gate3197(.O (g7844), .I (I12631));
INVX1 gate3198(.O (I17543), .I (g11499));
INVX1 gate3199(.O (I11068), .I (g6426));
INVX1 gate3200(.O (I13068), .I (g7906));
INVX1 gate3201(.O (g6680), .I (I10643));
INVX1 gate3202(.O (g6209), .I (I9956));
INVX1 gate3203(.O (g8985), .I (I14376));
INVX1 gate3204(.O (I11879), .I (g6893));
INVX1 gate3205(.O (g5994), .I (I9612));
INVX1 gate3206(.O (g10889), .I (I16629));
INVX1 gate3207(.O (I16850), .I (g10905));
INVX1 gate3208(.O (I11970), .I (g6918));
INVX1 gate3209(.O (g7394), .I (I11778));
INVX1 gate3210(.O (I10557), .I (g6197));
INVX1 gate3211(.O (g10354), .I (I15826));
INVX1 gate3212(.O (g2905), .I (I6068));
INVX1 gate3213(.O (g7089), .I (I11322));
INVX1 gate3214(.O (g7731), .I (I12376));
INVX1 gate3215(.O (g10888), .I (I16626));
INVX1 gate3216(.O (g6802), .I (I10816));
INVX1 gate3217(.O (g8239), .I (g7826));
INVX1 gate3218(.O (g4183), .I (I7366));
INVX1 gate3219(.O (g9273), .I (I14490));
INVX1 gate3220(.O (g4608), .I (g3829));
INVX1 gate3221(.O (g5816), .I (I9424));
INVX1 gate3222(.O (I5922), .I (g2170));
INVX1 gate3223(.O (I7465), .I (g3726));
INVX1 gate3224(.O (g7966), .I (I12762));
INVX1 gate3225(.O (g2100), .I (I4948));
INVX1 gate3226(.O (I10278), .I (g5815));
INVX1 gate3227(.O (g3940), .I (g2920));
INVX1 gate3228(.O (g6558), .I (I10484));
INVX1 gate3229(.O (I12009), .I (g6915));
INVX1 gate3230(.O (I6888), .I (g2960));
INVX1 gate3231(.O (I8262), .I (g4636));
INVX1 gate3232(.O (I11967), .I (g6911));
INVX1 gate3233(.O (g8020), .I (I12862));
INVX1 gate3234(.O (I10286), .I (g6237));
INVX1 gate3235(.O (g8420), .I (I13574));
INVX1 gate3236(.O (I5060), .I (g1191));
INVX1 gate3237(.O (g10931), .I (g10827));
INVX1 gate3238(.O (g3388), .I (I6590));
INVX1 gate3239(.O (I10039), .I (g5718));
INVX1 gate3240(.O (I14306), .I (g8812));
INVX1 gate3241(.O (I11459), .I (g6488));
INVX1 gate3242(.O (g11433), .I (I17350));
INVX1 gate3243(.O (g9572), .I (I14709));
INVX1 gate3244(.O (g5685), .I (I9208));
INVX1 gate3245(.O (g5197), .I (I8611));
INVX1 gate3246(.O (g5700), .I (I9237));
INVX1 gate3247(.O (g8794), .I (I14109));
INVX1 gate3248(.O (g5397), .I (I8835));
INVX1 gate3249(.O (g2750), .I (I5818));
INVX1 gate3250(.O (I8889), .I (g4553));
INVX1 gate3251(.O (g11620), .I (I17678));
INVX1 gate3252(.O (g10190), .I (I15548));
INVX1 gate3253(.O (I8476), .I (g4577));
INVX1 gate3254(.O (g4361), .I (I7648));
INVX1 gate3255(.O (I9766), .I (g5348));
INVX1 gate3256(.O (I15811), .I (g10200));
INVX1 gate3257(.O (g3428), .I (I6639));
INVX1 gate3258(.O (I7096), .I (g3186));
INVX1 gate3259(.O (I12454), .I (g7544));
INVX1 gate3260(.O (I9087), .I (g5113));
INVX1 gate3261(.O (I9105), .I (g5589));
INVX1 gate3262(.O (I9305), .I (g4970));
INVX1 gate3263(.O (I9801), .I (g5416));
INVX1 gate3264(.O (g3430), .I (I6643));
INVX1 gate3265(.O (g7814), .I (I12607));
INVX1 gate3266(.O (I12712), .I (g7441));
INVX1 gate3267(.O (g11646), .I (I17742));
INVX1 gate3268(.O (g4051), .I (I7166));
INVX1 gate3269(.O (I10601), .I (g5996));
INVX1 gate3270(.O (I13010), .I (g8047));
INVX1 gate3271(.O (g11343), .I (I17152));
INVX1 gate3272(.O (I13918), .I (g8451));
INVX1 gate3273(.O (I16379), .I (g10598));
INVX1 gate3274(.O (g4127), .I (I7276));
INVX1 gate3275(.O (g4451), .I (g3638));
INVX1 gate3276(.O (I15971), .I (g10408));
INVX1 gate3277(.O (g4327), .I (I7600));
INVX1 gate3278(.O (I17265), .I (g11352));
INVX1 gate3279(.O (g7350), .I (I11698));
INVX1 gate3280(.O (g2040), .I (g1786));
INVX1 gate3281(.O (g6574), .I (I10514));
INVX1 gate3282(.O (I12907), .I (g7959));
INVX1 gate3283(.O (I5995), .I (g2196));
INVX1 gate3284(.O (I11079), .I (g6649));
INVX1 gate3285(.O (g10546), .I (I16203));
INVX1 gate3286(.O (g7038), .I (I11201));
INVX1 gate3287(.O (I11444), .I (g6653));
INVX1 gate3288(.O (I17416), .I (g11420));
INVX1 gate3289(.O (g10211), .I (I15583));
INVX1 gate3290(.O (g9534), .I (I14687));
INVX1 gate3291(.O (g9961), .I (I15162));
INVX1 gate3292(.O (g6714), .I (g5867));
INVX1 gate3293(.O (g7438), .I (g7232));
INVX1 gate3294(.O (g7773), .I (I12484));
INVX1 gate3295(.O (I11599), .I (g6832));
INVX1 gate3296(.O (g7009), .I (I11152));
INVX1 gate3297(.O (g11369), .I (I17194));
INVX1 gate3298(.O (g2123), .I (I5047));
INVX1 gate3299(.O (I6639), .I (g2632));
INVX1 gate3300(.O (g4346), .I (I7625));
INVX1 gate3301(.O (g8515), .I (I13714));
INVX1 gate3302(.O (g10088), .I (I15317));
INVX1 gate3303(.O (I8285), .I (g4771));
INVX1 gate3304(.O (I10937), .I (g6552));
INVX1 gate3305(.O (I12239), .I (g7073));
INVX1 gate3306(.O (I5840), .I (g2432));
INVX1 gate3307(.O (I15368), .I (g9990));
INVX1 gate3308(.O (I17510), .I (g11481));
INVX1 gate3309(.O (I16742), .I (g10857));
INVX1 gate3310(.O (g8100), .I (g7947));
INVX1 gate3311(.O (I16944), .I (g11079));
INVX1 gate3312(.O (g3910), .I (g3015));
INVX1 gate3313(.O (I13086), .I (g7924));
INVX1 gate3314(.O (g7769), .I (I12472));
INVX1 gate3315(.O (I15412), .I (g10075));
INVX1 gate3316(.O (g3638), .I (I6821));
INVX1 gate3317(.O (I8139), .I (g3681));
INVX1 gate3318(.O (g7212), .I (I11444));
INVX1 gate3319(.O (g5723), .I (I9265));
INVX1 gate3320(.O (I14884), .I (g9454));
INVX1 gate3321(.O (g11412), .I (I17277));
INVX1 gate3322(.O (I11817), .I (g7246));
INVX1 gate3323(.O (I10168), .I (g5982));
INVX1 gate3324(.O (g5101), .I (I8473));
INVX1 gate3325(.O (g5817), .I (I9427));
INVX1 gate3326(.O (I11322), .I (g6652));
INVX1 gate3327(.O (g7918), .I (g7505));
INVX1 gate3328(.O (g5301), .I (g4373));
INVX1 gate3329(.O (g7967), .I (I12765));
INVX1 gate3330(.O (g6262), .I (I10045));
INVX1 gate3331(.O (I15229), .I (g9968));
INVX1 gate3332(.O (g2351), .I (I5427));
INVX1 gate3333(.O (I11159), .I (g6478));
INVX1 gate3334(.O (g10700), .I (I16379));
INVX1 gate3335(.O (g2648), .I (I5765));
INVX1 gate3336(.O (I9491), .I (g5072));
INVX1 gate3337(.O (g10126), .I (I15380));
INVX1 gate3338(.O (I8024), .I (g4117));
INVX1 gate3339(.O (I11901), .I (g6897));
INVX1 gate3340(.O (I16802), .I (g10902));
INVX1 gate3341(.O (g2530), .I (I5641));
INVX1 gate3342(.O (g6736), .I (I10739));
INVX1 gate3343(.O (I13125), .I (g7975));
INVX1 gate3344(.O (g8750), .I (I14045));
INVX1 gate3345(.O (I10666), .I (g6042));
INVX1 gate3346(.O (g4508), .I (g3946));
INVX1 gate3347(.O (g10250), .I (g10136));
INVX1 gate3348(.O (g2655), .I (g2013));
INVX1 gate3349(.O (g4944), .I (g4430));
INVX1 gate3350(.O (g4240), .I (g3664));
INVX1 gate3351(.O (I11783), .I (g7246));
INVX1 gate3352(.O (I16793), .I (g11014));
INVX1 gate3353(.O (I7342), .I (g4011));
INVX1 gate3354(.O (I9602), .I (g5013));
INVX1 gate3355(.O (g4472), .I (I7847));
INVX1 gate3356(.O (I10015), .I (g5641));
INVX1 gate3357(.O (I5704), .I (g2056));
INVX1 gate3358(.O (g7993), .I (I12813));
INVX1 gate3359(.O (I7255), .I (g3227));
INVX1 gate3360(.O (g6076), .I (I9717));
INVX1 gate3361(.O (I4906), .I (g119));
INVX1 gate3362(.O (I11656), .I (g7122));
INVX1 gate3363(.O (I6049), .I (g2219));
INVX1 gate3364(.O (g5751), .I (I9323));
INVX1 gate3365(.O (g3758), .I (I6955));
INVX1 gate3366(.O (g3066), .I (g2135));
INVX1 gate3367(.O (I8231), .I (g4170));
INVX1 gate3368(.O (g4443), .I (g3359));
INVX1 gate3369(.O (g10296), .I (I15708));
INVX1 gate3370(.O (g8440), .I (I13618));
INVX1 gate3371(.O (I11680), .I (g7064));
INVX1 gate3372(.O (g8969), .I (I14340));
INVX1 gate3373(.O (I17116), .I (g11229));
INVX1 gate3374(.O (g2410), .I (g1453));
INVX1 gate3375(.O (g9679), .I (g9452));
INVX1 gate3376(.O (I7726), .I (g3378));
INVX1 gate3377(.O (g6175), .I (g5320));
INVX1 gate3378(.O (g4116), .I (I7260));
INVX1 gate3379(.O (I7154), .I (g2617));
INVX1 gate3380(.O (g8323), .I (I13351));
INVX1 gate3381(.O (g6871), .I (g6724));
INVX1 gate3382(.O (g2884), .I (I6040));
INVX1 gate3383(.O (I7354), .I (g4066));
INVX1 gate3384(.O (g2839), .I (I5957));
INVX1 gate3385(.O (g3365), .I (I6553));
INVX1 gate3386(.O (g3861), .I (I7054));
INVX1 gate3387(.O (I6498), .I (g2958));
INVX1 gate3388(.O (I17746), .I (g11643));
INVX1 gate3389(.O (g3055), .I (g2135));
INVX1 gate3390(.O (I5053), .I (g1188));
INVX1 gate3391(.O (I15959), .I (g10402));
INVX1 gate3392(.O (g6285), .I (I10114));
INVX1 gate3393(.O (g11627), .I (I17695));
INVX1 gate3394(.O (g7921), .I (g7463));
INVX1 gate3395(.O (g10197), .I (I15565));
INVX1 gate3396(.O (g5673), .I (I9180));
INVX1 gate3397(.O (g4347), .I (g3880));
INVX1 gate3398(.O (I8551), .I (g4342));
INVX1 gate3399(.O (I10084), .I (g5742));
INVX1 gate3400(.O (g2172), .I (g43));
INVX1 gate3401(.O (g3333), .I (g2779));
INVX1 gate3402(.O (I9415), .I (g5047));
INVX1 gate3403(.O (g11112), .I (I16897));
INVX1 gate3404(.O (I17237), .I (g11394));
INVX1 gate3405(.O (g4681), .I (g3546));
INVX1 gate3406(.O (g10870), .I (I16580));
INVX1 gate3407(.O (g11050), .I (I16811));
INVX1 gate3408(.O (I8499), .I (g4330));
INVX1 gate3409(.O (I12577), .I (g7532));
INVX1 gate3410(.O (g8151), .I (g8036));
INVX1 gate3411(.O (g10527), .I (g10462));
INVX1 gate3412(.O (g3774), .I (I6999));
INVX1 gate3413(.O (g8351), .I (I13433));
INVX1 gate3414(.O (I17340), .I (g11366));
INVX1 gate3415(.O (g4533), .I (I7938));
INVX1 gate3416(.O (I13017), .I (g7848));
INVX1 gate3417(.O (I13364), .I (g8221));
INVX1 gate3418(.O (I15386), .I (g10101));
INVX1 gate3419(.O (g6184), .I (I9915));
INVX1 gate3420(.O (g2235), .I (g96));
INVX1 gate3421(.O (g2343), .I (g1927));
INVX1 gate3422(.O (I12439), .I (g7663));
INVX1 gate3423(.O (g5669), .I (I9168));
INVX1 gate3424(.O (I10531), .I (g6169));
INVX1 gate3425(.O (I17684), .I (g11609));
INVX1 gate3426(.O (g6339), .I (I10240));
INVX1 gate3427(.O (I14179), .I (g8785));
INVX1 gate3428(.O (g4210), .I (I7447));
INVX1 gate3429(.O (I14531), .I (g9273));
INVX1 gate3430(.O (I7112), .I (g3186));
INVX1 gate3431(.O (I17142), .I (g11301));
INVX1 gate3432(.O (g11096), .I (I16879));
INVX1 gate3433(.O (g7620), .I (I12208));
INVX1 gate3434(.O (g4596), .I (I8007));
INVX1 gate3435(.O (g3538), .I (I6726));
INVX1 gate3436(.O (I6019), .I (g2554));
INVX1 gate3437(.O (g4013), .I (I7157));
INVX1 gate3438(.O (g6424), .I (g6140));
INVX1 gate3439(.O (I16626), .I (g10859));
INVX1 gate3440(.O (I10186), .I (g6110));
INVX1 gate3441(.O (g6737), .I (g6016));
INVX1 gate3442(.O (g10867), .I (I16571));
INVX1 gate3443(.O (g2334), .I (I5388));
INVX1 gate3444(.O (g10894), .I (I16644));
INVX1 gate3445(.O (g6809), .I (I10837));
INVX1 gate3446(.O (I10685), .I (g6054));
INVX1 gate3447(.O (g5743), .I (I9311));
INVX1 gate3448(.O (g4413), .I (I7749));
INVX1 gate3449(.O (g5890), .I (g5361));
INVX1 gate3450(.O (I11289), .I (g6508));
INVX1 gate3451(.O (I6052), .I (g2220));
INVX1 gate3452(.O (g2548), .I (I5667));
INVX1 gate3453(.O (I14373), .I (g8956));
INVX1 gate3454(.O (I11309), .I (g6531));
INVX1 gate3455(.O (I5929), .I (g2225));
INVX1 gate3456(.O (I13023), .I (g8050));
INVX1 gate3457(.O (g8884), .I (I14224));
INVX1 gate3458(.O (I16298), .I (g10553));
INVX1 gate3459(.O (I13224), .I (g8261));
INVX1 gate3460(.O (g7788), .I (I12529));
INVX1 gate3461(.O (g6077), .I (I9720));
INVX1 gate3462(.O (g11429), .I (I17340));
INVX1 gate3463(.O (g5011), .I (I8385));
INVX1 gate3464(.O (I16775), .I (g10889));
INVX1 gate3465(.O (g3067), .I (I6273));
INVX1 gate3466(.O (I13571), .I (g8355));
INVX1 gate3467(.O (g10315), .I (g10243));
INVX1 gate3468(.O (g5856), .I (g5245));
INVX1 gate3469(.O (g5734), .I (I9290));
INVX1 gate3470(.O (g10819), .I (I16525));
INVX1 gate3471(.O (g11428), .I (I17337));
INVX1 gate3472(.O (g10910), .I (I16682));
INVX1 gate3473(.O (g3290), .I (I6461));
INVX1 gate3474(.O (I17362), .I (g11376));
INVX1 gate3475(.O (g10202), .I (g10171));
INVX1 gate3476(.O (I10334), .I (g6003));
INVX1 gate3477(.O (g10257), .I (g10197));
INVX1 gate3478(.O (g4317), .I (I7586));
INVX1 gate3479(.O (g8278), .I (I13206));
INVX1 gate3480(.O (I4876), .I (g580));
INVX1 gate3481(.O (g3093), .I (I6299));
INVX1 gate3482(.O (g1998), .I (g802));
INVX1 gate3483(.O (g5474), .I (I8889));
INVX1 gate3484(.O (g10111), .I (I15347));
INVX1 gate3485(.O (g7192), .I (g6742));
INVX1 gate3486(.O (g5992), .I (I9608));
INVX1 gate3487(.O (g7085), .I (I11318));
INVX1 gate3488(.O (g3256), .I (I6424));
INVX1 gate3489(.O (I7746), .I (g3763));
INVX1 gate3490(.O (g6634), .I (I10589));
INVX1 gate3491(.O (I9188), .I (g4908));
INVX1 gate3492(.O (I10762), .I (g6127));
INVX1 gate3493(.O (g8667), .I (I13952));
INVX1 gate3494(.O (g3816), .I (g3228));
INVX1 gate3495(.O (g8143), .I (g8029));
INVX1 gate3496(.O (I13816), .I (g8559));
INVX1 gate3497(.O (I15548), .I (g10083));
INVX1 gate3498(.O (I6504), .I (g3214));
INVX1 gate3499(.O (I9388), .I (g5576));
INVX1 gate3500(.O (g8235), .I (g7967));
INVX1 gate3501(.O (g8343), .I (I13409));
INVX1 gate3502(.O (g6742), .I (g5830));
INVX1 gate3503(.O (g11548), .I (g11519));
INVX1 gate3504(.O (g6104), .I (I9769));
INVX1 gate3505(.O (I14964), .I (g9762));
INVX1 gate3506(.O (g10590), .I (I16255));
INVX1 gate3507(.O (I9216), .I (g4935));
INVX1 gate3508(.O (I6385), .I (g2260));
INVX1 gate3509(.O (g6304), .I (I10171));
INVX1 gate3510(.O (I16856), .I (g10909));
INVX1 gate3511(.O (g8566), .I (I13791));
INVX1 gate3512(.O (g6499), .I (g5867));
INVX1 gate3513(.O (I16261), .I (g10556));
INVX1 gate3514(.O (g2202), .I (g148));
INVX1 gate3515(.O (g11504), .I (I17531));
INVX1 gate3516(.O (g8988), .I (I14385));
INVX1 gate3517(.O (g4775), .I (I8139));
INVX1 gate3518(.O (I11752), .I (g7032));
INVX1 gate3519(.O (g8134), .I (I13005));
INVX1 gate3520(.O (g7941), .I (g7406));
INVX1 gate3521(.O (I15317), .I (g10025));
INVX1 gate3522(.O (I6025), .I (g2259));
INVX1 gate3523(.O (g2908), .I (I6077));
INVX1 gate3524(.O (g8334), .I (I13382));
INVX1 gate3525(.O (g9265), .I (g8892));
INVX1 gate3526(.O (g6926), .I (I11046));
INVX1 gate3527(.O (g2094), .I (I4924));
INVX1 gate3528(.O (I12415), .I (g7631));
INVX1 gate3529(.O (g11317), .I (I17112));
INVX1 gate3530(.O (g10094), .I (I15329));
INVX1 gate3531(.O (g3397), .I (g2896));
INVX1 gate3532(.O (g8548), .I (g8390));
INVX1 gate3533(.O (g2518), .I (g590));
INVX1 gate3534(.O (g4060), .I (g3144));
INVX1 gate3535(.O (g4460), .I (g3820));
INVX1 gate3536(.O (I9564), .I (g5109));
INVX1 gate3537(.O (I7468), .I (g3697));
INVX1 gate3538(.O (g6273), .I (I10078));
INVX1 gate3539(.O (I8885), .I (g4548));
INVX1 gate3540(.O (g8804), .I (I14133));
INVX1 gate3541(.O (I14543), .I (g9311));
INVX1 gate3542(.O (I8414), .I (g4293));
INVX1 gate3543(.O (g10150), .I (I15448));
INVX1 gate3544(.O (g10801), .I (I16507));
INVX1 gate3545(.O (I9826), .I (g5390));
INVX1 gate3546(.O (I10117), .I (g6241));
INVX1 gate3547(.O (g7708), .I (I12339));
INVX1 gate3548(.O (I13669), .I (g8294));
INVX1 gate3549(.O (g10735), .I (I16416));
INVX1 gate3550(.O (g10877), .I (I16601));
INVX1 gate3551(.O (g11057), .I (g10937));
INVX1 gate3552(.O (g7520), .I (I11898));
INVX1 gate3553(.O (g8792), .I (I14105));
INVX1 gate3554(.O (I17347), .I (g11373));
INVX1 gate3555(.O (I7677), .I (g3735));
INVX1 gate3556(.O (I11668), .I (g7043));
INVX1 gate3557(.O (g6044), .I (I9665));
INVX1 gate3558(.O (g2593), .I (g1973));
INVX1 gate3559(.O (g7031), .I (g6413));
INVX1 gate3560(.O (g4739), .I (g4117));
INVX1 gate3561(.O (I8903), .I (g4561));
INVX1 gate3562(.O (g6444), .I (g6158));
INVX1 gate3563(.O (g11245), .I (g11112));
INVX1 gate3564(.O (g7431), .I (I11821));
INVX1 gate3565(.O (I15323), .I (g10019));
INVX1 gate3566(.O (g6269), .I (I10066));
INVX1 gate3567(.O (I15299), .I (g9995));
INVX1 gate3568(.O (g7812), .I (I12601));
INVX1 gate3569(.O (g11626), .I (I17692));
INVX1 gate3570(.O (g9770), .I (g9432));
INVX1 gate3571(.O (g10196), .I (I15562));
INVX1 gate3572(.O (I11489), .I (g6569));
INVX1 gate3573(.O (g10695), .I (I16366));
INVX1 gate3574(.O (g5688), .I (I9213));
INVX1 gate3575(.O (g11323), .I (I17124));
INVX1 gate3576(.O (I13489), .I (g8233));
INVX1 gate3577(.O (g2965), .I (I6196));
INVX1 gate3578(.O (I6406), .I (g2339));
INVX1 gate3579(.O (I5475), .I (g1289));
INVX1 gate3580(.O (I7716), .I (g3751));
INVX1 gate3581(.O (g6572), .I (g5805));
INVX1 gate3582(.O (g6862), .I (g6720));
INVX1 gate3583(.O (g7376), .I (I11756));
INVX1 gate3584(.O (I5949), .I (g2540));
INVX1 gate3585(.O (g10526), .I (g10460));
INVX1 gate3586(.O (g8313), .I (I13323));
INVX1 gate3587(.O (I12484), .I (g7580));
INVX1 gate3588(.O (I14242), .I (g8787));
INVX1 gate3589(.O (I9108), .I (g5593));
INVX1 gate3590(.O (I15775), .I (g10253));
INVX1 gate3591(.O (I13424), .I (g8200));
INVX1 gate3592(.O (g4479), .I (I7858));
INVX1 gate3593(.O (g9532), .I (I14681));
INVX1 gate3594(.O (I9308), .I (g5494));
INVX1 gate3595(.O (g6712), .I (g5984));
INVX1 gate3596(.O (I8036), .I (g3820));
INVX1 gate3597(.O (g4294), .I (g3664));
INVX1 gate3598(.O (I10123), .I (g5676));
INVX1 gate3599(.O (g6543), .I (g5888));
INVX1 gate3600(.O (g4840), .I (I8199));
INVX1 gate3601(.O (I8436), .I (g4462));
INVX1 gate3602(.O (g9553), .I (I14694));
INVX1 gate3603(.O (I5292), .I (g76));
INVX1 gate3604(.O (I9883), .I (g5557));
INVX1 gate3605(.O (I14123), .I (g8767));
INVX1 gate3606(.O (g3723), .I (g3071));
INVX1 gate3607(.O (g7765), .I (I12460));
INVX1 gate3608(.O (g7286), .I (I11534));
INVX1 gate3609(.O (g4190), .I (I7387));
INVX1 gate3610(.O (I5998), .I (g2197));
INVX1 gate3611(.O (g4390), .I (g3914));
INVX1 gate3612(.O (I10807), .I (g6396));
INVX1 gate3613(.O (g10457), .I (I15962));
INVX1 gate3614(.O (g3817), .I (I7043));
INVX1 gate3615(.O (g7911), .I (g7664));
INVX1 gate3616(.O (I5646), .I (g940));
INVX1 gate3617(.O (I10974), .I (g6563));
INVX1 gate3618(.O (g8094), .I (g7987));
INVX1 gate3619(.O (g2050), .I (g1861));
INVX1 gate3620(.O (g2641), .I (g1987));
INVX1 gate3621(.O (I8831), .I (g4480));
INVX1 gate3622(.O (I15232), .I (g9974));
INVX1 gate3623(.O (I10639), .I (g5830));
INVX1 gate3624(.O (I17516), .I (g11483));
INVX1 gate3625(.O (g2450), .I (g1351));
INVX1 gate3626(.O (I16432), .I (g10702));
INVX1 gate3627(.O (g4501), .I (g3946));
INVX1 gate3628(.O (g8518), .I (I13723));
INVX1 gate3629(.O (g6729), .I (I10724));
INVX1 gate3630(.O (g6961), .I (I11115));
INVX1 gate3631(.O (g8567), .I (I13794));
INVX1 gate3632(.O (I10293), .I (g5863));
INVX1 gate3633(.O (g4156), .I (I7295));
INVX1 gate3634(.O (I11713), .I (g7023));
INVX1 gate3635(.O (g7733), .I (I12380));
INVX1 gate3636(.O (I5850), .I (g2273));
INVX1 gate3637(.O (g7270), .I (I11515));
INVX1 gate3638(.O (g9990), .I (I15190));
INVX1 gate3639(.O (g6927), .I (I11049));
INVX1 gate3640(.O (g3751), .I (I6944));
INVX1 gate3641(.O (I9165), .I (g5037));
INVX1 gate3642(.O (I16461), .I (g10735));
INVX1 gate3643(.O (I9571), .I (g5509));
INVX1 gate3644(.O (I9365), .I (g5392));
INVX1 gate3645(.O (g7610), .I (I12180));
INVX1 gate3646(.O (g2179), .I (g89));
INVX1 gate3647(.O (g4942), .I (I8308));
INVX1 gate3648(.O (g9029), .I (I14424));
INVX1 gate3649(.O (g6014), .I (g5309));
INVX1 gate3650(.O (g7073), .I (I11296));
INVX1 gate3651(.O (I12799), .I (g7556));
INVX1 gate3652(.O (g7796), .I (I12553));
INVX1 gate3653(.O (I12813), .I (g7688));
INVX1 gate3654(.O (g6885), .I (I10979));
INVX1 gate3655(.O (g9429), .I (g9082));
INVX1 gate3656(.O (g22), .I (I4777));
INVX1 gate3657(.O (g7473), .I (g7148));
INVX1 gate3658(.O (I10391), .I (g5838));
INVX1 gate3659(.O (I17209), .I (g11289));
INVX1 gate3660(.O (g6660), .I (I10623));
INVX1 gate3661(.O (I11255), .I (g6547));
INVX1 gate3662(.O (g10256), .I (g10140));
INVX1 gate3663(.O (I6173), .I (g2125));
INVX1 gate3664(.O (g11512), .I (I17555));
INVX1 gate3665(.O (I13255), .I (g8270));
INVX1 gate3666(.O (I14391), .I (g8928));
INVX1 gate3667(.O (I16650), .I (g10776));
INVX1 gate3668(.O (I6373), .I (g2024));
INVX1 gate3669(.O (I6091), .I (g2270));
INVX1 gate3670(.O (g5183), .I (g4640));
INVX1 gate3671(.O (g7124), .I (I11363));
INVX1 gate3672(.O (g7980), .I (I12786));
INVX1 gate3673(.O (g7324), .I (I11620));
INVX1 gate3674(.O (g10280), .I (g10160));
INVX1 gate3675(.O (g6903), .I (I11005));
INVX1 gate3676(.O (g2777), .I (g2276));
INVX1 gate3677(.O (I5919), .I (g2530));
INVX1 gate3678(.O (I11188), .I (g6513));
INVX1 gate3679(.O (g7069), .I (I11286));
INVX1 gate3680(.O (I12805), .I (g7684));
INVX1 gate3681(.O (I13188), .I (g8171));
INVX1 gate3682(.O (g5779), .I (I9371));
INVX1 gate3683(.O (I13678), .I (g8306));
INVX1 gate3684(.O (I14579), .I (g9272));
INVX1 gate3685(.O (g4954), .I (g4509));
INVX1 gate3686(.O (g4250), .I (g3698));
INVX1 gate3687(.O (g4163), .I (I7308));
INVX1 gate3688(.O (I5952), .I (g2506));
INVX1 gate3689(.O (g2882), .I (I6034));
INVX1 gate3690(.O (g7540), .I (I11956));
INVX1 gate3691(.O (g8160), .I (I13057));
INVX1 gate3692(.O (g4363), .I (I7654));
INVX1 gate3693(.O (I11686), .I (g7039));
INVX1 gate3694(.O (I16528), .I (g10732));
INVX1 gate3695(.O (I7577), .I (g4124));
INVX1 gate3696(.O (I5276), .I (g1411));
INVX1 gate3697(.O (g8360), .I (I13460));
INVX1 gate3698(.O (I16843), .I (g10898));
INVX1 gate3699(.O (I6007), .I (g2199));
INVX1 gate3700(.O (g5423), .I (g4300));
INVX1 gate3701(.O (I13460), .I (g8155));
INVX1 gate3702(.O (I17453), .I (g11451));
INVX1 gate3703(.O (I11383), .I (g6385));
INVX1 gate3704(.O (g2271), .I (g877));
INVX1 gate3705(.O (g7377), .I (I11759));
INVX1 gate3706(.O (g7206), .I (I11436));
INVX1 gate3707(.O (g10157), .I (I15467));
INVX1 gate3708(.O (g11445), .I (I17384));
INVX1 gate3709(.O (g6036), .I (I9647));
INVX1 gate3710(.O (I5561), .I (g869));
INVX1 gate3711(.O (I13030), .I (g8052));
INVX1 gate3712(.O (g2611), .I (I5734));
INVX1 gate3713(.O (g4453), .I (I7810));
INVX1 gate3714(.O (g8450), .I (I13648));
INVX1 gate3715(.O (g6178), .I (g4977));
INVX1 gate3716(.O (I6767), .I (g2914));
INVX1 gate3717(.O (g11499), .I (I17516));
INVX1 gate3718(.O (I8495), .I (g4325));
INVX1 gate3719(.O (g3368), .I (g3138));
INVX1 gate3720(.O (g9745), .I (g9454));
INVX1 gate3721(.O (I11065), .I (g6750));
INVX1 gate3722(.O (I6535), .I (g2826));
INVX1 gate3723(.O (g1987), .I (g762));
INVX1 gate3724(.O (g9338), .I (I14519));
INVX1 gate3725(.O (g7287), .I (I11537));
INVX1 gate3726(.O (g2799), .I (g2276));
INVX1 gate3727(.O (g11498), .I (I17513));
INVX1 gate3728(.O (I5986), .I (g2194));
INVX1 gate3729(.O (g6135), .I (I9842));
INVX1 gate3730(.O (g5665), .I (I9156));
INVX1 gate3731(.O (g9109), .I (I14452));
INVX1 gate3732(.O (g6335), .I (I10228));
INVX1 gate3733(.O (I15989), .I (g10417));
INVX1 gate3734(.O (g9309), .I (g8892));
INVX1 gate3735(.O (g3531), .I (g2971));
INVX1 gate3736(.O (I8869), .I (g4421));
INVX1 gate3737(.O (g5127), .I (I8535));
INVX1 gate3738(.O (g3458), .I (g3144));
INVX1 gate3739(.O (g6182), .I (g5446));
INVX1 gate3740(.O (g6288), .I (I10123));
INVX1 gate3741(.O (I17274), .I (g11389));
INVX1 gate3742(.O (g6382), .I (I10278));
INVX1 gate3743(.O (I9662), .I (g5319));
INVX1 gate3744(.O (g8179), .I (I13086));
INVX1 gate3745(.O (g7849), .I (I12644));
INVX1 gate3746(.O (g10876), .I (I16598));
INVX1 gate3747(.O (g10885), .I (g10809));
INVX1 gate3748(.O (g11056), .I (g10950));
INVX1 gate3749(.O (g3743), .I (I6932));
INVX1 gate3750(.O (g8379), .I (I13485));
INVX1 gate3751(.O (g4912), .I (I8282));
INVX1 gate3752(.O (I14116), .I (g8766));
INVX1 gate3753(.O (g2997), .I (g2135));
INVX1 gate3754(.O (g11611), .I (I17657));
INVX1 gate3755(.O (I12400), .I (g7537));
INVX1 gate3756(.O (g2541), .I (I5658));
INVX1 gate3757(.O (g11080), .I (I16853));
INVX1 gate3758(.O (I7426), .I (g3334));
INVX1 gate3759(.O (I9290), .I (g5052));
INVX1 gate3760(.O (g5146), .I (g4596));
INVX1 gate3761(.O (g10854), .I (g10708));
INVX1 gate3762(.O (g6805), .I (I10825));
INVX1 gate3763(.O (g5633), .I (g4388));
INVX1 gate3764(.O (g3505), .I (I6694));
INVX1 gate3765(.O (g7781), .I (I12508));
INVX1 gate3766(.O (I5970), .I (g2185));
INVX1 gate3767(.O (g6749), .I (I10756));
INVX1 gate3768(.O (I16708), .I (g10822));
INVX1 gate3769(.O (g2238), .I (I5237));
INVX1 gate3770(.O (g11432), .I (I17347));
INVX1 gate3771(.O (I13837), .I (g8488));
INVX1 gate3772(.O (g3411), .I (I6616));
INVX1 gate3773(.O (I9093), .I (g5397));
INVX1 gate3774(.O (g7900), .I (g7712));
INVX1 gate3775(.O (I16258), .I (g10555));
INVX1 gate3776(.O (I4948), .I (g586));
INVX1 gate3777(.O (g2209), .I (g93));
INVX1 gate3778(.O (g7797), .I (I12556));
INVX1 gate3779(.O (I9256), .I (g5078));
INVX1 gate3780(.O (I8265), .I (g4602));
INVX1 gate3781(.O (I9816), .I (g5576));
INVX1 gate3782(.O (g5696), .I (I9229));
INVX1 gate3783(.O (I15461), .I (g10074));
INVX1 gate3784(.O (g6947), .I (I11085));
INVX1 gate3785(.O (I7984), .I (g3621));
INVX1 gate3786(.O (I5224), .I (g61));
INVX1 gate3787(.O (I7280), .I (g3208));
INVX1 gate3788(.O (I10237), .I (g6120));
INVX1 gate3789(.O (g6798), .I (I10804));
INVX1 gate3790(.O (I8442), .I (g4464));
INVX1 gate3791(.O (I12538), .I (g7658));
INVX1 gate3792(.O (g8271), .I (I13185));
INVX1 gate3793(.O (g2802), .I (g2276));
INVX1 gate3794(.O (g11342), .I (I17149));
INVX1 gate3795(.O (I10340), .I (g6205));
INVX1 gate3796(.O (g1991), .I (g778));
INVX1 gate3797(.O (I5120), .I (g622));
INVX1 gate3798(.O (g3474), .I (I6679));
INVX1 gate3799(.O (g9449), .I (g9094));
INVX1 gate3800(.O (g6560), .I (g5759));
INVX1 gate3801(.O (I14340), .I (g8820));
INVX1 gate3802(.O (g5753), .I (I9329));
INVX1 gate3803(.O (I8164), .I (g3566));
INVX1 gate3804(.O (I15736), .I (g10258));
INVX1 gate3805(.O (g10456), .I (I15959));
INVX1 gate3806(.O (g5508), .I (I8929));
INVX1 gate3807(.O (g11199), .I (g11112));
INVX1 gate3808(.O (I14684), .I (g9124));
INVX1 gate3809(.O (g11650), .I (I17752));
INVX1 gate3810(.O (g7144), .I (I11387));
INVX1 gate3811(.O (I11617), .I (g6839));
INVX1 gate3812(.O (g7344), .I (I11680));
INVX1 gate3813(.O (g5072), .I (I8442));
INVX1 gate3814(.O (I7636), .I (g3330));
INVX1 gate3815(.O (I13915), .I (g8451));
INVX1 gate3816(.O (g5472), .I (I8885));
INVX1 gate3817(.O (g8981), .I (I14364));
INVX1 gate3818(.O (I9421), .I (g5063));
INVX1 gate3819(.O (g8674), .I (I13959));
INVX1 gate3820(.O (I5789), .I (g2162));
INVX1 gate3821(.O (g5043), .I (g4840));
INVX1 gate3822(.O (I11201), .I (g6522));
INVX1 gate3823(.O (g10314), .I (I15744));
INVX1 gate3824(.O (g7259), .I (I11494));
INVX1 gate3825(.O (g5443), .I (I8872));
INVX1 gate3826(.O (g6208), .I (I9953));
INVX1 gate3827(.O (I7790), .I (g3782));
INVX1 gate3828(.O (I16879), .I (g10936));
INVX1 gate3829(.O (g6302), .I (I10165));
INVX1 gate3830(.O (g10307), .I (I15729));
INVX1 gate3831(.O (I15365), .I (g10025));
INVX1 gate3832(.O (I7061), .I (g3050));
INVX1 gate3833(.O (g6579), .I (g5949));
INVX1 gate3834(.O (g5116), .I (g4682));
INVX1 gate3835(.O (g6869), .I (I10949));
INVX1 gate3836(.O (g7852), .I (g7479));
INVX1 gate3837(.O (g7923), .I (g7527));
INVX1 gate3838(.O (I17164), .I (g11320));
INVX1 gate3839(.O (I7387), .I (g4083));
INVX1 gate3840(.O (g10596), .I (I16269));
INVX1 gate3841(.O (I11467), .I (g6488));
INVX1 gate3842(.O (I11494), .I (g6574));
INVX1 gate3843(.O (I13595), .I (g8339));
INVX1 gate3844(.O (g8132), .I (I12999));
INVX1 gate3845(.O (g6719), .I (I10710));
INVX1 gate3846(.O (I12235), .I (g7082));
INVX1 gate3847(.O (g8332), .I (I13376));
INVX1 gate3848(.O (g10243), .I (I15635));
INVX1 gate3849(.O (I11623), .I (g6841));
INVX1 gate3850(.O (I12683), .I (g7387));
INVX1 gate3851(.O (I6388), .I (g2329));
INVX1 gate3852(.O (g8680), .I (I13965));
INVX1 gate3853(.O (g10431), .I (g10328));
INVX1 gate3854(.O (I11037), .I (g6629));
INVX1 gate3855(.O (g8353), .I (I13439));
INVX1 gate3856(.O (I14130), .I (g8769));
INVX1 gate3857(.O (I10362), .I (g6224));
INVX1 gate3858(.O (g2864), .I (g2298));
INVX1 gate3859(.O (I10165), .I (g5948));
INVX1 gate3860(.O (I13782), .I (g8515));
INVX1 gate3861(.O (g6917), .I (I11029));
INVX1 gate3862(.O (g4894), .I (I8247));
INVX1 gate3863(.O (I6028), .I (g2208));
INVX1 gate3864(.O (g10269), .I (g10154));
INVX1 gate3865(.O (g8802), .I (I14127));
INVX1 gate3866(.O (I6671), .I (g2757));
INVX1 gate3867(.O (I6428), .I (g2348));
INVX1 gate3868(.O (g7886), .I (g7479));
INVX1 gate3869(.O (g4735), .I (g3546));
INVX1 gate3870(.O (I17327), .I (g11349));
INVX1 gate3871(.O (g6265), .I (I10054));
INVX1 gate3872(.O (g3976), .I (I7109));
INVX1 gate3873(.O (I6247), .I (g2462));
INVX1 gate3874(.O (g4782), .I (g4089));
INVX1 gate3875(.O (I11155), .I (g6470));
INVX1 gate3876(.O (g10156), .I (I15464));
INVX1 gate3877(.O (I15708), .I (g10241));
INVX1 gate3878(.O (I17537), .I (g11497));
INVX1 gate3879(.O (I13418), .I (g8145));
INVX1 gate3880(.O (I13822), .I (g8488));
INVX1 gate3881(.O (g5697), .I (I9232));
INVX1 gate3882(.O (I10006), .I (g5633));
INVX1 gate3883(.O (g6442), .I (I10362));
INVX1 gate3884(.O (g9452), .I (I14645));
INVX1 gate3885(.O (g7314), .I (I11590));
INVX1 gate3886(.O (g5210), .I (I8631));
INVX1 gate3887(.O (I17108), .I (g11225));
INVX1 gate3888(.O (g11471), .I (I17450));
INVX1 gate3889(.O (I7345), .I (g4050));
INVX1 gate3890(.O (I16458), .I (g10734));
INVX1 gate3891(.O (I8429), .I (g4458));
INVX1 gate3892(.O (I9605), .I (g5620));
INVX1 gate3893(.O (g4475), .I (I7852));
INVX1 gate3894(.O (g5596), .I (I9020));
INVX1 gate3895(.O (g6164), .I (g5426));
INVX1 gate3896(.O (I7763), .I (g3769));
INVX1 gate3897(.O (I7191), .I (g2646));
INVX1 gate3898(.O (g10734), .I (I16413));
INVX1 gate3899(.O (I10437), .I (g5755));
INVX1 gate3900(.O (g10335), .I (I15787));
INVX1 gate3901(.O (g7650), .I (I12261));
INVX1 gate3902(.O (g3326), .I (I6495));
INVX1 gate3903(.O (I15244), .I (g10031));
INVX1 gate3904(.O (g4292), .I (g3863));
INVX1 gate3905(.O (g10930), .I (g10827));
INVX1 gate3906(.O (g11043), .I (I16790));
INVX1 gate3907(.O (g6454), .I (I10388));
INVX1 gate3908(.O (g11244), .I (g11112));
INVX1 gate3909(.O (g4526), .I (I7931));
INVX1 gate3910(.O (I5478), .I (g1212));
INVX1 gate3911(.O (g6296), .I (I10147));
INVX1 gate3912(.O (I11194), .I (g6515));
INVX1 gate3913(.O (g3760), .I (g3003));
INVX1 gate3914(.O (g7008), .I (I11149));
INVX1 gate3915(.O (I13194), .I (g8140));
INVX1 gate3916(.O (I13589), .I (g8361));
INVX1 gate3917(.O (g2623), .I (g1999));
INVX1 gate3918(.O (I17381), .I (g11436));
INVX1 gate3919(.O (I7536), .I (g4098));
INVX1 gate3920(.O (I9585), .I (g5241));
INVX1 gate3921(.O (g2076), .I (I4886));
INVX1 gate3922(.O (g10131), .I (I15395));
INVX1 gate3923(.O (g2889), .I (I6049));
INVX1 gate3924(.O (I11524), .I (g6593));
INVX1 gate3925(.O (I16598), .I (g10804));
INVX1 gate3926(.O (g11069), .I (g10974));
INVX1 gate3927(.O (g4084), .I (g3119));
INVX1 gate3928(.O (I11836), .I (g7220));
INVX1 gate3929(.O (I5435), .I (g18));
INVX1 gate3930(.O (g4603), .I (g3829));
INVX1 gate3931(.O (g5936), .I (I9564));
INVX1 gate3932(.O (g7336), .I (I11656));
INVX1 gate3933(.O (g8600), .I (g8475));
INVX1 gate3934(.O (I15068), .I (g9710));
INVX1 gate3935(.O (g7768), .I (I12469));
INVX1 gate3936(.O (g4439), .I (I7793));
INVX1 gate3937(.O (g11657), .I (I17773));
INVX1 gate3938(.O (g5117), .I (g4682));
INVX1 gate3939(.O (g6553), .I (I10477));
INVX1 gate3940(.O (g8714), .I (I14005));
INVX1 gate3941(.O (g11068), .I (g10974));
INVX1 gate3942(.O (I7858), .I (g3631));
INVX1 gate3943(.O (I11477), .I (g6488));
INVX1 gate3944(.O (g7594), .I (I12120));
INVX1 gate3945(.O (g10487), .I (I16098));
INVX1 gate3946(.O (g7972), .I (I12770));
INVX1 gate3947(.O (g2175), .I (g44));
INVX1 gate3948(.O (I11119), .I (g6461));
INVX1 gate3949(.O (g9025), .I (I14412));
INVX1 gate3950(.O (g2871), .I (I6013));
INVX1 gate3951(.O (g10619), .I (I16292));
INVX1 gate3952(.O (I12759), .I (g7702));
INVX1 gate3953(.O (I7757), .I (g3767));
INVX1 gate3954(.O (I16817), .I (g10912));
INVX1 gate3955(.O (I9673), .I (g5182));
INVX1 gate3956(.O (I14236), .I (g8802));
INVX1 gate3957(.O (g7806), .I (I12583));
INVX1 gate3958(.O (I10952), .I (g6556));
INVX1 gate3959(.O (g3220), .I (I6398));
INVX1 gate3960(.O (I8109), .I (g3622));
INVX1 gate3961(.O (g2651), .I (g2007));
INVX1 gate3962(.O (I6217), .I (g2302));
INVX1 gate3963(.O (g4583), .I (g3880));
INVX1 gate3964(.O (g6412), .I (I10322));
INVX1 gate3965(.O (I17390), .I (g11430));
INVX1 gate3966(.O (g10279), .I (g10158));
INVX1 gate3967(.O (g7065), .I (I11272));
INVX1 gate3968(.O (I7315), .I (g2891));
INVX1 gate3969(.O (g6389), .I (I10289));
INVX1 gate3970(.O (I7642), .I (g3440));
INVX1 gate3971(.O (I9168), .I (g5040));
INVX1 gate3972(.O (g6706), .I (I10685));
INVX1 gate3973(.O (I9669), .I (g5426));
INVX1 gate3974(.O (g7887), .I (g7693));
INVX1 gate3975(.O (g7122), .I (I11357));
INVX1 gate3976(.O (I15792), .I (g10279));
INVX1 gate3977(.O (I9368), .I (g5288));
INVX1 gate3978(.O (g7322), .I (I11614));
INVX1 gate3979(.O (g4919), .I (I8290));
INVX1 gate3980(.O (I10063), .I (g5766));
INVX1 gate3981(.O (g6990), .I (I11132));
INVX1 gate3982(.O (I7447), .I (g3694));
INVX1 gate3983(.O (g10278), .I (g10182));
INVX1 gate3984(.O (g3977), .I (I7112));
INVX1 gate3985(.O (I6861), .I (g2942));
INVX1 gate3986(.O (g6888), .I (I10984));
INVX1 gate3987(.O (I16656), .I (g10791));
INVX1 gate3988(.O (I9531), .I (g5004));
INVX1 gate3989(.O (g6171), .I (g5446));
INVX1 gate3990(.O (g2184), .I (g1806));
INVX1 gate3991(.O (I16295), .I (g10552));
INVX1 gate3992(.O (I9458), .I (g5091));
INVX1 gate3993(.O (g3161), .I (I6367));
INVX1 gate3994(.O (I11704), .I (g7008));
INVX1 gate3995(.O (I12849), .I (g7632));
INVX1 gate3996(.O (I6055), .I (g2569));
INVX1 gate3997(.O (I17522), .I (g11485));
INVX1 gate3998(.O (g2339), .I (I5399));
INVX1 gate3999(.O (g7033), .I (I11188));
INVX1 gate4000(.O (g10039), .I (I15244));
INVX1 gate4001(.O (I10873), .I (g6331));
INVX1 gate4002(.O (g6956), .I (I11106));
INVX1 gate4003(.O (g5597), .I (I9023));
INVX1 gate4004(.O (I14873), .I (g9525));
INVX1 gate4005(.O (I7654), .I (g3728));
INVX1 gate4006(.O (I13809), .I (g8480));
INVX1 gate4007(.O (I6133), .I (g2253));
INVX1 gate4008(.O (g3051), .I (g2135));
INVX1 gate4009(.O (g2838), .I (g2165));
INVX1 gate4010(.O (g8076), .I (I12930));
INVX1 gate4011(.O (g2024), .I (g1718));
INVX1 gate4012(.O (I15458), .I (g10069));
INVX1 gate4013(.O (I13466), .I (g8160));
INVX1 gate4014(.O (I9505), .I (g5088));
INVX1 gate4015(.O (g6281), .I (I10102));
INVX1 gate4016(.O (g8476), .I (I13674));
INVX1 gate4017(.O (g3327), .I (I6498));
INVX1 gate4018(.O (g2424), .I (g1690));
INVX1 gate4019(.O (I8449), .I (g4469));
INVX1 gate4020(.O (I12652), .I (g7458));
INVX1 gate4021(.O (g9766), .I (g9432));
INVX1 gate4022(.O (g2809), .I (I5909));
INVX1 gate4023(.O (g5784), .I (I9380));
INVX1 gate4024(.O (g4004), .I (I7140));
INVX1 gate4025(.O (I9734), .I (g5257));
INVX1 gate4026(.O (I13036), .I (g8053));
INVX1 gate4027(.O (I5002), .I (g1173));
INVX1 gate4028(.O (I8865), .I (g4518));
INVX1 gate4029(.O (g7550), .I (g6974));
INVX1 gate4030(.O (g6297), .I (I10150));
INVX1 gate4031(.O (I11560), .I (g7037));
INVX1 gate4032(.O (g10187), .I (I15539));
INVX1 gate4033(.O (I6196), .I (g2462));
INVX1 gate4034(.O (I5824), .I (g2502));
INVX1 gate4035(.O (g7845), .I (I12634));
INVX1 gate4036(.O (I10834), .I (g6715));
INVX1 gate4037(.O (g8871), .I (I14185));
INVX1 gate4038(.O (g8375), .I (I13475));
INVX1 gate4039(.O (I15545), .I (g10075));
INVX1 gate4040(.O (g3633), .I (I6802));
INVX1 gate4041(.O (I15079), .I (g9745));
INVX1 gate4042(.O (I8098), .I (g3583));
INVX1 gate4043(.O (g2077), .I (g219));
INVX1 gate4044(.O (g2231), .I (I5218));
INVX1 gate4045(.O (g7195), .I (I11417));
INVX1 gate4046(.O (g11545), .I (g11519));
INVX1 gate4047(.O (g11079), .I (I16850));
INVX1 gate4048(.O (g11444), .I (I17381));
INVX1 gate4049(.O (g5937), .I (I9567));
INVX1 gate4050(.O (g7395), .I (g6941));
INVX1 gate4051(.O (I13642), .I (g8378));
INVX1 gate4052(.O (g7337), .I (I11659));
INVX1 gate4053(.O (g3103), .I (g2391));
INVX1 gate4054(.O (I9074), .I (g4764));
INVX1 gate4055(.O (g7913), .I (g7467));
INVX1 gate4056(.O (I6538), .I (g2827));
INVX1 gate4057(.O (g2523), .I (I5632));
INVX1 gate4058(.O (I7272), .I (g3253));
INVX1 gate4059(.O (g2643), .I (g1989));
INVX1 gate4060(.O (I9992), .I (g5633));
INVX1 gate4061(.O (g10143), .I (I15427));
INVX1 gate4062(.O (g5668), .I (I9165));
INVX1 gate4063(.O (g11078), .I (I16847));
INVX1 gate4064(.O (g6338), .I (I10237));
INVX1 gate4065(.O (I15598), .I (g10170));
INVX1 gate4066(.O (I10021), .I (g5692));
INVX1 gate4067(.O (g5840), .I (g5320));
INVX1 gate4068(.O (g4970), .I (g4411));
INVX1 gate4069(.O (g8500), .I (I13695));
INVX1 gate4070(.O (I7612), .I (g3817));
INVX1 gate4071(.O (g11598), .I (I17642));
INVX1 gate4072(.O (I7017), .I (g3068));
INVX1 gate4073(.O (g6109), .I (g5052));
INVX1 gate4074(.O (I12406), .I (g7464));
INVX1 gate4075(.O (g6309), .I (I10186));
INVX1 gate4076(.O (g11086), .I (I16867));
INVX1 gate4077(.O (g7807), .I (I12586));
INVX1 gate4078(.O (I7417), .I (g4160));
INVX1 gate4079(.O (g3732), .I (I6914));
INVX1 gate4080(.O (I17252), .I (g11343));
INVX1 gate4081(.O (g10169), .I (I15503));
INVX1 gate4082(.O (I7935), .I (g3440));
INVX1 gate4083(.O (I9080), .I (g4775));
INVX1 gate4084(.O (g8184), .I (I13105));
INVX1 gate4085(.O (g10884), .I (g10809));
INVX1 gate4086(.O (g6808), .I (I10834));
INVX1 gate4087(.O (I15817), .I (g10199));
INVX1 gate4088(.O (I9863), .I (g5557));
INVX1 gate4089(.O (g8139), .I (g8025));
INVX1 gate4090(.O (I16289), .I (g10541));
INVX1 gate4091(.O (g8339), .I (I13397));
INVX1 gate4092(.O (g2742), .I (I5798));
INVX1 gate4093(.O (g3944), .I (g2920));
INVX1 gate4094(.O (g10168), .I (I15500));
INVX1 gate4095(.O (I10607), .I (g5763));
INVX1 gate4096(.O (g6707), .I (g5949));
INVX1 gate4097(.O (I13630), .I (g8334));
INVX1 gate4098(.O (g2304), .I (I5348));
INVX1 gate4099(.O (g11322), .I (I17121));
INVX1 gate4100(.O (g9091), .I (g8892));
INVX1 gate4101(.O (g4320), .I (g4013));
INVX1 gate4102(.O (I15977), .I (g10411));
INVX1 gate4103(.O (g11159), .I (g10950));
INVX1 gate4104(.O (I10274), .I (g5811));
INVX1 gate4105(.O (I11166), .I (g6480));
INVX1 gate4106(.O (I11665), .I (g7038));
INVX1 gate4107(.O (I16571), .I (g10819));
INVX1 gate4108(.O (I13166), .I (g8009));
INVX1 gate4109(.O (I7330), .I (g3761));
INVX1 gate4110(.O (I8268), .I (g4674));
INVX1 gate4111(.O (g8424), .I (I13586));
INVX1 gate4112(.O (I5064), .I (g1690));
INVX1 gate4113(.O (g8795), .I (I14112));
INVX1 gate4114(.O (g10217), .I (I15589));
INVX1 gate4115(.O (g7142), .I (I11383));
INVX1 gate4116(.O (I6256), .I (g2462));
INVX1 gate4117(.O (g4277), .I (g3688));
INVX1 gate4118(.O (g6201), .I (I9938));
INVX1 gate4119(.O (g7342), .I (I11674));
INVX1 gate4120(.O (I11008), .I (g6795));
INVX1 gate4121(.O (g6957), .I (I11109));
INVX1 gate4122(.O (I15353), .I (g10007));
INVX1 gate4123(.O (g2754), .I (I5830));
INVX1 gate4124(.O (g4906), .I (I8275));
INVX1 gate4125(.O (g7815), .I (I12610));
INVX1 gate4126(.O (g11656), .I (I17770));
INVX1 gate4127(.O (g4789), .I (g3337));
INVX1 gate4128(.O (I7800), .I (g3791));
INVX1 gate4129(.O (g10486), .I (I16095));
INVX1 gate4130(.O (g11353), .I (I17176));
INVX1 gate4131(.O (g8077), .I (I12933));
INVX1 gate4132(.O (I15823), .I (g10201));
INVX1 gate4133(.O (g6449), .I (g6172));
INVX1 gate4134(.O (I13485), .I (g8194));
INVX1 gate4135(.O (g2273), .I (g881));
INVX1 gate4136(.O (g8477), .I (g8317));
INVX1 gate4137(.O (g6575), .I (g5949));
INVX1 gate4138(.O (g7692), .I (g7148));
INVX1 gate4139(.O (I12613), .I (g7525));
INVX1 gate4140(.O (g8523), .I (I13732));
INVX1 gate4141(.O (I6381), .I (g2257));
INVX1 gate4142(.O (g9767), .I (I14914));
INVX1 gate4143(.O (g7097), .I (I11330));
INVX1 gate4144(.O (I9688), .I (g5201));
INVX1 gate4145(.O (g7726), .I (I12363));
INVX1 gate4146(.O (I9857), .I (g5269));
INVX1 gate4147(.O (I13454), .I (g8183));
INVX1 gate4148(.O (g2613), .I (I5740));
INVX1 gate4149(.O (g7497), .I (g7148));
INVX1 gate4150(.O (g9535), .I (I14690));
INVX1 gate4151(.O (g6715), .I (I10702));
INVX1 gate4152(.O (g2044), .I (I4850));
INVX1 gate4153(.O (g7354), .I (I11710));
INVX1 gate4154(.O (g10580), .I (g10530));
INVX1 gate4155(.O (I10153), .I (g5947));
INVX1 gate4156(.O (g2444), .I (g876));
INVX1 gate4157(.O (I5237), .I (g1107));
INVX1 gate4158(.O (g5032), .I (I8403));
INVX1 gate4159(.O (g2269), .I (I5308));
INVX1 gate4160(.O (g10223), .I (I15595));
INVX1 gate4161(.O (I7213), .I (g2635));
INVX1 gate4162(.O (g9261), .I (g8892));
INVX1 gate4163(.O (I6421), .I (g2346));
INVX1 gate4164(.O (g4299), .I (g4144));
INVX1 gate4165(.O (I14409), .I (g8938));
INVX1 gate4166(.O (I12463), .I (g7579));
INVX1 gate4167(.O (g3697), .I (I6856));
INVX1 gate4168(.O (g8099), .I (g7990));
INVX1 gate4169(.O (I8385), .I (g4238));
INVX1 gate4170(.O (I14136), .I (g8775));
INVX1 gate4171(.O (g8304), .I (I13280));
INVX1 gate4172(.O (g3914), .I (g3015));
INVX1 gate4173(.O (I9126), .I (g4891));
INVX1 gate4174(.O (I13239), .I (g8266));
INVX1 gate4175(.O (g10110), .I (I15344));
INVX1 gate4176(.O (g11631), .I (I17707));
INVX1 gate4177(.O (I9326), .I (g5320));
INVX1 gate4178(.O (g2543), .I (I5662));
INVX1 gate4179(.O (g6584), .I (I10538));
INVX1 gate4180(.O (g11017), .I (I16742));
INVX1 gate4181(.O (g6539), .I (I10461));
INVX1 gate4182(.O (g6896), .I (I10996));
INVX1 gate4183(.O (g5568), .I (I8985));
INVX1 gate4184(.O (g10321), .I (I15759));
INVX1 gate4185(.O (I5089), .I (g1854));
INVX1 gate4186(.O (I5731), .I (g2089));
INVX1 gate4187(.O (I11238), .I (g6543));
INVX1 gate4188(.O (I17213), .I (g11290));
INVX1 gate4189(.O (g7783), .I (I12514));
INVX1 gate4190(.O (g10179), .I (g10041));
INVX1 gate4191(.O (g10531), .I (g10471));
INVX1 gate4192(.O (g7979), .I (I12783));
INVX1 gate4193(.O (g3413), .I (g2896));
INVX1 gate4194(.O (g5912), .I (I9544));
INVX1 gate4195(.O (g7312), .I (I11584));
INVX1 gate4196(.O (I7166), .I (g2620));
INVX1 gate4197(.O (I5966), .I (g2541));
INVX1 gate4198(.O (g10178), .I (I15526));
INVX1 gate4199(.O (I7366), .I (g4012));
INVX1 gate4200(.O (g4738), .I (g3440));
INVX1 gate4201(.O (I13941), .I (g8488));
INVX1 gate4202(.O (I13382), .I (g8134));
INVX1 gate4203(.O (g6268), .I (I10063));
INVX1 gate4204(.O (I11519), .I (g6591));
INVX1 gate4205(.O (I11176), .I (g6501));
INVX1 gate4206(.O (g10186), .I (I15536));
INVX1 gate4207(.O (g7001), .I (I11140));
INVX1 gate4208(.O (g8273), .I (I13191));
INVX1 gate4209(.O (g10676), .I (g10570));
INVX1 gate4210(.O (g6419), .I (I10331));
INVX1 gate4211(.O (I10891), .I (g6334));
INVX1 gate4212(.O (I13185), .I (g8192));
INVX1 gate4213(.O (g11289), .I (I17070));
INVX1 gate4214(.O (I7456), .I (g3716));
INVX1 gate4215(.O (g1993), .I (g786));
INVX1 gate4216(.O (g3820), .I (I7048));
INVX1 gate4217(.O (g7676), .I (I12303));
INVX1 gate4218(.O (g4140), .I (I7284));
INVX1 gate4219(.O (g6052), .I (g5426));
INVX1 gate4220(.O (g11309), .I (I17096));
INVX1 gate4221(.O (g4078), .I (I7205));
INVX1 gate4222(.O (I12514), .I (g7735));
INVX1 gate4223(.O (g8613), .I (g8484));
INVX1 gate4224(.O (I16525), .I (g10719));
INVX1 gate4225(.O (I7348), .I (g4056));
INVX1 gate4226(.O (g6452), .I (I10384));
INVX1 gate4227(.O (I9383), .I (g5296));
INVX1 gate4228(.O (I9608), .I (g5127));
INVX1 gate4229(.O (I15308), .I (g10019));
INVX1 gate4230(.O (g7329), .I (I11635));
INVX1 gate4231(.O (g4478), .I (g3820));
INVX1 gate4232(.O (g7761), .I (I12448));
INVX1 gate4233(.O (g2014), .I (g1104));
INVX1 gate4234(.O (g4907), .I (I8278));
INVX1 gate4235(.O (g8444), .I (I13630));
INVX1 gate4236(.O (g2885), .I (I6043));
INVX1 gate4237(.O (I9779), .I (g5391));
INVX1 gate4238(.O (g2946), .I (I6133));
INVX1 gate4239(.O (g4435), .I (g3914));
INVX1 gate4240(.O (I9023), .I (g4727));
INVX1 gate4241(.O (g8983), .I (I14370));
INVX1 gate4242(.O (g4082), .I (I7213));
INVX1 gate4243(.O (I12421), .I (g7634));
INVX1 gate4244(.O (I8406), .I (g4274));
INVX1 gate4245(.O (I5254), .I (g1700));
INVX1 gate4246(.O (I14109), .I (g8765));
INVX1 gate4247(.O (g8572), .I (I13809));
INVX1 gate4248(.O (g7727), .I (I12366));
INVX1 gate4249(.O (I7964), .I (g3433));
INVX1 gate4250(.O (g2903), .I (g2166));
INVX1 gate4251(.O (I7260), .I (g2844));
INVX1 gate4252(.O (I14537), .I (g9308));
INVX1 gate4253(.O (I10108), .I (g5743));
INVX1 gate4254(.O (g6086), .I (I9737));
INVX1 gate4255(.O (g8712), .I (g8680));
INVX1 gate4256(.O (g11495), .I (I17500));
INVX1 gate4257(.O (I12012), .I (g6916));
INVX1 gate4258(.O (I9588), .I (g5114));
INVX1 gate4259(.O (g7746), .I (I12403));
INVX1 gate4260(.O (I8487), .I (g4526));
INVX1 gate4261(.O (I5438), .I (g18));
INVX1 gate4262(.O (g3775), .I (I7002));
INVX1 gate4263(.O (g7221), .I (I11459));
INVX1 gate4264(.O (I17350), .I (g11377));
INVX1 gate4265(.O (I14303), .I (g8811));
INVX1 gate4266(.O (g6385), .I (g6119));
INVX1 gate4267(.O (g6881), .I (I10971));
INVX1 gate4268(.O (I12541), .I (g7662));
INVX1 gate4269(.O (g7703), .I (g7085));
INVX1 gate4270(.O (I9665), .I (g5174));
INVX1 gate4271(.O (I15752), .I (g10264));
INVX1 gate4272(.O (g4915), .I (g4413));
INVX1 gate4273(.O (g2178), .I (g45));
INVX1 gate4274(.O (g2436), .I (I5525));
INVX1 gate4275(.O (I15374), .I (g10007));
INVX1 gate4276(.O (g9028), .I (I14421));
INVX1 gate4277(.O (g8729), .I (g8595));
INVX1 gate4278(.O (g8961), .I (I14330));
INVX1 gate4279(.O (I4900), .I (g583));
INVX1 gate4280(.O (I11501), .I (g6581));
INVX1 gate4281(.O (I16610), .I (g10792));
INVX1 gate4282(.O (g9671), .I (I14802));
INVX1 gate4283(.O (I17152), .I (g11308));
INVX1 gate4284(.O (g3060), .I (g2135));
INVX1 gate4285(.O (I13729), .I (g8290));
INVX1 gate4286(.O (I13577), .I (g8330));
INVX1 gate4287(.O (I10381), .I (g5847));
INVX1 gate4288(.O (g4214), .I (I7459));
INVX1 gate4289(.O (I16255), .I (g10554));
INVX1 gate4290(.O (I14982), .I (g9672));
INVX1 gate4291(.O (g6425), .I (g6141));
INVX1 gate4292(.O (I11728), .I (g7010));
INVX1 gate4293(.O (g11643), .I (I17733));
INVX1 gate4294(.O (g2135), .I (I5064));
INVX1 gate4295(.O (I16679), .I (g10784));
INVX1 gate4296(.O (g2335), .I (I5391));
INVX1 gate4297(.O (g5683), .I (I9202));
INVX1 gate4298(.O (I13439), .I (g8187));
INVX1 gate4299(.O (I9346), .I (g5281));
INVX1 gate4300(.O (I7118), .I (g2979));
INVX1 gate4301(.O (g4310), .I (I7577));
INVX1 gate4302(.O (g2382), .I (g599));
INVX1 gate4303(.O (I7318), .I (g3266));
INVX1 gate4304(.O (I12829), .I (g7680));
INVX1 gate4305(.O (I16124), .I (g10396));
INVX1 gate4306(.O (g10909), .I (I16679));
INVX1 gate4307(.O (I12535), .I (g7656));
INVX1 gate4308(.O (g5778), .I (I9368));
INVX1 gate4309(.O (I10174), .I (g5994));
INVX1 gate4310(.O (I15669), .I (g10194));
INVX1 gate4311(.O (g10543), .I (I16196));
INVX1 gate4312(.O (g3784), .I (g2586));
INVX1 gate4313(.O (I17413), .I (g11425));
INVX1 gate4314(.O (g5894), .I (g5361));
INVX1 gate4315(.O (g9826), .I (I14979));
INVX1 gate4316(.O (g10117), .I (I15359));
INVX1 gate4317(.O (g8660), .I (I13945));
INVX1 gate4318(.O (g8946), .I (I14295));
INVX1 gate4319(.O (g10908), .I (I16676));
INVX1 gate4320(.O (g2916), .I (I6097));
INVX1 gate4321(.O (I7843), .I (g3440));
INVX1 gate4322(.O (g2022), .I (g1346));
INVX1 gate4323(.O (g5735), .I (I9293));
INVX1 gate4324(.O (I15392), .I (g10104));
INVX1 gate4325(.O (g7677), .I (g7148));
INVX1 gate4326(.O (g2749), .I (I5815));
INVX1 gate4327(.O (g3995), .I (g3121));
INVX1 gate4328(.O (g3937), .I (I7086));
INVX1 gate4329(.O (I10840), .I (g6719));
INVX1 gate4330(.O (g9741), .I (I14888));
INVX1 gate4331(.O (g4002), .I (g3121));
INVX1 gate4332(.O (I7393), .I (g4096));
INVX1 gate4333(.O (I16938), .I (g11086));
INVX1 gate4334(.O (I6531), .I (g3186));
INVX1 gate4335(.O (I11348), .I (g6695));
INVX1 gate4336(.O (I12344), .I (g7062));
INVX1 gate4337(.O (I13083), .I (g7921));
INVX1 gate4338(.O (g3479), .I (g2655));
INVX1 gate4339(.O (g11195), .I (g11112));
INVX1 gate4340(.O (g11489), .I (I17482));
INVX1 gate4341(.O (g6131), .I (g5548));
INVX1 gate4342(.O (g5661), .I (I9144));
INVX1 gate4343(.O (g10747), .I (I16432));
INVX1 gate4344(.O (I15559), .I (g10094));
INVX1 gate4345(.O (g5075), .I (g4439));
INVX1 gate4346(.O (g8513), .I (I13708));
INVX1 gate4347(.O (I15488), .I (g10116));
INVX1 gate4348(.O (I15424), .I (g10080));
INVX1 gate4349(.O (g6406), .I (I10314));
INVX1 gate4350(.O (g10242), .I (I15632));
INVX1 gate4351(.O (I8007), .I (g3829));
INVX1 gate4352(.O (g5475), .I (I8892));
INVX1 gate4353(.O (g4762), .I (I8116));
INVX1 gate4354(.O (g2798), .I (g2449));
INVX1 gate4355(.O (g5949), .I (I9591));
INVX1 gate4356(.O (g7349), .I (I11695));
INVX1 gate4357(.O (I10192), .I (g6115));
INVX1 gate4358(.O (g11424), .I (I17327));
INVX1 gate4359(.O (I9240), .I (g5069));
INVX1 gate4360(.O (g6635), .I (I10592));
INVX1 gate4361(.O (I11566), .I (g6820));
INVX1 gate4362(.O (g11016), .I (I16739));
INVX1 gate4363(.O (g9108), .I (I14449));
INVX1 gate4364(.O (g3390), .I (g3161));
INVX1 gate4365(.O (g9308), .I (I14499));
INVX1 gate4366(.O (g8036), .I (I12878));
INVX1 gate4367(.O (g2560), .I (I5684));
INVX1 gate4368(.O (g5627), .I (g4840));
INVX1 gate4369(.O (g8436), .I (I13606));
INVX1 gate4370(.O (g8178), .I (I13083));
INVX1 gate4371(.O (g6801), .I (I10813));
INVX1 gate4372(.O (g6305), .I (I10174));
INVX1 gate4373(.O (I6856), .I (g3318));
INVX1 gate4374(.O (g4590), .I (I7999));
INVX1 gate4375(.O (g7848), .I (I12641));
INVX1 gate4376(.O (g5292), .I (g4445));
INVX1 gate4377(.O (I10663), .I (g6040));
INVX1 gate4378(.O (g8378), .I (I13482));
INVX1 gate4379(.O (g9883), .I (I15060));
INVX1 gate4380(.O (I9043), .I (g4786));
INVX1 gate4381(.O (g3501), .I (g3077));
INVX1 gate4382(.O (I14522), .I (g9108));
INVX1 gate4383(.O (I8535), .I (g4340));
INVX1 gate4384(.O (I9443), .I (g5557));
INVX1 gate4385(.O (g7747), .I (I12406));
INVX1 gate4386(.O (g5998), .I (I9620));
INVX1 gate4387(.O (g5646), .I (I9099));
INVX1 gate4388(.O (g10974), .I (I16723));
INVX1 gate4389(.O (g8335), .I (I13385));
INVX1 gate4390(.O (g2873), .I (I6019));
INVX1 gate4391(.O (g6748), .I (I10753));
INVX1 gate4392(.O (g2632), .I (g2002));
INVX1 gate4393(.O (I6074), .I (g2228));
INVX1 gate4394(.O (g2095), .I (g143));
INVX1 gate4395(.O (I11653), .I (g6954));
INVX1 gate4396(.O (g2037), .I (g1771));
INVX1 gate4397(.O (g8182), .I (I13099));
INVX1 gate4398(.O (I4886), .I (g257));
INVX1 gate4399(.O (g4222), .I (g3638));
INVX1 gate4400(.O (g5603), .I (I9029));
INVX1 gate4401(.O (I6474), .I (g2297));
INVX1 gate4402(.O (I7625), .I (g4164));
INVX1 gate4403(.O (g5039), .I (I8418));
INVX1 gate4404(.O (I4951), .I (g262));
INVX1 gate4405(.O (g10293), .I (I15701));
INVX1 gate4406(.O (g2653), .I (g2011));
INVX1 gate4407(.O (g2208), .I (g84));
INVX1 gate4408(.O (g2302), .I (g29));
INVX1 gate4409(.O (I12029), .I (g6922));
INVX1 gate4410(.O (g5850), .I (g5320));
INVX1 gate4411(.O (g6226), .I (I9973));
INVX1 gate4412(.O (I10553), .I (g6192));
INVX1 gate4413(.O (g3704), .I (I6861));
INVX1 gate4414(.O (g8805), .I (I14136));
INVX1 gate4415(.O (g10265), .I (g10143));
INVX1 gate4416(.O (g2579), .I (g1969));
INVX1 gate4417(.O (I5837), .I (g2507));
INVX1 gate4418(.O (I7938), .I (g3406));
INVX1 gate4419(.O (I9147), .I (g5011));
INVX1 gate4420(.O (I13636), .I (g8357));
INVX1 gate4421(.O (g8422), .I (I13580));
INVX1 gate4422(.O (I10949), .I (g6747));
INVX1 gate4423(.O (I17302), .I (g11391));
INVX1 gate4424(.O (g4899), .I (I8262));
INVX1 gate4425(.O (I11333), .I (g6670));
INVX1 gate4426(.O (I13415), .I (g8144));
INVX1 gate4427(.O (g4464), .I (I7829));
INVX1 gate4428(.O (g2719), .I (g2043));
INVX1 gate4429(.O (g9448), .I (g9091));
INVX1 gate4430(.O (I7909), .I (g3387));
INVX1 gate4431(.O (I6080), .I (g2108));
INVX1 gate4432(.O (I14326), .I (g8818));
INVX1 gate4433(.O (g4785), .I (g3337));
INVX1 gate4434(.O (g11042), .I (I16787));
INVX1 gate4435(.O (g10391), .I (g10313));
INVX1 gate4436(.O (I6480), .I (g2462));
INVX1 gate4437(.O (g5702), .I (I9243));
INVX1 gate4438(.O (g6445), .I (I10367));
INVX1 gate4439(.O (g2752), .I (I5824));
INVX1 gate4440(.O (I14040), .I (g8649));
INVX1 gate4441(.O (I14948), .I (g9555));
INVX1 gate4442(.O (g9827), .I (I14982));
INVX1 gate4443(.O (g6091), .I (I9744));
INVX1 gate4444(.O (I10702), .I (g6071));
INVX1 gate4445(.O (g3810), .I (g3228));
INVX1 gate4446(.O (g3363), .I (I6549));
INVX1 gate4447(.O (I10904), .I (g6558));
INVX1 gate4448(.O (g8798), .I (I14119));
INVX1 gate4449(.O (g7119), .I (I11354));
INVX1 gate4450(.O (g7319), .I (I11605));
INVX1 gate4451(.O (g3432), .I (g3144));
INVX1 gate4452(.O (I6569), .I (g3186));
INVX1 gate4453(.O (g10579), .I (g10528));
INVX1 gate4454(.O (g4563), .I (g3946));
INVX1 gate4455(.O (g9774), .I (g9474));
INVX1 gate4456(.O (I7606), .I (g4166));
INVX1 gate4457(.O (g8560), .I (I13773));
INVX1 gate4458(.O (I14252), .I (g8783));
INVX1 gate4459(.O (g6169), .I (I9896));
INVX1 gate4460(.O (I15383), .I (g10107));
INVX1 gate4461(.O (I16277), .I (g10536));
INVX1 gate4462(.O (g6283), .I (I10108));
INVX1 gate4463(.O (g7352), .I (I11704));
INVX1 gate4464(.O (g2042), .I (g1796));
INVX1 gate4465(.O (g4295), .I (I7556));
INVX1 gate4466(.O (g10578), .I (g10527));
INVX1 gate4467(.O (I9013), .I (g4767));
INVX1 gate4468(.O (g4237), .I (g4013));
INVX1 gate4469(.O (g6407), .I (I10317));
INVX1 gate4470(.O (I14564), .I (g9026));
INVX1 gate4471(.O (g6920), .I (I11034));
INVX1 gate4472(.O (g6578), .I (I10526));
INVX1 gate4473(.O (g6868), .I (I10946));
INVX1 gate4474(.O (g5616), .I (I9046));
INVX1 gate4475(.O (I16595), .I (g10783));
INVX1 gate4476(.O (g8873), .I (I14191));
INVX1 gate4477(.O (g8632), .I (I13915));
INVX1 gate4478(.O (g8095), .I (g7942));
INVX1 gate4479(.O (g2164), .I (I5095));
INVX1 gate4480(.O (g6718), .I (g5949));
INVX1 gate4481(.O (g2364), .I (g611));
INVX1 gate4482(.O (g2233), .I (I5224));
INVX1 gate4483(.O (g9780), .I (g9474));
INVX1 gate4484(.O (g4194), .I (I7399));
INVX1 gate4485(.O (I16623), .I (g10858));
INVX1 gate4486(.O (g8437), .I (I13609));
INVX1 gate4487(.O (I10183), .I (g6108));
INVX1 gate4488(.O (I7586), .I (g4127));
INVX1 gate4489(.O (g11065), .I (g10974));
INVX1 gate4490(.O (g4394), .I (I7729));
INVX1 gate4491(.O (I5192), .I (g55));
INVX1 gate4492(.O (I6976), .I (g2884));
INVX1 gate4493(.O (g2054), .I (g1864));
INVX1 gate4494(.O (g6582), .I (g5949));
INVX1 gate4495(.O (I13609), .I (g8312));
INVX1 gate4496(.O (I14397), .I (g8888));
INVX1 gate4497(.O (g7386), .I (I11767));
INVX1 gate4498(.O (g4731), .I (I8085));
INVX1 gate4499(.O (I11312), .I (g6488));
INVX1 gate4500(.O (g5647), .I (I9102));
INVX1 gate4501(.O (g2454), .I (I5549));
INVX1 gate4502(.O (g8579), .I (I13822));
INVX1 gate4503(.O (g8869), .I (I14179));
INVX1 gate4504(.O (g7975), .I (I12773));
INVX1 gate4505(.O (I13200), .I (g8251));
INVX1 gate4506(.O (g6261), .I (I10042));
INVX1 gate4507(.O (I11608), .I (g6903));
INVX1 gate4508(.O (g2296), .I (I5332));
INVX1 gate4509(.O (I11115), .I (g6462));
INVX1 gate4510(.O (I12604), .I (g7630));
INVX1 gate4511(.O (g10116), .I (I15356));
INVX1 gate4512(.O (I9117), .I (g5615));
INVX1 gate4513(.O (g6793), .I (I10795));
INVX1 gate4514(.O (g8719), .I (g8579));
INVX1 gate4515(.O (g4557), .I (g3946));
INVX1 gate4516(.O (I9317), .I (g5576));
INVX1 gate4517(.O (g2725), .I (g2018));
INVX1 gate4518(.O (g1974), .I (g627));
INVX1 gate4519(.O (I14509), .I (g8926));
INVX1 gate4520(.O (g5546), .I (I8973));
INVX1 gate4521(.O (g7026), .I (I11173));
INVX1 gate4522(.O (I5854), .I (g2523));
INVX1 gate4523(.O (I8388), .I (g4239));
INVX1 gate4524(.O (g4966), .I (I8340));
INVX1 gate4525(.O (I12770), .I (g7638));
INVX1 gate4526(.O (I14933), .I (g9454));
INVX1 gate4527(.O (g7426), .I (I11814));
INVX1 gate4528(.O (g9994), .I (I15196));
INVX1 gate4529(.O (g9290), .I (I14494));
INVX1 gate4530(.O (I11921), .I (g6904));
INVX1 gate4531(.O (I17662), .I (g11602));
INVX1 gate4532(.O (I12981), .I (g8041));
INVX1 gate4533(.O (g8752), .I (g8635));
INVX1 gate4534(.O (g6227), .I (g5446));
INVX1 gate4535(.O (g10041), .I (I15250));
INVX1 gate4536(.O (g5503), .I (g4515));
INVX1 gate4537(.O (I7710), .I (g3749));
INVX1 gate4538(.O (g7614), .I (I12190));
INVX1 gate4539(.O (g10275), .I (I15669));
INVX1 gate4540(.O (g4242), .I (g3664));
INVX1 gate4541(.O (g10493), .I (I16114));
INVX1 gate4542(.O (g7325), .I (I11623));
INVX1 gate4543(.O (I17249), .I (g11342));
INVX1 gate4544(.O (g4948), .I (I8315));
INVX1 gate4545(.O (I7691), .I (g3363));
INVX1 gate4546(.O (g9816), .I (g9490));
INVX1 gate4547(.O (I17482), .I (g11479));
INVX1 gate4548(.O (g10465), .I (I15986));
INVX1 gate4549(.O (g1980), .I (g646));
INVX1 gate4550(.O (I8247), .I (g4615));
INVX1 gate4551(.O (g7984), .I (I12796));
INVX1 gate4552(.O (g2012), .I (g981));
INVX1 gate4553(.O (g11160), .I (g10950));
INVX1 gate4554(.O (g8442), .I (I13624));
INVX1 gate4555(.O (I17710), .I (g11620));
INVX1 gate4556(.O (g6203), .I (g5446));
INVX1 gate4557(.O (I17552), .I (g11502));
INVX1 gate4558(.O (I16853), .I (g10907));
INVX1 gate4559(.O (I9581), .I (g5111));
INVX1 gate4560(.O (g10035), .I (I15241));
INVX1 gate4561(.O (g5120), .I (I8520));
INVX1 gate4562(.O (I5031), .I (g928));
INVX1 gate4563(.O (g5320), .I (g4418));
INVX1 gate4564(.O (g4254), .I (g4013));
INVX1 gate4565(.O (I16589), .I (g10820));
INVX1 gate4566(.O (I11674), .I (g7051));
INVX1 gate4567(.O (g10806), .I (I16518));
INVX1 gate4568(.O (g7544), .I (I11964));
INVX1 gate4569(.O (g8164), .I (g7872));
INVX1 gate4570(.O (I13674), .I (g8304));
INVX1 gate4571(.O (I15470), .I (g10111));
INVX1 gate4572(.O (I5812), .I (g2090));
INVX1 gate4573(.O (g8233), .I (g7872));
INVX1 gate4574(.O (g11617), .I (I17669));
INVX1 gate4575(.O (I6183), .I (g2131));
INVX1 gate4576(.O (g11470), .I (I17447));
INVX1 gate4577(.O (I7659), .I (g3731));
INVX1 gate4578(.O (g10142), .I (I15424));
INVX1 gate4579(.O (g2888), .I (I6046));
INVX1 gate4580(.O (I6924), .I (g2843));
INVX1 gate4581(.O (g7636), .I (I12248));
INVX1 gate4582(.O (I6220), .I (g883));
INVX1 gate4583(.O (I4891), .I (g582));
INVX1 gate4584(.O (g2171), .I (I5116));
INVX1 gate4585(.O (g4438), .I (I7790));
INVX1 gate4586(.O (I14452), .I (g8922));
INVX1 gate4587(.O (g4773), .I (I8133));
INVX1 gate4588(.O (g7306), .I (I11566));
INVX1 gate4589(.O (I13732), .I (g8291));
INVX1 gate4590(.O (g8296), .I (I13242));
INVX1 gate4591(.O (g2956), .I (I6159));
INVX1 gate4592(.O (I15075), .I (g9761));
INVX1 gate4593(.O (g8725), .I (g8589));
INVX1 gate4594(.O (g7790), .I (I12535));
INVX1 gate4595(.O (g9263), .I (g8892));
INVX1 gate4596(.O (g3683), .I (I6844));
INVX1 gate4597(.O (g11075), .I (g10937));
INVX1 gate4598(.O (I5765), .I (g2004));
INVX1 gate4599(.O (I15595), .I (g10165));
INVX1 gate4600(.O (I15467), .I (g10079));
INVX1 gate4601(.O (I15494), .I (g10117));
INVX1 gate4602(.O (I17356), .I (g11384));
INVX1 gate4603(.O (g8532), .I (I13741));
INVX1 gate4604(.O (I8308), .I (g4443));
INVX1 gate4605(.O (g7187), .I (I11405));
INVX1 gate4606(.O (I7311), .I (g2803));
INVX1 gate4607(.O (g4769), .I (g3586));
INVX1 gate4608(.O (g5987), .I (I9605));
INVX1 gate4609(.O (I11692), .I (g7048));
INVX1 gate4610(.O (g7387), .I (I11770));
INVX1 gate4611(.O (g11467), .I (I17438));
INVX1 gate4612(.O (I9995), .I (g5536));
INVX1 gate4613(.O (I12832), .I (g7681));
INVX1 gate4614(.O (I4859), .I (g578));
INVX1 gate4615(.O (I10051), .I (g5702));
INVX1 gate4616(.O (I10072), .I (g5719));
INVX1 gate4617(.O (g4212), .I (I7453));
INVX1 gate4618(.O (I9479), .I (g4954));
INVX1 gate4619(.O (g6689), .I (g5830));
INVX1 gate4620(.O (g10130), .I (I15392));
INVX1 gate4621(.O (g7756), .I (I12433));
INVX1 gate4622(.O (g2297), .I (g865));
INVX1 gate4623(.O (g11623), .I (I17687));
INVX1 gate4624(.O (g6388), .I (I10286));
INVX1 gate4625(.O (g10193), .I (g10057));
INVX1 gate4626(.O (I16616), .I (g10796));
INVX1 gate4627(.O (g11037), .I (I16772));
INVX1 gate4628(.O (I10592), .I (g5865));
INVX1 gate4629(.O (g5299), .I (g4393));
INVX1 gate4630(.O (I10756), .I (g5810));
INVX1 gate4631(.O (I15782), .I (g10259));
INVX1 gate4632(.O (g7622), .I (g7067));
INVX1 gate4633(.O (g3735), .I (I6921));
INVX1 gate4634(.O (g7027), .I (I11176));
INVX1 gate4635(.O (g7427), .I (I11817));
INVX1 gate4636(.O (I17182), .I (g11309));
INVX1 gate4637(.O (g10165), .I (I15491));
INVX1 gate4638(.O (I13400), .I (g8236));
INVX1 gate4639(.O (g10523), .I (g10456));
INVX1 gate4640(.O (I17672), .I (g11605));
INVX1 gate4641(.O (g3782), .I (I7006));
INVX1 gate4642(.O (I13013), .I (g8048));
INVX1 gate4643(.O (g5892), .I (I9519));
INVX1 gate4644(.O (I11214), .I (g6528));
INVX1 gate4645(.O (g7904), .I (I12690));
INVX1 gate4646(.O (g11419), .I (I17312));
INVX1 gate4647(.O (g2745), .I (I5809));
INVX1 gate4648(.O (g2639), .I (I5754));
INVX1 gate4649(.O (g6030), .I (I9639));
INVX1 gate4650(.O (g2338), .I (g1909));
INVX1 gate4651(.O (g11352), .I (I17173));
INVX1 gate4652(.O (I15418), .I (g10083));
INVX1 gate4653(.O (I5073), .I (g34));
INVX1 gate4654(.O (I13329), .I (g8116));
INVX1 gate4655(.O (I11207), .I (g6524));
INVX1 gate4656(.O (g7446), .I (g7148));
INVX1 gate4657(.O (g3475), .I (g3056));
INVX1 gate4658(.O (I6999), .I (g2905));
INVX1 gate4659(.O (g11155), .I (g10950));
INVX1 gate4660(.O (I7284), .I (g3255));
INVX1 gate4661(.O (I15266), .I (g10001));
INVX1 gate4662(.O (g8990), .I (I14391));
INVX1 gate4663(.O (I9156), .I (g5032));
INVX1 gate4664(.O (I12099), .I (g7258));
INVX1 gate4665(.O (I11005), .I (g6386));
INVX1 gate4666(.O (I12388), .I (g7219));
INVX1 gate4667(.O (I17331), .I (g11357));
INVX1 gate4668(.O (I13005), .I (g8046));
INVX1 gate4669(.O (g8888), .I (I14232));
INVX1 gate4670(.O (g7403), .I (I11783));
INVX1 gate4671(.O (g3627), .I (I6784));
INVX1 gate4672(.O (g4822), .I (g3706));
INVX1 gate4673(.O (g8029), .I (I12871));
INVX1 gate4674(.O (g6564), .I (g5784));
INVX1 gate4675(.O (I16808), .I (g10906));
INVX1 gate4676(.O (g8171), .I (I13068));
INVX1 gate4677(.O (g7345), .I (I11683));
INVX1 gate4678(.O (I17513), .I (g11482));
INVX1 gate4679(.O (I8711), .I (g4530));
INVX1 gate4680(.O (g2808), .I (g2156));
INVX1 gate4681(.O (g3292), .I (g2373));
INVX1 gate4682(.O (I10846), .I (g6729));
INVX1 gate4683(.O (g8787), .I (I14094));
INVX1 gate4684(.O (I12251), .I (g7076));
INVX1 gate4685(.O (g7763), .I (I12454));
INVX1 gate4686(.O (I16101), .I (g10381));
INVX1 gate4687(.O (g8956), .I (I14319));
INVX1 gate4688(.O (g2707), .I (g2041));
INVX1 gate4689(.O (I8827), .I (g4477));
INVX1 gate4690(.O (g10437), .I (g10333));
INVX1 gate4691(.O (I8133), .I (g3632));
INVX1 gate4692(.O (g2759), .I (I5843));
INVX1 gate4693(.O (I8333), .I (g4456));
INVX1 gate4694(.O (I7420), .I (g4167));
INVX1 gate4695(.O (g7637), .I (I12251));
INVX1 gate4696(.O (I15589), .I (g10161));
INVX1 gate4697(.O (g5078), .I (g4372));
INVX1 gate4698(.O (g3039), .I (g2310));
INVX1 gate4699(.O (g2201), .I (g102));
INVX1 gate4700(.O (g3439), .I (g3144));
INVX1 gate4701(.O (g7107), .I (I11342));
INVX1 gate4702(.O (I7559), .I (g4116));
INVX1 gate4703(.O (g7307), .I (I11569));
INVX1 gate4704(.O (I12032), .I (g6923));
INVX1 gate4705(.O (g8297), .I (I13245));
INVX1 gate4706(.O (g10347), .I (I15807));
INVX1 gate4707(.O (g5035), .I (I8410));
INVX1 gate4708(.O (I6944), .I (g2859));
INVX1 gate4709(.O (I8396), .I (g4255));
INVX1 gate4710(.O (g10253), .I (g10138));
INVX1 gate4711(.O (I6240), .I (g878));
INVX1 gate4712(.O (I7931), .I (g3624));
INVX1 gate4713(.O (g7359), .I (I11725));
INVX1 gate4714(.O (g6108), .I (I9779));
INVX1 gate4715(.O (g6308), .I (I10183));
INVX1 gate4716(.O (I9810), .I (g5576));
INVX1 gate4717(.O (g5082), .I (g4840));
INVX1 gate4718(.O (g2449), .I (g790));
INVX1 gate4719(.O (I9032), .I (g4732));
INVX1 gate4720(.O (I11100), .I (g6442));
INVX1 gate4721(.O (g5482), .I (I8903));
INVX1 gate4722(.O (I14405), .I (g8937));
INVX1 gate4723(.O (g10600), .I (I16277));
INVX1 gate4724(.O (g11401), .I (I17246));
INVX1 gate4725(.O (g10781), .I (I16475));
INVX1 gate4726(.O (I4783), .I (g873));
INVX1 gate4727(.O (I6043), .I (g2267));
INVX1 gate4728(.O (I9053), .I (g4752));
INVX1 gate4729(.O (g8684), .I (I13969));
INVX1 gate4730(.O (g3583), .I (I6742));
INVX1 gate4731(.O (g4895), .I (I8250));
INVX1 gate4732(.O (g5876), .I (g5361));
INVX1 gate4733(.O (g8138), .I (I13013));
INVX1 gate4734(.O (I6443), .I (g2363));
INVX1 gate4735(.O (I11235), .I (g6538));
INVX1 gate4736(.O (g8338), .I (I13394));
INVX1 gate4737(.O (g10236), .I (g10190));
INVX1 gate4738(.O (g7757), .I (I12436));
INVX1 gate4739(.O (g2604), .I (I5713));
INVX1 gate4740(.O (g4062), .I (I7185));
INVX1 gate4741(.O (g2098), .I (I4938));
INVX1 gate4742(.O (I11683), .I (g7069));
INVX1 gate4743(.O (g5656), .I (I9129));
INVX1 gate4744(.O (g7416), .I (I11800));
INVX1 gate4745(.O (g4620), .I (I8031));
INVX1 gate4746(.O (g10351), .I (I15817));
INVX1 gate4747(.O (g4462), .I (I7825));
INVX1 gate4748(.O (I15864), .I (g10339));
INVX1 gate4749(.O (I5399), .I (g895));
INVX1 gate4750(.O (g6589), .I (I10549));
INVX1 gate4751(.O (I12871), .I (g7638));
INVX1 gate4752(.O (g10175), .I (I15517));
INVX1 gate4753(.O (g10821), .I (I16531));
INVX1 gate4754(.O (I7630), .I (g3524));
INVX1 gate4755(.O (I15749), .I (g10263));
INVX1 gate4756(.O (g2833), .I (I5949));
INVX1 gate4757(.O (I6034), .I (g2210));
INVX1 gate4758(.O (g7522), .I (I11904));
INVX1 gate4759(.O (I8418), .I (g4794));
INVX1 gate4760(.O (g7811), .I (I12598));
INVX1 gate4761(.O (g7315), .I (I11593));
INVX1 gate4762(.O (g11616), .I (I17666));
INVX1 gate4763(.O (I17149), .I (g11306));
INVX1 gate4764(.O (I6565), .I (g2614));
INVX1 gate4765(.O (g7047), .I (I11222));
INVX1 gate4766(.O (I7300), .I (g2883));
INVX1 gate4767(.O (g11313), .I (I17104));
INVX1 gate4768(.O (I12360), .I (g7183));
INVX1 gate4769(.O (I8290), .I (g4778));
INVX1 gate4770(.O (g10063), .I (I15287));
INVX1 gate4771(.O (I17387), .I (g11438));
INVX1 gate4772(.O (g8707), .I (g8671));
INVX1 gate4773(.O (g6165), .I (g5446));
INVX1 gate4774(.O (g10264), .I (g10128));
INVX1 gate4775(.O (g6571), .I (I10503));
INVX1 gate4776(.O (g6365), .I (I10274));
INVX1 gate4777(.O (g6861), .I (I10941));
INVX1 gate4778(.O (g5214), .I (g4640));
INVX1 gate4779(.O (g10137), .I (I15409));
INVX1 gate4780(.O (g6048), .I (I9673));
INVX1 gate4781(.O (I11515), .I (g6589));
INVX1 gate4782(.O (g9772), .I (g9432));
INVX1 gate4783(.O (I11882), .I (g6895));
INVX1 gate4784(.O (I5510), .I (g588));
INVX1 gate4785(.O (g2539), .I (I5652));
INVX1 gate4786(.O (g2896), .I (g2356));
INVX1 gate4787(.O (I6347), .I (g2462));
INVX1 gate4788(.O (I15704), .I (g10238));
INVX1 gate4789(.O (I5245), .I (g925));
INVX1 gate4790(.O (g6448), .I (I10374));
INVX1 gate4791(.O (g9531), .I (I14678));
INVX1 gate4792(.O (I15305), .I (g10001));
INVX1 gate4793(.O (g6711), .I (g5949));
INVX1 gate4794(.O (g6055), .I (I9688));
INVX1 gate4795(.O (I12162), .I (g7146));
INVX1 gate4796(.O (I17104), .I (g11223));
INVX1 gate4797(.O (g10873), .I (I16589));
INVX1 gate4798(.O (g11053), .I (g10950));
INVX1 gate4799(.O (I8256), .I (g4711));
INVX1 gate4800(.O (g9890), .I (I15075));
INVX1 gate4801(.O (I10282), .I (g6163));
INVX1 gate4802(.O (g3404), .I (g3121));
INVX1 gate4803(.O (g6133), .I (I9836));
INVX1 gate4804(.O (g11466), .I (I17435));
INVX1 gate4805(.O (g5663), .I (I9150));
INVX1 gate4806(.O (I10302), .I (g6179));
INVX1 gate4807(.O (I6914), .I (g2828));
INVX1 gate4808(.O (g9505), .I (g9052));
INVX1 gate4809(.O (g2162), .I (I5089));
INVX1 gate4810(.O (I7973), .I (g3437));
INVX1 gate4811(.O (I15036), .I (g9721));
INVX1 gate4812(.O (g2268), .I (g654));
INVX1 gate4813(.O (g8449), .I (I13645));
INVX1 gate4814(.O (g4192), .I (I7393));
INVX1 gate4815(.O (I10105), .I (g5736));
INVX1 gate4816(.O (g4298), .I (g4130));
INVX1 gate4817(.O (g3764), .I (I6971));
INVX1 gate4818(.O (I12451), .I (g7538));
INVX1 gate4819(.O (g6846), .I (I10910));
INVX1 gate4820(.O (g11036), .I (I16769));
INVX1 gate4821(.O (I12472), .I (g7539));
INVX1 gate4822(.O (g8575), .I (I13816));
INVX1 gate4823(.O (g3546), .I (g3307));
INVX1 gate4824(.O (I14105), .I (g8776));
INVX1 gate4825(.O (g4485), .I (g3546));
INVX1 gate4826(.O (I6013), .I (g2200));
INVX1 gate4827(.O (g5402), .I (I8842));
INVX1 gate4828(.O (g6196), .I (g5446));
INVX1 gate4829(.O (g7880), .I (g7479));
INVX1 gate4830(.O (g6396), .I (I10296));
INVX1 gate4831(.O (g7595), .I (I12123));
INVX1 gate4832(.O (g6803), .I (I10819));
INVX1 gate4833(.O (g7537), .I (I11947));
INVX1 gate4834(.O (g5236), .I (g4361));
INVX1 gate4835(.O (I17368), .I (g11423));
INVX1 gate4836(.O (g8604), .I (g8479));
INVX1 gate4837(.O (g10208), .I (I15580));
INVX1 gate4838(.O (I16239), .I (g10525));
INVX1 gate4839(.O (g11642), .I (I17730));
INVX1 gate4840(.O (g8498), .I (g8353));
INVX1 gate4841(.O (I11584), .I (g6827));
INVX1 gate4842(.O (g1972), .I (g461));
INVX1 gate4843(.O (I8421), .I (g4309));
INVX1 gate4844(.O (g9474), .I (g9331));
INVX1 gate4845(.O (g7272), .I (I11519));
INVX1 gate4846(.O (I13206), .I (g8197));
INVX1 gate4847(.O (g10542), .I (I16193));
INVX1 gate4848(.O (g6509), .I (I10427));
INVX1 gate4849(.O (g11064), .I (g10974));
INVX1 gate4850(.O (I15733), .I (g10257));
INVX1 gate4851(.O (g7612), .I (I12186));
INVX1 gate4852(.O (g7243), .I (I11483));
INVX1 gate4853(.O (g2086), .I (I4906));
INVX1 gate4854(.O (I11759), .I (g7244));
INVX1 gate4855(.O (I11725), .I (g7040));
INVX1 gate4856(.O (I12776), .I (g7586));
INVX1 gate4857(.O (g5657), .I (I9132));
INVX1 gate4858(.O (g10913), .I (I16691));
INVX1 gate4859(.O (I16941), .I (g11076));
INVX1 gate4860(.O (g2728), .I (g2025));
INVX1 gate4861(.O (I13114), .I (g7930));
INVX1 gate4862(.O (g6418), .I (g6137));
INVX1 gate4863(.O (I11082), .I (g6749));
INVX1 gate4864(.O (g7982), .I (I12790));
INVX1 gate4865(.O (g4520), .I (I7923));
INVX1 gate4866(.O (g5222), .I (g4640));
INVX1 gate4867(.O (I17228), .I (g11300));
INVX1 gate4868(.O (g11630), .I (I17704));
INVX1 gate4869(.O (g2185), .I (g46));
INVX1 gate4870(.O (g4219), .I (g3635));
INVX1 gate4871(.O (g6290), .I (I10129));
INVX1 gate4872(.O (I7151), .I (g2642));
INVX1 gate4873(.O (g2881), .I (I6031));
INVX1 gate4874(.O (I7351), .I (g4061));
INVX1 gate4875(.O (I16518), .I (g10718));
INVX1 gate4876(.O (I6601), .I (g3186));
INVX1 gate4877(.O (I7648), .I (g3727));
INVX1 gate4878(.O (I12825), .I (g7696));
INVX1 gate4879(.O (g10320), .I (I15756));
INVX1 gate4880(.O (g10905), .I (I16667));
INVX1 gate4881(.O (g7629), .I (I12229));
INVX1 gate4882(.O (I15665), .I (g10193));
INVX1 gate4883(.O (g7328), .I (I11632));
INVX1 gate4884(.O (g2070), .I (g213));
INVX1 gate4885(.O (g10530), .I (g10466));
INVX1 gate4886(.O (g3906), .I (g3015));
INVX1 gate4887(.O (I17716), .I (g11622));
INVX1 gate4888(.O (g7330), .I (I11638));
INVX1 gate4889(.O (g10593), .I (I16264));
INVX1 gate4890(.O (I4866), .I (g579));
INVX1 gate4891(.O (g8362), .I (I13466));
INVX1 gate4892(.O (I13744), .I (g8297));
INVX1 gate4893(.O (g2025), .I (g1696));
INVX1 gate4894(.O (I11345), .I (g6692));
INVX1 gate4895(.O (g10346), .I (I15804));
INVX1 gate4896(.O (I8631), .I (g4425));
INVX1 gate4897(.O (g5899), .I (g5361));
INVX1 gate4898(.O (g8419), .I (I13571));
INVX1 gate4899(.O (g4958), .I (I8328));
INVX1 gate4900(.O (g6256), .I (I10027));
INVX1 gate4901(.O (g4176), .I (I7345));
INVX1 gate4902(.O (g6816), .I (I10858));
INVX1 gate4903(.O (g10122), .I (I15374));
INVX1 gate4904(.O (g4376), .I (I7691));
INVX1 gate4905(.O (g4005), .I (I7143));
INVX1 gate4906(.O (g10464), .I (I15983));
INVX1 gate4907(.O (I10027), .I (g5751));
INVX1 gate4908(.O (I15476), .I (g10114));
INVX1 gate4909(.O (I15485), .I (g10092));
INVX1 gate4910(.O (g7800), .I (I12565));
INVX1 gate4911(.O (g10034), .I (I15238));
INVX1 gate4912(.O (g6181), .I (g5426));
INVX1 gate4913(.O (I11804), .I (g7190));
INVX1 gate4914(.O (I14249), .I (g8804));
INVX1 gate4915(.O (g11454), .I (I17419));
INVX1 gate4916(.O (g6847), .I (g6482));
INVX1 gate4917(.O (g10292), .I (I15698));
INVX1 gate4918(.O (I9475), .I (g5445));
INVX1 gate4919(.O (I10248), .I (g6125));
INVX1 gate4920(.O (g6685), .I (I10648));
INVX1 gate4921(.O (g6197), .I (I9930));
INVX1 gate4922(.O (g6700), .I (g5949));
INVX1 gate4923(.O (I17112), .I (g11227));
INVX1 gate4924(.O (I10710), .I (g6088));
INVX1 gate4925(.O (g6397), .I (I10299));
INVX1 gate4926(.O (I10003), .I (g4908));
INVX1 gate4927(.O (g7213), .I (I11447));
INVX1 gate4928(.O (I10204), .I (g6031));
INVX1 gate4929(.O (I14552), .I (g9264));
INVX1 gate4930(.O (I5336), .I (g1700));
INVX1 gate4931(.O (g2131), .I (I5060));
INVX1 gate4932(.O (g8486), .I (g8348));
INVX1 gate4933(.O (I6784), .I (g2742));
INVX1 gate4934(.O (g2006), .I (g932));
INVX1 gate4935(.O (g2331), .I (g658));
INVX1 gate4936(.O (I16577), .I (g10825));
INVX1 gate4937(.O (g4733), .I (I8089));
INVX1 gate4938(.O (g2406), .I (g1365));
INVX1 gate4939(.O (g5844), .I (I9461));
INVX1 gate4940(.O (I13332), .I (g8206));
INVX1 gate4941(.O (g6263), .I (I10048));
INVX1 gate4942(.O (g4270), .I (g4013));
INVX1 gate4943(.O (I11135), .I (g6679));
INVX1 gate4944(.O (I7372), .I (g4057));
INVX1 gate4945(.O (g10136), .I (I15406));
INVX1 gate4946(.O (g2635), .I (g2003));
INVX1 gate4947(.O (I16439), .I (g10702));
INVX1 gate4948(.O (I17742), .I (g11636));
INVX1 gate4949(.O (I12318), .I (g6862));
INVX1 gate4950(.O (g11074), .I (g10901));
INVX1 gate4951(.O (g6950), .I (I11094));
INVX1 gate4952(.O (g11239), .I (g11112));
INVX1 gate4953(.O (I10081), .I (g5735));
INVX1 gate4954(.O (I17096), .I (g11219));
INVX1 gate4955(.O (g4225), .I (I7478));
INVX1 gate4956(.O (I15238), .I (g9974));
INVX1 gate4957(.O (g2087), .I (g225));
INVX1 gate4958(.O (g11594), .I (I17636));
INVX1 gate4959(.O (g3945), .I (I7096));
INVX1 gate4960(.O (I7143), .I (g2614));
INVX1 gate4961(.O (I5943), .I (g2233));
INVX1 gate4962(.O (g2801), .I (g2117));
INVX1 gate4963(.O (g5089), .I (g4840));
INVX1 gate4964(.O (I13406), .I (g8179));
INVX1 gate4965(.O (I9084), .I (g4886));
INVX1 gate4966(.O (g3738), .I (g3062));
INVX1 gate4967(.O (I13962), .I (g8451));
INVX1 gate4968(.O (I14786), .I (g9266));
INVX1 gate4969(.O (g7512), .I (g7148));
INVX1 gate4970(.O (g8025), .I (I12867));
INVX1 gate4971(.O (g9760), .I (g9454));
INVX1 gate4972(.O (I6294), .I (g2238));
INVX1 gate4973(.O (I17681), .I (g11608));
INVX1 gate4974(.O (g8425), .I (I13589));
INVX1 gate4975(.O (g3709), .I (I6870));
INVX1 gate4976(.O (g4124), .I (I7269));
INVX1 gate4977(.O (g4324), .I (g4144));
INVX1 gate4978(.O (g2748), .I (I5812));
INVX1 gate4979(.O (g6562), .I (g5774));
INVX1 gate4980(.O (g7366), .I (I11746));
INVX1 gate4981(.O (g10164), .I (I15488));
INVX1 gate4982(.O (I11833), .I (g7077));
INVX1 gate4983(.O (I11049), .I (g6635));
INVX1 gate4984(.O (I15675), .I (g10133));
INVX1 gate4985(.O (g4469), .I (I7840));
INVX1 gate4986(.O (g5705), .I (I9248));
INVX1 gate4987(.O (g5471), .I (g4370));
INVX1 gate4988(.O (g2755), .I (I5833));
INVX1 gate4989(.O (g11185), .I (I16956));
INVX1 gate4990(.O (g7056), .I (I11249));
INVX1 gate4991(.O (I17730), .I (g11638));
INVX1 gate4992(.O (g3907), .I (I7076));
INVX1 gate4993(.O (g10891), .I (I16635));
INVX1 gate4994(.O (g2226), .I (g86));
INVX1 gate4995(.O (I6501), .I (g2578));
INVX1 gate4996(.O (I10090), .I (g5767));
INVX1 gate4997(.O (g6723), .I (I10716));
INVX1 gate4998(.O (I13048), .I (g8059));
INVX1 gate4999(.O (g6257), .I (I10030));
INVX1 gate5000(.O (I14090), .I (g8771));
INVX1 gate5001(.O (g11518), .I (I17563));
INVX1 gate5002(.O (g4177), .I (I7348));
INVX1 gate5003(.O (I6156), .I (g2119));
INVX1 gate5004(.O (g6101), .I (I9762));
INVX1 gate5005(.O (g7148), .I (I11397));
INVX1 gate5006(.O (g6817), .I (I10861));
INVX1 gate5007(.O (g7649), .I (I12258));
INVX1 gate5008(.O (g5948), .I (I9588));
INVX1 gate5009(.O (g6301), .I (I10162));
INVX1 gate5010(.O (g7348), .I (I11692));
INVX1 gate5011(.O (I6356), .I (g2459));
INVX1 gate5012(.O (g4377), .I (I7694));
INVX1 gate5013(.O (g4206), .I (I7435));
INVX1 gate5014(.O (I10651), .I (g6035));
INVX1 gate5015(.O (g3517), .I (I6702));
INVX1 gate5016(.O (g10575), .I (g10523));
INVX1 gate5017(.O (I14182), .I (g8788));
INVX1 gate5018(.O (I14672), .I (g9261));
INVX1 gate5019(.O (g7355), .I (I11713));
INVX1 gate5020(.O (g2045), .I (g1811));
INVX1 gate5021(.O (g7851), .I (g7479));
INVX1 gate5022(.O (I17549), .I (g11501));
INVX1 gate5023(.O (g3876), .I (I7061));
INVX1 gate5024(.O (g8131), .I (g8020));
INVX1 gate5025(.O (g10327), .I (I15771));
INVX1 gate5026(.O (g8331), .I (I13373));
INVX1 gate5027(.O (g2173), .I (I5120));
INVX1 gate5028(.O (I12120), .I (g7106));
INVX1 gate5029(.O (g2373), .I (g471));
INVX1 gate5030(.O (g4287), .I (I7546));
INVX1 gate5031(.O (I9276), .I (g5241));
INVX1 gate5032(.O (g10537), .I (I16178));
INVX1 gate5033(.O (I10331), .I (g6198));
INVX1 gate5034(.O (g7964), .I (g7651));
INVX1 gate5035(.O (g8635), .I (I13918));
INVX1 gate5036(.O (g6751), .I (I10762));
INVX1 gate5037(.O (I12562), .I (g7377));
INVX1 gate5038(.O (I8011), .I (g3820));
INVX1 gate5039(.O (I11947), .I (g6905));
INVX1 gate5040(.O (g8105), .I (g7992));
INVX1 gate5041(.O (g2169), .I (g42));
INVX1 gate5042(.O (I5395), .I (g892));
INVX1 gate5043(.O (I14449), .I (g8973));
INVX1 gate5044(.O (g10283), .I (g10166));
INVX1 gate5045(.O (g2369), .I (g617));
INVX1 gate5046(.O (I5913), .I (g2169));
INVX1 gate5047(.O (I11106), .I (g6667));
INVX1 gate5048(.O (g8487), .I (g8350));
INVX1 gate5049(.O (g2602), .I (I5707));
INVX1 gate5050(.O (I11605), .I (g6834));
INVX1 gate5051(.O (g4199), .I (I7414));
INVX1 gate5052(.O (g6585), .I (I10541));
INVX1 gate5053(.O (g2007), .I (g936));
INVX1 gate5054(.O (g5773), .I (I9359));
INVX1 gate5055(.O (g10492), .I (I16111));
INVX1 gate5056(.O (g4399), .I (g3638));
INVX1 gate5057(.O (g7463), .I (g6921));
INVX1 gate5058(.O (g2407), .I (g197));
INVX1 gate5059(.O (I6163), .I (g2547));
INVX1 gate5060(.O (g2920), .I (g2462));
INVX1 gate5061(.O (I14961), .I (g9769));
INVX1 gate5062(.O (g2578), .I (g1962));
INVX1 gate5063(.O (g2868), .I (I6010));
INVX1 gate5064(.O (g3214), .I (I6391));
INVX1 gate5065(.O (g4781), .I (I8147));
INVX1 gate5066(.O (g6041), .I (I9658));
INVX1 gate5067(.O (I6363), .I (g2459));
INVX1 gate5068(.O (I7202), .I (g2647));
INVX1 gate5069(.O (I15729), .I (g10254));
INVX1 gate5070(.O (I13812), .I (g8519));
INVX1 gate5071(.O (I9647), .I (g5148));
INVX1 gate5072(.O (g4898), .I (I8259));
INVX1 gate5073(.O (g6441), .I (g6151));
INVX1 gate5074(.O (I13463), .I (g8156));
INVX1 gate5075(.O (g9451), .I (I14642));
INVX1 gate5076(.O (g4900), .I (I8265));
INVX1 gate5077(.O (I6432), .I (g2350));
INVX1 gate5078(.O (g11501), .I (I17522));
INVX1 gate5079(.O (g3110), .I (g2482));
INVX1 gate5080(.O (g11577), .I (I17613));
INVX1 gate5081(.O (g7279), .I (g6382));
INVX1 gate5082(.O (g5836), .I (g5320));
INVX1 gate5083(.O (g4510), .I (I7909));
INVX1 gate5084(.O (g11439), .I (I17368));
INVX1 gate5085(.O (g3663), .I (I6832));
INVX1 gate5086(.O (I12427), .I (g7636));
INVX1 gate5087(.O (g10091), .I (I15320));
INVX1 gate5088(.O (g9346), .I (I14543));
INVX1 gate5089(.O (I12366), .I (g7134));
INVX1 gate5090(.O (g2261), .I (g1713));
INVX1 gate5091(.O (g7619), .I (I12205));
INVX1 gate5092(.O (g7318), .I (I11602));
INVX1 gate5093(.O (g2793), .I (g2276));
INVX1 gate5094(.O (g4291), .I (g4013));
INVX1 gate5095(.O (g7872), .I (I12655));
INVX1 gate5096(.O (g11438), .I (I17365));
INVX1 gate5097(.O (g10174), .I (I15514));
INVX1 gate5098(.O (g10796), .I (I16500));
INVX1 gate5099(.O (I16664), .I (g10795));
INVX1 gate5100(.O (g9103), .I (g8892));
INVX1 gate5101(.O (I8080), .I (g3538));
INVX1 gate5102(.O (g2015), .I (g1107));
INVX1 gate5103(.O (g6368), .I (g5987));
INVX1 gate5104(.O (g8445), .I (I13633));
INVX1 gate5105(.O (I7776), .I (g3773));
INVX1 gate5106(.O (g7057), .I (I11252));
INVX1 gate5107(.O (g2227), .I (g95));
INVX1 gate5108(.O (g4344), .I (g3946));
INVX1 gate5109(.O (I5142), .I (g639));
INVX1 gate5110(.O (I7593), .I (g4142));
INVX1 gate5111(.O (I5248), .I (g1110));
INVX1 gate5112(.O (g7989), .I (I12805));
INVX1 gate5113(.O (I9224), .I (g5063));
INVX1 gate5114(.O (I15284), .I (g10034));
INVX1 gate5115(.O (g3762), .I (I6965));
INVX1 gate5116(.O (I12403), .I (g7611));
INVX1 gate5117(.O (I12547), .I (g7673));
INVX1 gate5118(.O (g4207), .I (I7438));
INVX1 gate5119(.O (g11083), .I (g10913));
INVX1 gate5120(.O (g11348), .I (g11276));
INVX1 gate5121(.O (g10390), .I (g10309));
INVX1 gate5122(.O (I16484), .I (g10770));
INVX1 gate5123(.O (g9732), .I (I14873));
INVX1 gate5124(.O (I5815), .I (g1994));
INVX1 gate5125(.O (I9120), .I (g5218));
INVX1 gate5126(.O (g11284), .I (g11208));
INVX1 gate5127(.O (I9320), .I (g5013));
INVX1 gate5128(.O (g2246), .I (g1810));
INVX1 gate5129(.O (g5822), .I (g5320));
INVX1 gate5130(.O (g4819), .I (g3354));
INVX1 gate5131(.O (g3877), .I (I7064));
INVX1 gate5132(.O (g9508), .I (g9271));
INVX1 gate5133(.O (I12226), .I (g7066));
INVX1 gate5134(.O (g8007), .I (I12843));
INVX1 gate5135(.O (I7264), .I (g3252));
INVX1 gate5136(.O (g11622), .I (I17684));
INVX1 gate5137(.O (g2203), .I (g677));
INVX1 gate5138(.O (g7686), .I (g7148));
INVX1 gate5139(.O (g10192), .I (I15554));
INVX1 gate5140(.O (I10620), .I (g5884));
INVX1 gate5141(.O (I5497), .I (g587));
INVX1 gate5142(.O (I6929), .I (g2846));
INVX1 gate5143(.O (I12481), .I (g7570));
INVX1 gate5144(.O (I13421), .I (g8200));
INVX1 gate5145(.O (I16200), .I (g10494));
INVX1 gate5146(.O (g8868), .I (I14176));
INVX1 gate5147(.O (I5960), .I (g2239));
INVX1 gate5148(.O (I7360), .I (g4081));
INVX1 gate5149(.O (I14097), .I (g8773));
INVX1 gate5150(.O (I9617), .I (g5405));
INVX1 gate5151(.O (g6856), .I (I10924));
INVX1 gate5152(.O (g6411), .I (g6135));
INVX1 gate5153(.O (g6734), .I (I10733));
INVX1 gate5154(.O (I9789), .I (g5401));
INVX1 gate5155(.O (I10343), .I (g6003));
INVX1 gate5156(.O (g8535), .I (I13744));
INVX1 gate5157(.O (I7450), .I (g3704));
INVX1 gate5158(.O (I10971), .I (g6344));
INVX1 gate5159(.O (g7321), .I (I11611));
INVX1 gate5160(.O (g8582), .I (I13825));
INVX1 gate5161(.O (g7670), .I (I12289));
INVX1 gate5162(.O (I17261), .I (g11346));
INVX1 gate5163(.O (g4215), .I (I7462));
INVX1 gate5164(.O (I7996), .I (g3462));
INVX1 gate5165(.O (g11653), .I (I17761));
INVX1 gate5166(.O (g2502), .I (I5579));
INVX1 gate5167(.O (g4886), .I (I8231));
INVX1 gate5168(.O (g4951), .I (I8320));
INVX1 gate5169(.O (I16799), .I (g11017));
INVX1 gate5170(.O (g7232), .I (I11472));
INVX1 gate5171(.O (I12490), .I (g7637));
INVX1 gate5172(.O (g10553), .I (I16220));
INVX1 gate5173(.O (g8015), .I (I12857));
INVX1 gate5174(.O (I15415), .I (g10075));
INVX1 gate5175(.O (g5895), .I (g5361));
INVX1 gate5176(.O (g7938), .I (g7403));
INVX1 gate5177(.O (I8126), .I (g3662));
INVX1 gate5178(.O (g7813), .I (I12604));
INVX1 gate5179(.O (I5979), .I (g2543));
INVX1 gate5180(.O (g4314), .I (g4013));
INVX1 gate5181(.O (I5218), .I (g1104));
INVX1 gate5182(.O (g5062), .I (g4840));
INVX1 gate5183(.O (I13788), .I (g8517));
INVX1 gate5184(.O (g9347), .I (I14546));
INVX1 gate5185(.O (I12376), .I (g7195));
INVX1 gate5186(.O (g10326), .I (I15768));
INVX1 gate5187(.O (g5620), .I (g4417));
INVX1 gate5188(.O (g7909), .I (g7664));
INVX1 gate5189(.O (g2689), .I (g2038));
INVX1 gate5190(.O (I12103), .I (g6859));
INVX1 gate5191(.O (I11829), .I (g7213));
INVX1 gate5192(.O (g6863), .I (g6740));
INVX1 gate5193(.O (I16184), .I (g10484));
INVX1 gate5194(.O (I16805), .I (g10904));
INVX1 gate5195(.O (g10536), .I (I16175));
INVX1 gate5196(.O (g8664), .I (I13949));
INVX1 gate5197(.O (g10040), .I (I15247));
INVX1 gate5198(.O (I10412), .I (g5821));
INVX1 gate5199(.O (I12354), .I (g7143));
INVX1 gate5200(.O (g2216), .I (g41));
INVX1 gate5201(.O (g9533), .I (I14684));
INVX1 gate5202(.O (g6713), .I (I10698));
INVX1 gate5203(.O (I14412), .I (g8939));
INVX1 gate5204(.O (g7519), .I (g6956));
INVX1 gate5205(.O (I13828), .I (g8488));
INVX1 gate5206(.O (g10904), .I (I16664));
INVX1 gate5207(.O (g2028), .I (g1703));
INVX1 gate5208(.O (I14133), .I (g8772));
INVX1 gate5209(.O (g10252), .I (g10137));
INVX1 gate5210(.O (g8721), .I (g8582));
INVX1 gate5211(.O (g6569), .I (I10499));
INVX1 gate5212(.O (g10621), .I (I16298));
INVX1 gate5213(.O (g7606), .I (I12168));
INVX1 gate5214(.O (I6894), .I (g2813));
INVX1 gate5215(.O (I13344), .I (g8121));
INVX1 gate5216(.O (I10228), .I (g6113));
INVX1 gate5217(.O (g2247), .I (I5258));
INVX1 gate5218(.O (I14228), .I (g8797));
INVX1 gate5219(.O (g4336), .I (g4130));
INVX1 gate5220(.O (g3394), .I (I6598));
INVX1 gate5221(.O (I5830), .I (g2067));
INVX1 gate5222(.O (g2564), .I (g1814));
INVX1 gate5223(.O (g7687), .I (I12318));
INVX1 gate5224(.O (g4768), .I (I8126));
INVX1 gate5225(.O (g11576), .I (I17610));
INVX1 gate5226(.O (I10716), .I (g6093));
INVX1 gate5227(.O (I13682), .I (g8310));
INVX1 gate5228(.O (g3731), .I (I6911));
INVX1 gate5229(.O (I15554), .I (g10088));
INVX1 gate5230(.O (g2826), .I (g2163));
INVX1 gate5231(.O (I6661), .I (g2752));
INVX1 gate5232(.O (g6688), .I (I10655));
INVX1 gate5233(.O (I11173), .I (g6500));
INVX1 gate5234(.O (g10183), .I (g10042));
INVX1 gate5235(.O (g6857), .I (I10927));
INVX1 gate5236(.O (g5192), .I (g4640));
INVX1 gate5237(.O (g5085), .I (g4377));
INVX1 gate5238(.O (I5221), .I (g1407));
INVX1 gate5239(.O (g9820), .I (I14961));
INVX1 gate5240(.O (g4943), .I (I8311));
INVX1 gate5241(.O (I12190), .I (g7268));
INVX1 gate5242(.O (I7674), .I (g3352));
INVX1 gate5243(.O (g11200), .I (g11112));
INVX1 gate5244(.O (g10062), .I (I15284));
INVX1 gate5245(.O (g3705), .I (g3113));
INVX1 gate5246(.O (I16214), .I (g10500));
INVX1 gate5247(.O (I17271), .I (g11388));
INVX1 gate5248(.O (I12520), .I (g7415));
INVX1 gate5249(.O (g2638), .I (I5751));
INVX1 gate5250(.O (g4065), .I (g2794));
INVX1 gate5251(.O (I8161), .I (g3637));
INVX1 gate5252(.O (g4887), .I (I8234));
INVX1 gate5253(.O (g4228), .I (g3914));
INVX1 gate5254(.O (g4322), .I (I7593));
INVX1 gate5255(.O (g7570), .I (I12032));
INVX1 gate5256(.O (g2108), .I (I4992));
INVX1 gate5257(.O (g5941), .I (I9571));
INVX1 gate5258(.O (I14379), .I (g8961));
INVX1 gate5259(.O (g2609), .I (I5728));
INVX1 gate5260(.O (g4934), .I (g4243));
INVX1 gate5261(.O (g7341), .I (I11671));
INVX1 gate5262(.O (I11029), .I (g6485));
INVX1 gate5263(.O (g10851), .I (I16553));
INVX1 gate5264(.O (g10872), .I (I16586));
INVX1 gate5265(.O (g11052), .I (I16817));
INVX1 gate5266(.O (I5932), .I (g2539));
INVX1 gate5267(.O (I10958), .I (g6559));
INVX1 gate5268(.O (g6400), .I (I10308));
INVX1 gate5269(.O (I14112), .I (g8777));
INVX1 gate5270(.O (I10378), .I (g6244));
INVX1 gate5271(.O (g7525), .I (I11921));
INVX1 gate5272(.O (I7680), .I (g3736));
INVX1 gate5273(.O (I14958), .I (g9767));
INVX1 gate5274(.O (g2883), .I (I6037));
INVX1 gate5275(.O (g8671), .I (I13956));
INVX1 gate5276(.O (I6484), .I (g2073));
INVX1 gate5277(.O (I6439), .I (g2352));
INVX1 gate5278(.O (I9915), .I (g5304));
INVX1 gate5279(.O (g3254), .I (g2322));
INVX1 gate5280(.O (g9775), .I (g9474));
INVX1 gate5281(.O (I17736), .I (g11640));
INVX1 gate5282(.O (I15798), .I (g10281));
INVX1 gate5283(.O (g3814), .I (g3228));
INVX1 gate5284(.O (g5708), .I (I9253));
INVX1 gate5285(.O (I10096), .I (g5794));
INVX1 gate5286(.O (g2217), .I (I5192));
INVX1 gate5287(.O (g2758), .I (I5840));
INVX1 gate5288(.O (g5520), .I (I8943));
INVX1 gate5289(.O (I14944), .I (g9454));
INVX1 gate5290(.O (I17198), .I (g11319));
INVX1 gate5291(.O (I15184), .I (g9974));
INVX1 gate5292(.O (g4096), .I (I7236));
INVX1 gate5293(.O (g8564), .I (I13785));
INVX1 gate5294(.O (g3038), .I (g1982));
INVX1 gate5295(.O (g4496), .I (I7889));
INVX1 gate5296(.O (I8303), .I (g4784));
INVX1 gate5297(.O (g11184), .I (I16953));
INVX1 gate5298(.O (g5252), .I (g4640));
INVX1 gate5299(.O (g7607), .I (I12171));
INVX1 gate5300(.O (I17528), .I (g11487));
INVX1 gate5301(.O (I6702), .I (g2801));
INVX1 gate5302(.O (g3773), .I (I6996));
INVX1 gate5303(.O (g5812), .I (g5320));
INVX1 gate5304(.O (g3009), .I (g2135));
INVX1 gate5305(.O (I14681), .I (g9110));
INVX1 gate5306(.O (g2165), .I (I5098));
INVX1 gate5307(.O (g6183), .I (g5320));
INVX1 gate5308(.O (g2571), .I (g1822));
INVX1 gate5309(.O (g7659), .I (I12274));
INVX1 gate5310(.O (g2861), .I (I6001));
INVX1 gate5311(.O (g7358), .I (I11722));
INVX1 gate5312(.O (g4195), .I (I7402));
INVX1 gate5313(.O (g5176), .I (g4682));
INVX1 gate5314(.O (g6220), .I (g5446));
INVX1 gate5315(.O (I5716), .I (g2068));
INVX1 gate5316(.O (g10574), .I (I16239));
INVX1 gate5317(.O (I17764), .I (g11651));
INVX1 gate5318(.O (I5149), .I (g1453));
INVX1 gate5319(.O (g4395), .I (I7732));
INVX1 gate5320(.O (g10047), .I (I15266));
INVX1 gate5321(.O (g4337), .I (g4144));
INVX1 gate5322(.O (g4913), .I (I8285));
INVX1 gate5323(.O (I17365), .I (g11380));
INVX1 gate5324(.O (I14802), .I (g9666));
INVX1 gate5325(.O (g10205), .I (g10176));
INVX1 gate5326(.O (g2055), .I (g1950));
INVX1 gate5327(.O (g3769), .I (I6982));
INVX1 gate5328(.O (g10912), .I (I16688));
INVX1 gate5329(.O (g10311), .I (g10242));
INVX1 gate5330(.O (g2455), .I (g826));
INVX1 gate5331(.O (g9739), .I (I14884));
INVX1 gate5332(.O (g2827), .I (g2164));
INVX1 gate5333(.O (I6952), .I (g2867));
INVX1 gate5334(.O (I14793), .I (g9269));
INVX1 gate5335(.O (g3212), .I (I6385));
INVX1 gate5336(.O (I9402), .I (g5107));
INVX1 gate5337(.O (I12339), .I (g7054));
INVX1 gate5338(.O (I8240), .I (g4380));
INVX1 gate5339(.O (g1975), .I (g622));
INVX1 gate5340(.O (I5198), .I (g143));
INVX1 gate5341(.O (I12296), .I (g7236));
INVX1 gate5342(.O (g7311), .I (I11581));
INVX1 gate5343(.O (g2774), .I (g2276));
INVX1 gate5344(.O (I6616), .I (g3186));
INVX1 gate5345(.O (g3967), .I (g3247));
INVX1 gate5346(.O (I17161), .I (g11314));
INVX1 gate5347(.O (g6588), .I (I10546));
INVX1 gate5348(.O (I4935), .I (g585));
INVX1 gate5349(.O (I12644), .I (g7729));
INVX1 gate5350(.O (g2846), .I (I5970));
INVX1 gate5351(.O (I9762), .I (g5276));
INVX1 gate5352(.O (I10549), .I (g6184));
INVX1 gate5353(.O (g9079), .I (g8892));
INVX1 gate5354(.O (I13648), .I (g8376));
INVX1 gate5355(.O (g10051), .I (I15272));
INVX1 gate5356(.O (I14690), .I (g9150));
INVX1 gate5357(.O (g6161), .I (I9886));
INVX1 gate5358(.O (I14549), .I (g9262));
INVX1 gate5359(.O (g7615), .I (I12193));
INVX1 gate5360(.O (g6361), .I (g5867));
INVX1 gate5361(.O (g2196), .I (g91));
INVX1 gate5362(.O (g4266), .I (g3688));
INVX1 gate5363(.O (I7600), .I (g4159));
INVX1 gate5364(.O (g9668), .I (g9490));
INVX1 gate5365(.O (g2396), .I (g1389));
INVX1 gate5366(.O (g10592), .I (I16261));
INVX1 gate5367(.O (I15400), .I (g10069));
INVX1 gate5368(.O (g2803), .I (g2154));
INVX1 gate5369(.O (g5733), .I (I9287));
INVX1 gate5370(.O (I17225), .I (g11298));
INVX1 gate5371(.O (g11400), .I (I17243));
INVX1 gate5372(.O (g6051), .I (I9680));
INVX1 gate5373(.O (I11770), .I (g7202));
INVX1 gate5374(.O (g5270), .I (g4367));
INVX1 gate5375(.O (g7374), .I (I11752));
INVX1 gate5376(.O (I11563), .I (g6819));
INVX1 gate5377(.O (I8116), .I (g3627));
INVX1 gate5378(.O (g6127), .I (I9826));
INVX1 gate5379(.O (g6451), .I (I10381));
INVX1 gate5380(.O (g8758), .I (I14055));
INVX1 gate5381(.O (g8066), .I (I12916));
INVX1 gate5382(.O (g8589), .I (I13834));
INVX1 gate5383(.O (I15329), .I (g9995));
INVX1 gate5384(.O (g7985), .I (I12799));
INVX1 gate5385(.O (I17258), .I (g11345));
INVX1 gate5386(.O (g4142), .I (I7288));
INVX1 gate5387(.O (g2509), .I (I5588));
INVX1 gate5388(.O (I16407), .I (g10696));
INVX1 gate5389(.O (I15539), .I (g10069));
INVX1 gate5390(.O (I6546), .I (g2987));
INVX1 gate5391(.O (g5073), .I (g4840));
INVX1 gate5392(.O (g10350), .I (I15814));
INVX1 gate5393(.O (g11207), .I (I16982));
INVX1 gate5394(.O (g1984), .I (g758));
INVX1 gate5395(.O (I10317), .I (g6003));
INVX1 gate5396(.O (g7284), .I (I11528));
INVX1 gate5397(.O (g11539), .I (g11519));
INVX1 gate5398(.O (g6146), .I (I9863));
INVX1 gate5399(.O (g10820), .I (I16528));
INVX1 gate5400(.O (g4081), .I (I7210));
INVX1 gate5401(.O (g7545), .I (I11967));
INVX1 gate5402(.O (g9356), .I (I14573));
INVX1 gate5403(.O (g8571), .I (I13806));
INVX1 gate5404(.O (I8147), .I (g3633));
INVX1 gate5405(.O (g2662), .I (g2014));
INVX1 gate5406(.O (g5124), .I (g4596));
INVX1 gate5407(.O (g2018), .I (g1336));
INVX1 gate5408(.O (g5980), .I (I9594));
INVX1 gate5409(.O (g2067), .I (g108));
INVX1 gate5410(.O (g7380), .I (g7279));
INVX1 gate5411(.O (g8448), .I (I13642));
INVX1 gate5412(.O (g6103), .I (I9766));
INVX1 gate5413(.O (I10129), .I (g5688));
INVX1 gate5414(.O (I9930), .I (g5317));
INVX1 gate5415(.O (I11767), .I (g7201));
INVX1 gate5416(.O (I11794), .I (g7188));
INVX1 gate5417(.O (g8711), .I (g8677));
INVX1 gate5418(.O (g7591), .I (I12103));
INVX1 gate5419(.O (g6303), .I (I10168));
INVX1 gate5420(.O (g2418), .I (I5497));
INVX1 gate5421(.O (I11845), .I (g6869));
INVX1 gate5422(.O (g5069), .I (g4368));
INVX1 gate5423(.O (I13794), .I (g8472));
INVX1 gate5424(.O (I10057), .I (g5741));
INVX1 gate5425(.O (g4726), .I (g3546));
INVX1 gate5426(.O (g2994), .I (g2057));
INVX1 gate5427(.O (g5469), .I (I8880));
INVX1 gate5428(.O (g7853), .I (I12652));
INVX1 gate5429(.O (g4354), .I (I7639));
INVX1 gate5430(.O (I5258), .I (g67));
INVX1 gate5431(.O (g7020), .I (I11159));
INVX1 gate5432(.O (I5818), .I (g2098));
INVX1 gate5433(.O (g8133), .I (I13002));
INVX1 gate5434(.O (g8333), .I (I13379));
INVX1 gate5435(.O (g7420), .I (I11804));
INVX1 gate5436(.O (I15241), .I (g10013));
INVX1 gate5437(.O (I11898), .I (g6896));
INVX1 gate5438(.O (g5177), .I (g4596));
INVX1 gate5439(.O (g6732), .I (I10729));
INVX1 gate5440(.O (I12867), .I (g7638));
INVX1 gate5441(.O (I17657), .I (g11598));
INVX1 gate5442(.O (I13633), .I (g8346));
INVX1 gate5443(.O (g11241), .I (g11112));
INVX1 gate5444(.O (I16206), .I (g10453));
INVX1 gate5445(.O (I10299), .I (g6243));
INVX1 gate5446(.O (g2256), .I (I5279));
INVX1 gate5447(.O (I11191), .I (g6514));
INVX1 gate5448(.O (I11719), .I (g7029));
INVX1 gate5449(.O (g7559), .I (I12009));
INVX1 gate5450(.O (I14323), .I (g8817));
INVX1 gate5451(.O (g10691), .I (I16360));
INVX1 gate5452(.O (g7794), .I (I12547));
INVX1 gate5453(.O (I7076), .I (g2985));
INVX1 gate5454(.O (I13191), .I (g8132));
INVX1 gate5455(.O (I14299), .I (g8810));
INVX1 gate5456(.O (I7889), .I (g3373));
INVX1 gate5457(.O (g8196), .I (I13125));
INVX1 gate5458(.O (g6944), .I (I11082));
INVX1 gate5459(.O (g8803), .I (I14130));
INVX1 gate5460(.O (I6277), .I (g1206));
INVX1 gate5461(.O (g6072), .I (g4977));
INVX1 gate5462(.O (I15771), .I (g10250));
INVX1 gate5463(.O (I9237), .I (g5205));
INVX1 gate5464(.O (I17337), .I (g11363));
INVX1 gate5465(.O (g2181), .I (I5142));
INVX1 gate5466(.O (g8538), .I (I13747));
INVX1 gate5467(.O (g2381), .I (g1368));
INVX1 gate5468(.O (g9432), .I (g9313));
INVX1 gate5469(.O (I15235), .I (g9968));
INVX1 gate5470(.O (I6789), .I (g2748));
INVX1 gate5471(.O (I16114), .I (g10387));
INVX1 gate5472(.O (g4783), .I (g3829));
INVX1 gate5473(.O (g6043), .I (I9662));
INVX1 gate5474(.O (I12910), .I (g7922));
INVX1 gate5475(.O (I7375), .I (g4062));
INVX1 gate5476(.O (g2847), .I (I5973));
INVX1 gate5477(.O (g8780), .I (I14077));
INVX1 gate5478(.O (g6443), .I (g6157));
INVX1 gate5479(.O (I12202), .I (g6983));
INVX1 gate5480(.O (g8509), .I (g8366));
INVX1 gate5481(.O (g9453), .I (g9100));
INVX1 gate5482(.O (g4112), .I (g2994));
INVX1 gate5483(.O (g7905), .I (g7450));
INVX1 gate5484(.O (g2197), .I (g101));
INVX1 gate5485(.O (I7651), .I (g3332));
INVX1 gate5486(.O (g4312), .I (g4144));
INVX1 gate5487(.O (I8820), .I (g4473));
INVX1 gate5488(.O (I11440), .I (g6577));
INVX1 gate5489(.O (g10929), .I (g10827));
INVX1 gate5490(.O (I12496), .I (g7724));
INVX1 gate5491(.O (g2021), .I (g1341));
INVX1 gate5492(.O (I9194), .I (g5236));
INVX1 gate5493(.O (g7628), .I (I12226));
INVX1 gate5494(.O (I9394), .I (g5195));
INVX1 gate5495(.O (g6116), .I (I9801));
INVX1 gate5496(.O (g2421), .I (g1374));
INVX1 gate5497(.O (g7630), .I (I12232));
INVX1 gate5498(.O (g4001), .I (g3200));
INVX1 gate5499(.O (I12978), .I (g8040));
INVX1 gate5500(.O (I14232), .I (g8800));
INVX1 gate5501(.O (g10928), .I (g10827));
INVX1 gate5502(.O (g8067), .I (I12919));
INVX1 gate5503(.O (I9731), .I (g5255));
INVX1 gate5504(.O (g5898), .I (g5361));
INVX1 gate5505(.O (g8418), .I (I13568));
INVX1 gate5506(.O (g6434), .I (I10352));
INVX1 gate5507(.O (g4676), .I (g3354));
INVX1 gate5508(.O (g5900), .I (I9531));
INVX1 gate5509(.O (g6565), .I (g5790));
INVX1 gate5510(.O (I5821), .I (g2101));
INVX1 gate5511(.O (I6299), .I (g2242));
INVX1 gate5512(.O (I11926), .I (g6900));
INVX1 gate5513(.O (g8290), .I (I13224));
INVX1 gate5514(.O (I12986), .I (g8042));
INVX1 gate5515(.O (g4129), .I (I7280));
INVX1 gate5516(.O (g5797), .I (I9399));
INVX1 gate5517(.O (g4329), .I (g4144));
INVX1 gate5518(.O (I14697), .I (g9260));
INVX1 gate5519(.O (g4761), .I (g3440));
INVX1 gate5520(.O (g11515), .I (g11490));
INVX1 gate5521(.O (I7384), .I (g4082));
INVX1 gate5522(.O (I13612), .I (g8325));
INVX1 gate5523(.O (g5245), .I (g4369));
INVX1 gate5524(.O (I7339), .I (g4004));
INVX1 gate5525(.O (I13099), .I (g7927));
INVX1 gate5526(.O (I12384), .I (g7212));
INVX1 gate5527(.O (g8093), .I (I12948));
INVX1 gate5528(.O (I13388), .I (g8230));
INVX1 gate5529(.O (g6681), .I (g5830));
INVX1 gate5530(.O (I11701), .I (g7065));
INVX1 gate5531(.O (I11534), .I (g6917));
INVX1 gate5532(.O (g10787), .I (I16487));
INVX1 gate5533(.O (g5291), .I (g4384));
INVX1 gate5534(.O (g3392), .I (g3121));
INVX1 gate5535(.O (I11272), .I (g6546));
INVX1 gate5536(.O (g10282), .I (g10164));
INVX1 gate5537(.O (g7750), .I (I12415));
INVX1 gate5538(.O (g3485), .I (g2662));
INVX1 gate5539(.O (g2562), .I (g1383));
INVX1 gate5540(.O (g6697), .I (g5949));
INVX1 gate5541(.O (g5144), .I (g4682));
INVX1 gate5542(.O (g4592), .I (g3829));
INVX1 gate5543(.O (g6914), .I (I11024));
INVX1 gate5544(.O (I17444), .I (g11446));
INVX1 gate5545(.O (g5344), .I (I8811));
INVX1 gate5546(.O (g6210), .I (g5205));
INVX1 gate5547(.O (I12150), .I (g7074));
INVX1 gate5548(.O (g4746), .I (I8098));
INVX1 gate5549(.O (g8181), .I (I13096));
INVX1 gate5550(.O (g10827), .I (I16543));
INVX1 gate5551(.O (g6596), .I (I10566));
INVX1 gate5552(.O (I6738), .I (g3113));
INVX1 gate5553(.O (g4221), .I (g3914));
INVX1 gate5554(.O (g8381), .I (I13489));
INVX1 gate5555(.O (g2101), .I (I4951));
INVX1 gate5556(.O (g2817), .I (I5919));
INVX1 gate5557(.O (g3941), .I (g3015));
INVX1 gate5558(.O (g7040), .I (I11207));
INVX1 gate5559(.O (g6413), .I (I10325));
INVX1 gate5560(.O (I10831), .I (g6710));
INVX1 gate5561(.O (g7440), .I (I11836));
INVX1 gate5562(.O (g8197), .I (I13128));
INVX1 gate5563(.O (g8700), .I (g8574));
INVX1 gate5564(.O (I10445), .I (g5770));
INVX1 gate5565(.O (I7523), .I (g4095));
INVX1 gate5566(.O (I11140), .I (g6448));
INVX1 gate5567(.O (I12196), .I (g7272));
INVX1 gate5568(.O (g2605), .I (I5716));
INVX1 gate5569(.O (g11441), .I (I17374));
INVX1 gate5570(.O (I9150), .I (g5012));
INVX1 gate5571(.O (I10499), .I (g6149));
INVX1 gate5572(.O (g8421), .I (I13577));
INVX1 gate5573(.O (g7123), .I (I11360));
INVX1 gate5574(.O (g5088), .I (I8456));
INVX1 gate5575(.O (g11206), .I (I16979));
INVX1 gate5576(.O (g7323), .I (I11617));
INVX1 gate5577(.O (I14499), .I (g8889));
INVX1 gate5578(.O (I6907), .I (g2994));
INVX1 gate5579(.O (I12526), .I (g7648));
INVX1 gate5580(.O (g10803), .I (g10708));
INVX1 gate5581(.O (I7205), .I (g2632));
INVX1 gate5582(.O (I9773), .I (g4934));
INVX1 gate5583(.O (I15759), .I (g10267));
INVX1 gate5584(.O (I11061), .I (g6641));
INVX1 gate5585(.O (I15725), .I (g10251));
INVX1 gate5586(.O (g5701), .I (I9240));
INVX1 gate5587(.O (g3708), .I (I6867));
INVX1 gate5588(.O (g4953), .I (I8324));
INVX1 gate5589(.O (g2751), .I (I5821));
INVX1 gate5590(.O (g3520), .I (g2779));
INVX1 gate5591(.O (g8950), .I (I14303));
INVX1 gate5592(.O (I16500), .I (g10711));
INVX1 gate5593(.O (g3219), .I (I6395));
INVX1 gate5594(.O (I6517), .I (g3271));
INVX1 gate5595(.O (I6690), .I (g2743));
INVX1 gate5596(.O (I9409), .I (g5013));
INVX1 gate5597(.O (I15114), .I (g9875));
INVX1 gate5598(.O (I5427), .I (g913));
INVX1 gate5599(.O (g4468), .I (I7837));
INVX1 gate5600(.O (I15082), .I (g9719));
INVX1 gate5601(.O (g6117), .I (I9804));
INVX1 gate5602(.O (I14989), .I (g9813));
INVX1 gate5603(.O (I17158), .I (g11312));
INVX1 gate5604(.O (g3252), .I (I6414));
INVX1 gate5605(.O (g10881), .I (I16613));
INVX1 gate5606(.O (I7104), .I (g3186));
INVX1 gate5607(.O (g11435), .I (I17356));
INVX1 gate5608(.O (I6876), .I (g2956));
INVX1 gate5609(.O (I9769), .I (g5287));
INVX1 gate5610(.O (g11082), .I (I16859));
INVX1 gate5611(.O (g3812), .I (g3228));
INVX1 gate5612(.O (I7099), .I (g3228));
INVX1 gate5613(.O (I12457), .I (g7559));
INVX1 gate5614(.O (I10924), .I (g6736));
INVX1 gate5615(.O (g5886), .I (g5361));
INVX1 gate5616(.O (g11107), .I (g10974));
INVX1 gate5617(.O (I9836), .I (g5405));
INVX1 gate5618(.O (I14080), .I (g8714));
INVX1 gate5619(.O (g7351), .I (I11701));
INVX1 gate5620(.O (g2041), .I (g1791));
INVX1 gate5621(.O (g7648), .I (I12255));
INVX1 gate5622(.O (g7530), .I (I11926));
INVX1 gate5623(.O (I11360), .I (g6351));
INVX1 gate5624(.O (g8562), .I (I13779));
INVX1 gate5625(.O (I15744), .I (g10261));
INVX1 gate5626(.O (I13360), .I (g8126));
INVX1 gate5627(.O (I17353), .I (g11381));
INVX1 gate5628(.O (g3405), .I (g3144));
INVX1 gate5629(.O (g5114), .I (I8506));
INVX1 gate5630(.O (I5403), .I (g636));
INVX1 gate5631(.O (g9778), .I (g9474));
INVX1 gate5632(.O (g5314), .I (g4387));
INVX1 gate5633(.O (I11447), .I (g6431));
INVX1 gate5634(.O (g11345), .I (I17158));
INVX1 gate5635(.O (g9894), .I (I15085));
INVX1 gate5636(.O (g8723), .I (g8585));
INVX1 gate5637(.O (g4716), .I (g3546));
INVX1 gate5638(.O (I11162), .I (g6479));
INVX1 gate5639(.O (I16613), .I (g10794));
INVX1 gate5640(.O (g11399), .I (I17240));
INVX1 gate5641(.O (g3765), .I (g3120));
INVX1 gate5642(.O (I10753), .I (g5814));
INVX1 gate5643(.O (I10461), .I (g5849));
INVX1 gate5644(.O (I5391), .I (g1101));
INVX1 gate5645(.O (g3911), .I (g3015));
INVX1 gate5646(.O (I9229), .I (g4954));
INVX1 gate5647(.O (g7010), .I (I11155));
INVX1 gate5648(.O (g6581), .I (I10531));
INVX1 gate5649(.O (g10890), .I (I16632));
INVX1 gate5650(.O (g5650), .I (I9111));
INVX1 gate5651(.O (g7410), .I (I11790));
INVX1 gate5652(.O (g9782), .I (I14933));
INVX1 gate5653(.O (g11398), .I (I17237));
INVX1 gate5654(.O (I15804), .I (g10283));
INVX1 gate5655(.O (I16947), .I (g11080));
INVX1 gate5656(.O (I5695), .I (g575));
INVX1 gate5657(.O (g10249), .I (g10135));
INVX1 gate5658(.O (g2168), .I (I5111));
INVX1 gate5659(.O (g2669), .I (g2015));
INVX1 gate5660(.O (g6060), .I (I9695));
INVX1 gate5661(.O (I16273), .I (g10559));
INVX1 gate5662(.O (g2368), .I (I5445));
INVX1 gate5663(.O (I11629), .I (g6914));
INVX1 gate5664(.O (g11652), .I (I17758));
INVX1 gate5665(.O (I9822), .I (g5219));
INVX1 gate5666(.O (g9661), .I (I14786));
INVX1 gate5667(.O (g4198), .I (I7411));
INVX1 gate5668(.O (g4747), .I (g3586));
INVX1 gate5669(.O (I11472), .I (g6488));
INVX1 gate5670(.O (I10736), .I (g6104));
INVX1 gate5671(.O (g4398), .I (g3914));
INVX1 gate5672(.O (I13451), .I (g8152));
INVX1 gate5673(.O (g3733), .I (I6917));
INVX1 gate5674(.O (I7444), .I (g3683));
INVX1 gate5675(.O (g10248), .I (g10134));
INVX1 gate5676(.O (g2772), .I (g2508));
INVX1 gate5677(.O (I7269), .I (g2851));
INVX1 gate5678(.O (I15263), .I (g9995));
INVX1 gate5679(.O (I10198), .I (g6118));
INVX1 gate5680(.O (I12300), .I (g7240));
INVX1 gate5681(.O (g10552), .I (I16217));
INVX1 gate5682(.O (g8751), .I (g8632));
INVX1 gate5683(.O (I15332), .I (g10001));
INVX1 gate5684(.O (g10204), .I (g10174));
INVX1 gate5685(.O (g2743), .I (I5801));
INVX1 gate5686(.O (g4241), .I (g3664));
INVX1 gate5687(.O (g2890), .I (I6052));
INVX1 gate5688(.O (g5768), .I (I9352));
INVX1 gate5689(.O (I10843), .I (g6723));
INVX1 gate5690(.O (g8585), .I (I13828));
INVX1 gate5691(.O (I5858), .I (g2529));
INVX1 gate5692(.O (g5594), .I (I9016));
INVX1 gate5693(.O (I14528), .I (g9270));
INVX1 gate5694(.O (g3473), .I (I6676));
INVX1 gate5695(.O (g7278), .I (I11524));
INVX1 gate5696(.O (I14330), .I (g8819));
INVX1 gate5697(.O (g9526), .I (g9256));
INVX1 gate5698(.O (I4938), .I (g261));
INVX1 gate5699(.O (I8250), .I (g4589));
INVX1 gate5700(.O (I11071), .I (g6656));
INVX1 gate5701(.O (I15406), .I (g10065));
INVX1 gate5702(.O (I15962), .I (g10405));
INVX1 gate5703(.O (g2011), .I (g976));
INVX1 gate5704(.O (g6995), .I (g6482));
INVX1 gate5705(.O (g7618), .I (I12202));
INVX1 gate5706(.O (g3980), .I (g3121));
INVX1 gate5707(.O (g8441), .I (I13621));
INVX1 gate5708(.O (g11406), .I (I17261));
INVX1 gate5709(.O (g5943), .I (I9581));
INVX1 gate5710(.O (g7343), .I (I11677));
INVX1 gate5711(.O (g2411), .I (I5494));
INVX1 gate5712(.O (I10132), .I (g5696));
INVX1 gate5713(.O (g10786), .I (I16484));
INVX1 gate5714(.O (g3069), .I (I6277));
INVX1 gate5715(.O (I13776), .I (g8513));
INVX1 gate5716(.O (I13785), .I (g8516));
INVX1 gate5717(.O (g1982), .I (g736));
INVX1 gate5718(.O (g4524), .I (g3946));
INVX1 gate5719(.O (g6294), .I (I10141));
INVX1 gate5720(.O (I15500), .I (g10051));
INVX1 gate5721(.O (I5251), .I (g1424));
INVX1 gate5722(.O (I6590), .I (g3186));
INVX1 gate5723(.O (g3540), .I (g3307));
INVX1 gate5724(.O (I7729), .I (g3757));
INVX1 gate5725(.O (g5887), .I (I9510));
INVX1 gate5726(.O (g10356), .I (I15832));
INVX1 gate5727(.O (I5047), .I (g1185));
INVX1 gate5728(.O (g5122), .I (g4682));
INVX1 gate5729(.O (g11500), .I (I17519));
INVX1 gate5730(.O (g6190), .I (g5426));
INVX1 gate5731(.O (g2074), .I (g1377));
INVX1 gate5732(.O (g4319), .I (g4144));
INVX1 gate5733(.O (g7693), .I (I12326));
INVX1 gate5734(.O (g11049), .I (I16808));
INVX1 gate5735(.O (I11950), .I (g6906));
INVX1 gate5736(.O (I16514), .I (g10717));
INVX1 gate5737(.O (g10826), .I (I16540));
INVX1 gate5738(.O (I9062), .I (g4759));
INVX1 gate5739(.O (g7334), .I (I11650));
INVX1 gate5740(.O (g10380), .I (I15864));
INVX1 gate5741(.O (g3206), .I (g2055));
INVX1 gate5742(.O (I13825), .I (g8488));
INVX1 gate5743(.O (I13370), .I (g8128));
INVX1 gate5744(.O (I9620), .I (g5189));
INVX1 gate5745(.O (g4258), .I (I7509));
INVX1 gate5746(.O (I16507), .I (g10712));
INVX1 gate5747(.O (g4352), .I (I7633));
INVX1 gate5748(.O (I11858), .I (g6888));
INVX1 gate5749(.O (g11048), .I (I16805));
INVX1 gate5750(.O (g4577), .I (I7984));
INVX1 gate5751(.O (g4867), .I (I8204));
INVX1 gate5752(.O (I14709), .I (g9267));
INVX1 gate5753(.O (g5033), .I (I8406));
INVX1 gate5754(.O (g10233), .I (g10187));
INVX1 gate5755(.O (g6156), .I (g5426));
INVX1 gate5756(.O (g4717), .I (g3829));
INVX1 gate5757(.O (I7014), .I (g2919));
INVX1 gate5758(.O (I12511), .I (g7733));
INVX1 gate5759(.O (g10182), .I (I15530));
INVX1 gate5760(.O (g7555), .I (I11989));
INVX1 gate5761(.O (g7804), .I (I12577));
INVX1 gate5762(.O (I7414), .I (g4156));
INVX1 gate5763(.O (I10087), .I (g5753));
INVX1 gate5764(.O (g9919), .I (I15114));
INVX1 gate5765(.O (g2080), .I (I4894));
INVX1 gate5766(.O (I7946), .I (g3417));
INVX1 gate5767(.O (I10258), .I (g6134));
INVX1 gate5768(.O (I14087), .I (g8770));
INVX1 gate5769(.O (g7792), .I (I12541));
INVX1 gate5770(.O (g2480), .I (I5561));
INVX1 gate5771(.O (I11367), .I (g6392));
INVX1 gate5772(.O (I11394), .I (g6621));
INVX1 gate5773(.O (g5096), .I (g4840));
INVX1 gate5774(.O (g6942), .I (I11076));
INVX1 gate5775(.O (g8890), .I (I14236));
INVX1 gate5776(.O (g2713), .I (g2042));
INVX1 gate5777(.O (I13367), .I (g8221));
INVX1 gate5778(.O (I13394), .I (g8137));
INVX1 gate5779(.O (g4211), .I (I7450));
INVX1 gate5780(.O (g4186), .I (I7375));
INVX1 gate5781(.O (g6704), .I (g5949));
INVX1 gate5782(.O (I17687), .I (g11610));
INVX1 gate5783(.O (g4386), .I (I7713));
INVX1 gate5784(.O (g10932), .I (g10827));
INVX1 gate5785(.O (I8929), .I (g4582));
INVX1 gate5786(.O (g5845), .I (g5320));
INVX1 gate5787(.O (g4975), .I (I8351));
INVX1 gate5788(.O (g2569), .I (I5695));
INVX1 gate5789(.O (I7513), .I (g4144));
INVX1 gate5790(.O (g8011), .I (I12853));
INVX1 gate5791(.O (I17752), .I (g11645));
INVX1 gate5792(.O (g5195), .I (g4453));
INVX1 gate5793(.O (g5395), .I (I8831));
INVX1 gate5794(.O (g5891), .I (g5361));
INVX1 gate5795(.O (I9842), .I (g5405));
INVX1 gate5796(.O (I17374), .I (g11411));
INVX1 gate5797(.O (g7113), .I (I11348));
INVX1 gate5798(.O (g11106), .I (g10974));
INVX1 gate5799(.O (g7313), .I (I11587));
INVX1 gate5800(.O (I11420), .I (g6417));
INVX1 gate5801(.O (g4426), .I (g3914));
INVX1 gate5802(.O (g10897), .I (g10827));
INVX1 gate5803(.O (I12916), .I (g7849));
INVX1 gate5804(.O (I10069), .I (g5787));
INVX1 gate5805(.O (g6954), .I (I11100));
INVX1 gate5806(.O (g6250), .I (I10009));
INVX1 gate5807(.O (g4170), .I (g3328));
INVX1 gate5808(.O (g6810), .I (I10840));
INVX1 gate5809(.O (g4614), .I (g3829));
INVX1 gate5810(.O (g9527), .I (I14668));
INVX1 gate5811(.O (g4370), .I (I7671));
INVX1 gate5812(.O (I12550), .I (g7675));
INVX1 gate5813(.O (I7378), .I (g4067));
INVX1 gate5814(.O (I10810), .I (g6539));
INVX1 gate5815(.O (I11318), .I (g6488));
INVX1 gate5816(.O (g4125), .I (I7272));
INVX1 gate5817(.O (I15371), .I (g9990));
INVX1 gate5818(.O (g6432), .I (g6146));
INVX1 gate5819(.O (g7908), .I (g7454));
INVX1 gate5820(.O (I13227), .I (g8264));
INVX1 gate5821(.O (g6053), .I (I9684));
INVX1 gate5822(.O (I14955), .I (g9765));
INVX1 gate5823(.O (I17669), .I (g11604));
INVX1 gate5824(.O (g8992), .I (I14397));
INVX1 gate5825(.O (g9764), .I (g9432));
INVX1 gate5826(.O (I16920), .I (g11084));
INVX1 gate5827(.O (g11033), .I (I16760));
INVX1 gate5828(.O (g3291), .I (g2161));
INVX1 gate5829(.O (I12307), .I (g7245));
INVX1 gate5830(.O (I5935), .I (g2174));
INVX1 gate5831(.O (I6844), .I (g2915));
INVX1 gate5832(.O (g6453), .I (g5817));
INVX1 gate5833(.O (I9854), .I (g5557));
INVX1 gate5834(.O (I14970), .I (g9732));
INVX1 gate5835(.O (g4280), .I (g4013));
INVX1 gate5836(.O (I7182), .I (g2645));
INVX1 gate5837(.O (I7288), .I (g2873));
INVX1 gate5838(.O (g4939), .I (I8303));
INVX1 gate5839(.O (I11540), .I (g6877));
INVX1 gate5840(.O (I5982), .I (g2510));
INVX1 gate5841(.O (g3144), .I (g2462));
INVX1 gate5842(.O (I11058), .I (g6641));
INVX1 gate5843(.O (I15795), .I (g10280));
INVX1 gate5844(.O (g3344), .I (I6528));
INVX1 gate5845(.O (I16121), .I (g10396));
INVX1 gate5846(.O (g6568), .I (g5797));
INVX1 gate5847(.O (I10171), .I (g5992));
INVX1 gate5848(.O (g4083), .I (I7216));
INVX1 gate5849(.O (g8080), .I (I12942));
INVX1 gate5850(.O (I4879), .I (g256));
INVX1 gate5851(.O (g4544), .I (g3880));
INVX1 gate5852(.O (g3207), .I (g2439));
INVX1 gate5853(.O (g8573), .I (I13812));
INVX1 gate5854(.O (I7916), .I (g3664));
INVX1 gate5855(.O (I7022), .I (g2941));
INVX1 gate5856(.O (I13203), .I (g8196));
INVX1 gate5857(.O (g8480), .I (I13682));
INVX1 gate5858(.O (g7776), .I (I12493));
INVX1 gate5859(.O (g2000), .I (g810));
INVX1 gate5860(.O (I7749), .I (g3764));
INVX1 gate5861(.O (I6557), .I (g3086));
INVX1 gate5862(.O (g8713), .I (g8684));
INVX1 gate5863(.O (I17525), .I (g11486));
INVX1 gate5864(.O (g2126), .I (g12));
INVX1 gate5865(.O (g4636), .I (I8036));
INVX1 gate5866(.O (I15514), .I (g10122));
INVX1 gate5867(.O (I17424), .I (g11424));
INVX1 gate5868(.O (g3694), .I (I6851));
INVX1 gate5869(.O (g6157), .I (I9880));
INVX1 gate5870(.O (I6071), .I (g2269));
INVX1 gate5871(.O (I14967), .I (g9763));
INVX1 gate5872(.O (I12773), .I (g7581));
INVX1 gate5873(.O (I16682), .I (g10799));
INVX1 gate5874(.O (I17558), .I (g11504));
INVX1 gate5875(.O (I15507), .I (g10047));
INVX1 gate5876(.O (g5081), .I (I8449));
INVX1 gate5877(.O (I12942), .I (g7982));
INVX1 gate5878(.O (g3088), .I (I6294));
INVX1 gate5879(.O (g5815), .I (I9421));
INVX1 gate5880(.O (g8569), .I (I13800));
INVX1 gate5881(.O (g4306), .I (g3586));
INVX1 gate5882(.O (g7965), .I (I12759));
INVX1 gate5883(.O (I12268), .I (g7107));
INVX1 gate5884(.O (g5481), .I (I8900));
INVX1 gate5885(.O (g11507), .I (I17540));
INVX1 gate5886(.O (I12156), .I (g6878));
INVX1 gate5887(.O (g4790), .I (g3337));
INVX1 gate5888(.O (I12655), .I (g7402));
INVX1 gate5889(.O (g5692), .I (I9221));
INVX1 gate5890(.O (I15421), .I (g10083));
INVX1 gate5891(.O (g1964), .I (g114));
INVX1 gate5892(.O (g10387), .I (g10357));
INVX1 gate5893(.O (g97), .I (I4780));
INVX1 gate5894(.O (g7264), .I (I11501));
INVX1 gate5895(.O (I12180), .I (g7263));
INVX1 gate5896(.O (g10620), .I (I16295));
INVX1 gate5897(.O (g4187), .I (I7378));
INVX1 gate5898(.O (g4061), .I (I7182));
INVX1 gate5899(.O (g10148), .I (g10121));
INVX1 gate5900(.O (g11421), .I (I17318));
INVX1 gate5901(.O (g4387), .I (I7716));
INVX1 gate5902(.O (g4461), .I (g3829));
INVX1 gate5903(.O (I6955), .I (g2871));
INVX1 gate5904(.O (g7360), .I (I11728));
INVX1 gate5905(.O (g11163), .I (I16920));
INVX1 gate5906(.O (g10104), .I (I15338));
INVX1 gate5907(.O (I11146), .I (g6439));
INVX1 gate5908(.O (g4756), .I (g3440));
INVX1 gate5909(.O (I17713), .I (g11621));
INVX1 gate5910(.O (I13738), .I (g8295));
INVX1 gate5911(.O (I13645), .I (g8379));
INVX1 gate5912(.O (g8688), .I (g8507));
INVX1 gate5913(.O (I12335), .I (g7133));
INVX1 gate5914(.O (g7521), .I (I11901));
INVX1 gate5915(.O (g10343), .I (I15795));
INVX1 gate5916(.O (I14010), .I (g8642));
INVX1 gate5917(.O (I14918), .I (g9535));
INVX1 gate5918(.O (g8976), .I (I14349));
INVX1 gate5919(.O (g2608), .I (I5725));
INVX1 gate5920(.O (I9829), .I (g5013));
INVX1 gate5921(.O (I16760), .I (g10888));
INVX1 gate5922(.O (g2220), .I (g104));
INVX1 gate5923(.O (g4427), .I (g3638));
INVX1 gate5924(.O (I12930), .I (g7896));
INVX1 gate5925(.O (g7450), .I (g7148));
INVX1 gate5926(.O (I12993), .I (g8044));
INVX1 gate5927(.O (I15473), .I (g10087));
INVX1 gate5928(.O (I13290), .I (g8254));
INVX1 gate5929(.O (g2779), .I (g1974));
INVX1 gate5930(.O (I6150), .I (g2122));
INVX1 gate5931(.O (g9987), .I (I15187));
INVX1 gate5932(.O (g11541), .I (g11519));
INVX1 gate5933(.O (I17610), .I (g11549));
INVX1 gate5934(.O (I11698), .I (g7057));
INVX1 gate5935(.O (g4200), .I (I7417));
INVX1 gate5936(.O (g9771), .I (g9432));
INVX1 gate5937(.O (I12694), .I (g7374));
INVX1 gate5938(.O (I12838), .I (g7682));
INVX1 gate5939(.O (g11473), .I (I17456));
INVX1 gate5940(.O (g2023), .I (g1357));
INVX1 gate5941(.O (I10078), .I (g5729));
INVX1 gate5942(.O (I17255), .I (g11344));
INVX1 gate5943(.O (g4514), .I (g3946));
INVX1 gate5944(.O (I10598), .I (g5874));
INVX1 gate5945(.O (g5783), .I (I9377));
INVX1 gate5946(.O (g4003), .I (g3144));
INVX1 gate5947(.O (g7724), .I (I12357));
INVX1 gate5948(.O (I15359), .I (g10019));
INVX1 gate5949(.O (I6409), .I (g2356));
INVX1 gate5950(.O (g8126), .I (I12989));
INVX1 gate5951(.O (I7719), .I (g3752));
INVX1 gate5952(.O (g5112), .I (g4682));
INVX1 gate5953(.O (g7379), .I (g6863));
INVX1 gate5954(.O (g5218), .I (I8647));
INVX1 gate5955(.O (g8326), .I (I13360));
INVX1 gate5956(.O (I17188), .I (g11313));
INVX1 gate5957(.O (I17124), .I (g11232));
INVX1 gate5958(.O (g5267), .I (I8711));
INVX1 gate5959(.O (I17678), .I (g11607));
INVX1 gate5960(.O (I11427), .I (g6573));
INVX1 gate5961(.O (I12487), .I (g7723));
INVX1 gate5962(.O (I15829), .I (g10203));
INVX1 gate5963(.O (I13427), .I (g8241));
INVX1 gate5964(.O (g9892), .I (I15079));
INVX1 gate5965(.O (I8039), .I (g3506));
INVX1 gate5966(.O (I7752), .I (g3407));
INVX1 gate5967(.O (g4763), .I (g3586));
INVX1 gate5968(.O (I12502), .I (g7726));
INVX1 gate5969(.O (g4191), .I (I7390));
INVX1 gate5970(.O (I11632), .I (g6931));
INVX1 gate5971(.O (g7878), .I (g7479));
INVX1 gate5972(.O (g10850), .I (I16550));
INVX1 gate5973(.O (g8760), .I (g8670));
INVX1 gate5974(.O (g11434), .I (I17353));
INVX1 gate5975(.O (g4391), .I (g3638));
INVX1 gate5976(.O (g1989), .I (g770));
INVX1 gate5977(.O (I10322), .I (g6193));
INVX1 gate5978(.O (g7289), .I (I11543));
INVX1 gate5979(.O (g7777), .I (I12496));
INVX1 gate5980(.O (g7658), .I (I12271));
INVX1 gate5981(.O (g5401), .I (I8839));
INVX1 gate5982(.O (g3408), .I (g3108));
INVX1 gate5983(.O (I10159), .I (g5936));
INVX1 gate5984(.O (g10133), .I (g10064));
INVX1 gate5985(.O (g5676), .I (I9185));
INVX1 gate5986(.O (g2451), .I (g248));
INVX1 gate5987(.O (I10901), .I (g6620));
INVX1 gate5988(.O (g4637), .I (I8039));
INVX1 gate5989(.O (I12279), .I (g7225));
INVX1 gate5990(.O (I5348), .I (g746));
INVX1 gate5991(.O (g3336), .I (I6523));
INVX1 gate5992(.O (I15344), .I (g10025));
INVX1 gate5993(.O (g6778), .I (g5987));
INVX1 gate5994(.O (g7882), .I (g7479));
INVX1 gate5995(.O (g3768), .I (I6979));
INVX1 gate5996(.O (g10896), .I (I16650));
INVX1 gate5997(.O (I13403), .I (g8236));
INVX1 gate5998(.O (g11344), .I (I17155));
INVX1 gate5999(.O (g4307), .I (g4013));
INVX1 gate6000(.O (g4536), .I (g3880));
INVX1 gate6001(.O (g10228), .I (I15604));
INVX1 gate6002(.O (g4159), .I (I7300));
INVX1 gate6003(.O (g2346), .I (I5414));
INVX1 gate6004(.O (g4359), .I (g3880));
INVX1 gate6005(.O (I12469), .I (g7531));
INVX1 gate6006(.O (g6735), .I (I10736));
INVX1 gate6007(.O (g8183), .I (I13102));
INVX1 gate6008(.O (g8608), .I (g8482));
INVX1 gate6009(.O (g8924), .I (I14249));
INVX1 gate6010(.O (g5830), .I (I9446));
INVX1 gate6011(.O (g7611), .I (I12183));
INVX1 gate6012(.O (g8220), .I (g7826));
INVX1 gate6013(.O (I12286), .I (g7231));
INVX1 gate6014(.O (I14561), .I (g9025));
INVX1 gate6015(.O (g5727), .I (I9273));
INVX1 gate6016(.O (g2103), .I (I4961));
INVX1 gate6017(.O (I8919), .I (g4576));
INVX1 gate6018(.O (g3943), .I (g2779));
INVX1 gate6019(.O (I9177), .I (g4904));
INVX1 gate6020(.O (I7233), .I (g2817));
INVX1 gate6021(.O (I10144), .I (g5689));
INVX1 gate6022(.O (g9340), .I (I14525));
INVX1 gate6023(.O (I14295), .I (g8806));
INVX1 gate6024(.O (I9377), .I (g5576));
INVX1 gate6025(.O (I17219), .I (g11292));
INVX1 gate6026(.O (g7799), .I (I12562));
INVX1 gate6027(.O (g4757), .I (I8109));
INVX1 gate6028(.O (I16604), .I (g10786));
INVX1 gate6029(.O (I7054), .I (g3093));
INVX1 gate6030(.O (I11572), .I (g6822));
INVX1 gate6031(.O (g8423), .I (I13583));
INVX1 gate6032(.O (g6475), .I (g5987));
INVX1 gate6033(.O (g4416), .I (g3638));
INVX1 gate6034(.O (g7981), .I (g7624));
INVX1 gate6035(.O (g6949), .I (I11091));
INVX1 gate6036(.O (g3228), .I (I6409));
INVX1 gate6037(.O (g8977), .I (I14352));
INVX1 gate6038(.O (g2732), .I (I5792));
INVX1 gate6039(.O (I9287), .I (g5576));
INVX1 gate6040(.O (g9082), .I (g8892));
INVX1 gate6041(.O (g10310), .I (I15736));
INVX1 gate6042(.O (g8588), .I (I13831));
INVX1 gate6043(.O (g7997), .I (g7697));
INVX1 gate6044(.O (g2753), .I (I5827));
INVX1 gate6045(.O (I12601), .I (g7629));
INVX1 gate6046(.O (g6292), .I (I10135));
INVX1 gate6047(.O (I11127), .I (g6452));
INVX1 gate6048(.O (g4315), .I (g3863));
INVX1 gate6049(.O (g4811), .I (g3661));
INVX1 gate6050(.O (g2508), .I (g940));
INVX1 gate6051(.O (g8361), .I (I13463));
INVX1 gate6052(.O (g10379), .I (I15861));
INVX1 gate6053(.O (I10966), .I (g6561));
INVX1 gate6054(.O (g2240), .I (g88));
INVX1 gate6055(.O (I8004), .I (g3967));
INVX1 gate6056(.O (g2072), .I (I4876));
INVX1 gate6057(.O (g3433), .I (I6648));
INVX1 gate6058(.O (I6921), .I (g2839));
INVX1 gate6059(.O (I5279), .I (g73));
INVX1 gate6060(.O (g7332), .I (I11644));
INVX1 gate6061(.O (g10050), .I (I15269));
INVX1 gate6062(.O (I9199), .I (g4935));
INVX1 gate6063(.O (g10378), .I (I15858));
INVX1 gate6064(.O (I8647), .I (g4219));
INVX1 gate6065(.O (I9399), .I (g5013));
INVX1 gate6066(.O (g5624), .I (I9056));
INVX1 gate6067(.O (g7680), .I (g7148));
INVX1 gate6068(.O (g11506), .I (I17537));
INVX1 gate6069(.O (g7353), .I (I11707));
INVX1 gate6070(.O (g2043), .I (g1801));
INVX1 gate6071(.O (g6084), .I (I9731));
INVX1 gate6072(.O (g8327), .I (g8164));
INVX1 gate6073(.O (I14364), .I (g8952));
INVX1 gate6074(.O (g4874), .I (I8215));
INVX1 gate6075(.O (g6039), .I (I9652));
INVX1 gate6076(.O (g5068), .I (g4840));
INVX1 gate6077(.O (I11956), .I (g6912));
INVX1 gate6078(.O (g3096), .I (g2482));
INVX1 gate6079(.O (I13956), .I (g8451));
INVX1 gate6080(.O (I13376), .I (g8226));
INVX1 gate6081(.O (I13385), .I (g8230));
INVX1 gate6082(.O (I11103), .I (g6667));
INVX1 gate6083(.O (g3496), .I (I6686));
INVX1 gate6084(.O (g7744), .I (I12397));
INVX1 gate6085(.O (I11889), .I (g6898));
INVX1 gate6086(.O (I17470), .I (g11452));
INVX1 gate6087(.O (g7802), .I (I12571));
INVX1 gate6088(.O (I5652), .I (g554));
INVX1 gate6089(.O (g8146), .I (g8033));
INVX1 gate6090(.O (I5057), .I (g1961));
INVX1 gate6091(.O (I11354), .I (g6553));
INVX1 gate6092(.O (g2116), .I (I5020));
INVX1 gate6093(.O (g8346), .I (I13418));
INVX1 gate6094(.O (I5843), .I (g2509));
INVX1 gate6095(.O (I13354), .I (g8214));
INVX1 gate6096(.O (I8503), .I (g4445));
INVX1 gate6097(.O (I5989), .I (g2252));
INVX1 gate6098(.O (I9510), .I (g5421));
INVX1 gate6099(.O (I11824), .I (g7246));
INVX1 gate6100(.O (g2034), .I (g1766));
INVX1 gate6101(.O (g5677), .I (I9188));
INVX1 gate6102(.O (g8103), .I (g7994));
INVX1 gate6103(.O (g3395), .I (I6601));
INVX1 gate6104(.O (g2434), .I (g1362));
INVX1 gate6105(.O (g3337), .I (g2745));
INVX1 gate6106(.O (g3913), .I (g2920));
INVX1 gate6107(.O (I10289), .I (g6003));
INVX1 gate6108(.O (I17277), .I (g11390));
INVX1 gate6109(.O (I12168), .I (g7256));
INVX1 gate6110(.O (I11671), .I (g7047));
INVX1 gate6111(.O (g9310), .I (I14503));
INVX1 gate6112(.O (g6583), .I (I10535));
INVX1 gate6113(.O (g6702), .I (g5949));
INVX1 gate6114(.O (g4880), .I (g3638));
INVX1 gate6115(.O (g5866), .I (g5361));
INVX1 gate6116(.O (g8696), .I (g8656));
INVX1 gate6117(.O (I5549), .I (g868));
INVX1 gate6118(.O (I7029), .I (g2946));
INVX1 gate6119(.O (I14309), .I (g8813));
INVX1 gate6120(.O (g2347), .I (g1945));
INVX1 gate6121(.O (I7429), .I (g3344));
INVX1 gate6122(.O (g10802), .I (I16510));
INVX1 gate6123(.O (g5149), .I (I8551));
INVX1 gate6124(.O (I9144), .I (g5007));
INVX1 gate6125(.O (I14224), .I (g8794));
INVX1 gate6126(.O (g6919), .I (g6453));
INVX1 gate6127(.O (I10308), .I (g6003));
INVX1 gate6128(.O (I12363), .I (g7187));
INVX1 gate6129(.O (I7956), .I (g3428));
INVX1 gate6130(.O (g7901), .I (g7712));
INVX1 gate6131(.O (g4272), .I (g3586));
INVX1 gate6132(.O (I8320), .I (g4452));
INVX1 gate6133(.O (g10730), .I (I16407));
INVX1 gate6134(.O (I12478), .I (g7560));
INVX1 gate6135(.O (I12015), .I (g6924));
INVX1 gate6136(.O (g6276), .I (I10087));
INVX1 gate6137(.O (g11649), .I (I17749));
INVX1 gate6138(.O (g9824), .I (I14973));
INVX1 gate6139(.O (g4243), .I (g3524));
INVX1 gate6140(.O (g3266), .I (I6436));
INVX1 gate6141(.O (I9259), .I (g5301));
INVX1 gate6142(.O (g8240), .I (g7972));
INVX1 gate6143(.O (g2914), .I (I6091));
INVX1 gate6144(.O (g5198), .I (I8614));
INVX1 gate6145(.O (g5747), .I (I9317));
INVX1 gate6146(.O (I15491), .I (g10093));
INVX1 gate6147(.O (g2210), .I (g103));
INVX1 gate6148(.O (g4417), .I (I7757));
INVX1 gate6149(.O (I10495), .I (g6144));
INVX1 gate6150(.O (g8472), .I (I13666));
INVX1 gate6151(.O (g6561), .I (g5773));
INVX1 gate6152(.O (g11648), .I (I17746));
INVX1 gate6153(.O (g4935), .I (g4420));
INVX1 gate6154(.O (g9762), .I (I14903));
INVX1 gate6155(.O (I17419), .I (g11421));
INVX1 gate6156(.O (I12556), .I (g7678));
INVX1 gate6157(.O (I15604), .I (g10148));
INVX1 gate6158(.O (I10816), .I (g6406));
INVX1 gate6159(.O (I9923), .I (g5308));
INVX1 gate6160(.O (g2013), .I (g1101));
INVX1 gate6161(.O (g8443), .I (I13627));
INVX1 gate6162(.O (g7600), .I (I12150));
INVX1 gate6163(.O (I12580), .I (g7540));
INVX1 gate6164(.O (g7574), .I (g6995));
INVX1 gate6165(.O (I6085), .I (g2234));
INVX1 gate6166(.O (g10548), .I (I16209));
INVX1 gate6167(.O (I17155), .I (g11310));
INVX1 gate6168(.O (g3142), .I (I6360));
INVX1 gate6169(.O (g5241), .I (g4386));
INVX1 gate6170(.O (g6527), .I (I10445));
INVX1 gate6171(.O (I12223), .I (g7049));
INVX1 gate6172(.O (g4328), .I (g4130));
INVX1 gate6173(.O (I14687), .I (g9258));
INVX1 gate6174(.O (I17170), .I (g11294));
INVX1 gate6175(.O (I14976), .I (g9670));
INVX1 gate6176(.O (g8116), .I (I12971));
INVX1 gate6177(.O (g3255), .I (I6421));
INVX1 gate6178(.O (I7639), .I (g3722));
INVX1 gate6179(.O (g8316), .I (I13332));
INVX1 gate6180(.O (g3815), .I (g3228));
INVX1 gate6181(.O (I11211), .I (g6527));
INVX1 gate6182(.O (I10374), .I (g5852));
INVX1 gate6183(.O (g6764), .I (g5987));
INVX1 gate6184(.O (I7109), .I (g2970));
INVX1 gate6185(.O (I5909), .I (g2207));
INVX1 gate6186(.O (I16534), .I (g10747));
INVX1 gate6187(.O (I10643), .I (g6026));
INVX1 gate6188(.O (I11088), .I (g6434));
INVX1 gate6189(.O (I11024), .I (g6399));
INVX1 gate6190(.O (g9556), .I (I14701));
INVX1 gate6191(.O (I16098), .I (g10369));
INVX1 gate6192(.O (g10317), .I (I15749));
INVX1 gate6193(.O (g8565), .I (I13788));
INVX1 gate6194(.O (g2820), .I (I5926));
INVX1 gate6195(.O (g3097), .I (g2482));
INVX1 gate6196(.O (I9886), .I (g5286));
INVX1 gate6197(.O (I6941), .I (g2858));
INVX1 gate6198(.O (g3726), .I (I6898));
INVX1 gate6199(.O (g7580), .I (I12056));
INVX1 gate6200(.O (g6503), .I (I10421));
INVX1 gate6201(.O (g5644), .I (I9093));
INVX1 gate6202(.O (I5740), .I (g2341));
INVX1 gate6203(.O (g6970), .I (I11122));
INVX1 gate6204(.O (g8347), .I (I13421));
INVX1 gate6205(.O (I15395), .I (g10058));
INVX1 gate6206(.O (g2317), .I (g622));
INVX1 gate6207(.O (I8892), .I (g4554));
INVX1 gate6208(.O (g10129), .I (I15389));
INVX1 gate6209(.O (g9930), .I (I15127));
INVX1 gate6210(.O (I9114), .I (g5603));
INVX1 gate6211(.O (g6925), .I (I11043));
INVX1 gate6212(.O (I17194), .I (g11317));
INVX1 gate6213(.O (I7707), .I (g3370));
INVX1 gate6214(.O (g11395), .I (I17228));
INVX1 gate6215(.O (g1962), .I (g27));
INVX1 gate6216(.O (g10057), .I (I15278));
INVX1 gate6217(.O (g2601), .I (I5704));
INVX1 gate6218(.O (g10128), .I (I15386));
INVX1 gate6219(.O (g5818), .I (g5320));
INVX1 gate6220(.O (g8697), .I (g8660));
INVX1 gate6221(.O (I6520), .I (g3186));
INVX1 gate6222(.O (I14668), .I (g9309));
INVX1 gate6223(.O (g4213), .I (I7456));
INVX1 gate6224(.O (g11633), .I (I17713));
INVX1 gate6225(.O (I11659), .I (g7097));
INVX1 gate6226(.O (I12186), .I (g7264));
INVX1 gate6227(.O (g6120), .I (I9813));
INVX1 gate6228(.O (I10195), .I (g6116));
INVX1 gate6229(.O (I6031), .I (g2209));
INVX1 gate6230(.O (I12953), .I (g8024));
INVX1 gate6231(.O (g10323), .I (I15763));
INVX1 gate6232(.O (g11191), .I (g11112));
INVX1 gate6233(.O (g2775), .I (I5862));
INVX1 gate6234(.O (g7076), .I (I11303));
INVX1 gate6235(.O (I6812), .I (g3290));
INVX1 gate6236(.O (g3783), .I (I7009));
INVX1 gate6237(.O (g7476), .I (g6933));
INVX1 gate6238(.O (I6958), .I (g2872));
INVX1 gate6239(.O (g5893), .I (g5106));
INVX1 gate6240(.O (g6277), .I (I10090));
INVX1 gate6241(.O (I14525), .I (g9109));
INVX1 gate6242(.O (I14424), .I (g8945));
INVX1 gate6243(.O (g3112), .I (g2482));
INVX1 gate6244(.O (g3267), .I (I6439));
INVX1 gate6245(.O (g10775), .I (I16461));
INVX1 gate6246(.O (I16766), .I (g10892));
INVX1 gate6247(.O (I12936), .I (g7983));
INVX1 gate6248(.O (I15832), .I (g10206));
INVX1 gate6249(.O (I8340), .I (g4804));
INVX1 gate6250(.O (I11296), .I (g6525));
INVX1 gate6251(.O (g2060), .I (g1380));
INVX1 gate6252(.O (g6617), .I (g6019));
INVX1 gate6253(.O (I14558), .I (g9024));
INVX1 gate6254(.O (g6789), .I (I10789));
INVX1 gate6255(.O (I17749), .I (g11644));
INVX1 gate6256(.O (I11644), .I (g6970));
INVX1 gate6257(.O (I17616), .I (g11561));
INVX1 gate6258(.O (I16871), .I (g10973));
INVX1 gate6259(.O (I11338), .I (g6680));
INVX1 gate6260(.O (I13338), .I (g8210));
INVX1 gate6261(.O (I9594), .I (g5083));
INVX1 gate6262(.O (g4166), .I (I7315));
INVX1 gate6263(.O (g11440), .I (I17371));
INVX1 gate6264(.O (g4366), .I (I7659));
INVX1 gate6265(.O (g5426), .I (I8869));
INVX1 gate6266(.O (I15861), .I (g10339));
INVX1 gate6267(.O (I16360), .I (g10590));
INVX1 gate6268(.O (I6911), .I (g2825));
INVX1 gate6269(.O (I13969), .I (g8451));
INVX1 gate6270(.O (I7833), .I (g3585));
INVX1 gate6271(.O (g7285), .I (I11531));
INVX1 gate6272(.O (g3329), .I (I6504));
INVX1 gate6273(.O (I15247), .I (g10032));
INVX1 gate6274(.O (g11573), .I (g11561));
INVX1 gate6275(.O (I5525), .I (g589));
INVX1 gate6276(.O (I5710), .I (g2431));
INVX1 gate6277(.O (g3761), .I (I6962));
INVX1 gate6278(.O (g5614), .I (I9040));
INVX1 gate6279(.O (I12762), .I (g7541));
INVX1 gate6280(.O (I17704), .I (g11618));
INVX1 gate6281(.O (g4056), .I (I7173));
INVX1 gate6282(.O (g7500), .I (g6943));
INVX1 gate6283(.O (I10713), .I (g6003));
INVX1 gate6284(.O (g8317), .I (I13335));
INVX1 gate6285(.O (I15389), .I (g10110));
INVX1 gate6286(.O (g4456), .I (g3375));
INVX1 gate6287(.O (I14713), .I (g9052));
INVX1 gate6288(.O (g6299), .I (I10156));
INVX1 gate6289(.O (g5821), .I (I9433));
INVX1 gate6290(.O (g3828), .I (g2920));
INVX1 gate6291(.O (g10697), .I (I16370));
INVX1 gate6292(.O (g6547), .I (g5893));
INVX1 gate6293(.O (I13197), .I (g8186));
INVX1 gate6294(.O (g11389), .I (I17216));
INVX1 gate6295(.O (g11045), .I (I16796));
INVX1 gate6296(.O (I6733), .I (g3321));
INVX1 gate6297(.O (I9065), .I (g4760));
INVX1 gate6298(.O (I17466), .I (g11447));
INVX1 gate6299(.O (g8601), .I (g8477));
INVX1 gate6300(.O (g10261), .I (g10126));
INVX1 gate6301(.O (g2937), .I (I6106));
INVX1 gate6302(.O (g3727), .I (I6901));
INVX1 gate6303(.O (g2079), .I (I4891));
INVX1 gate6304(.O (g5984), .I (I9602));
INVX1 gate6305(.O (I10610), .I (g5879));
INVX1 gate6306(.O (g10880), .I (I16610));
INVX1 gate6307(.O (I15701), .I (g10236));
INVX1 gate6308(.O (g4355), .I (I7642));
INVX1 gate6309(.O (g11388), .I (I17213));
INVX1 gate6310(.O (g7339), .I (I11665));
INVX1 gate6311(.O (g2479), .I (g26));
INVX1 gate6312(.O (I10042), .I (g5723));
INVX1 gate6313(.O (I15272), .I (g10019));
INVX1 gate6314(.O (I16629), .I (g10860));
INVX1 gate6315(.O (g2840), .I (I5960));
INVX1 gate6316(.O (I10189), .I (g6112));
INVX1 gate6317(.O (g7024), .I (I11169));
INVX1 gate6318(.O (I16220), .I (g10502));
INVX1 gate6319(.O (g2190), .I (I5149));
INVX1 gate6320(.O (g4260), .I (I7513));
INVX1 gate6321(.O (g2390), .I (I5475));
INVX1 gate6322(.O (g7795), .I (I12550));
INVX1 gate6323(.O (I9433), .I (g5069));
INVX1 gate6324(.O (I17642), .I (g11579));
INVX1 gate6325(.O (I10678), .I (g5777));
INVX1 gate6326(.O (g7737), .I (I12388));
INVX1 gate6327(.O (g7809), .I (I12592));
INVX1 gate6328(.O (g3703), .I (g2920));
INVX1 gate6329(.O (I14188), .I (g8792));
INVX1 gate6330(.O (I14678), .I (g9265));
INVX1 gate6331(.O (g5106), .I (I8490));
INVX1 gate6332(.O (g4463), .I (g3829));
INVX1 gate6333(.O (I9096), .I (g5568));
INVX1 gate6334(.O (g2156), .I (I5073));
INVX1 gate6335(.O (g7672), .I (I12293));
INVX1 gate6336(.O (I14939), .I (g9454));
INVX1 gate6337(.O (g2356), .I (I5438));
INVX1 gate6338(.O (g7077), .I (I11306));
INVX1 gate6339(.O (g6709), .I (g5949));
INVX1 gate6340(.O (I17733), .I (g11639));
INVX1 gate6341(.O (g9814), .I (g9490));
INVX1 gate6342(.O (g5790), .I (I9388));
INVX1 gate6343(.O (I9550), .I (g5030));
INVX1 gate6344(.O (I10030), .I (g5685));
INVX1 gate6345(.O (g7477), .I (I11869));
INVX1 gate6346(.O (I10093), .I (g5779));
INVX1 gate6347(.O (I9845), .I (g5405));
INVX1 gate6348(.O (g3624), .I (I6767));
INVX1 gate6349(.O (g6140), .I (I9851));
INVX1 gate6350(.O (g6340), .I (I10243));
INVX1 gate6351(.O (I5111), .I (g39));
INVX1 gate6352(.O (I11581), .I (g6826));
INVX1 gate6353(.O (I11450), .I (g6488));
INVX1 gate6354(.O (I12568), .I (g7502));
INVX1 gate6355(.O (g9350), .I (I14555));
INVX1 gate6356(.O (g10499), .I (I16124));
INVX1 gate6357(.O (I5311), .I (g98));
INVX1 gate6358(.O (g3068), .I (g2303));
INVX1 gate6359(.O (I13714), .I (g8351));
INVX1 gate6360(.O (I11315), .I (g6644));
INVX1 gate6361(.O (g8784), .I (I14087));
INVX1 gate6362(.O (g2942), .I (I6121));
INVX1 gate6363(.O (g8739), .I (g8640));
INVX1 gate6364(.O (I12242), .I (g7089));
INVX1 gate6365(.O (g4279), .I (I7536));
INVX1 gate6366(.O (I11707), .I (g7009));
INVX1 gate6367(.O (g7205), .I (I11433));
INVX1 gate6368(.O (g9773), .I (g9474));
INVX1 gate6369(.O (I7086), .I (g3142));
INVX1 gate6370(.O (I13819), .I (g8488));
INVX1 gate6371(.O (g11061), .I (g10974));
INVX1 gate6372(.O (g10498), .I (I16121));
INVX1 gate6373(.O (g9009), .I (I14405));
INVX1 gate6374(.O (g6435), .I (I10355));
INVX1 gate6375(.O (g4167), .I (I7318));
INVX1 gate6376(.O (g5027), .I (I8396));
INVX1 gate6377(.O (g6517), .I (I10434));
INVX1 gate6378(.O (g6082), .I (I9727));
INVX1 gate6379(.O (I12123), .I (g6861));
INVX1 gate6380(.O (g4318), .I (g4130));
INVX1 gate6381(.O (g4367), .I (I7662));
INVX1 gate6382(.O (I16859), .I (g10911));
INVX1 gate6383(.O (g4872), .I (I8211));
INVX1 gate6384(.O (g7634), .I (I12242));
INVX1 gate6385(.O (I5174), .I (g52));
INVX1 gate6386(.O (I16950), .I (g11081));
INVX1 gate6387(.O (g8079), .I (I12939));
INVX1 gate6388(.O (I16370), .I (g10592));
INVX1 gate6389(.O (g6482), .I (I10412));
INVX1 gate6390(.O (I11055), .I (g6419));
INVX1 gate6391(.O (g10056), .I (I15275));
INVX1 gate6392(.O (I9807), .I (g5419));
INVX1 gate6393(.O (g8479), .I (g8319));
INVX1 gate6394(.O (I7185), .I (g2626));
INVX1 gate6395(.O (I12751), .I (g7626));
INVX1 gate6396(.O (g9769), .I (I14918));
INVX1 gate6397(.O (g4057), .I (I7176));
INVX1 gate6398(.O (g5904), .I (I9539));
INVX1 gate6399(.O (g7304), .I (I11560));
INVX1 gate6400(.O (g5200), .I (g4567));
INVX1 gate6401(.O (g10080), .I (I15308));
INVX1 gate6402(.O (g8294), .I (I13236));
INVX1 gate6403(.O (I13978), .I (g8575));
INVX1 gate6404(.O (g4457), .I (g3829));
INVX1 gate6405(.O (g2163), .I (I5092));
INVX1 gate6406(.O (I8877), .I (g4421));
INVX1 gate6407(.O (g2363), .I (I5441));
INVX1 gate6408(.O (I7070), .I (g3138));
INVX1 gate6409(.O (g5446), .I (I8877));
INVX1 gate6410(.O (I11590), .I (g6829));
INVX1 gate6411(.O (I16172), .I (g10498));
INVX1 gate6412(.O (g4193), .I (I7396));
INVX1 gate6413(.O (g3716), .I (I6876));
INVX1 gate6414(.O (g11360), .I (I17185));
INVX1 gate6415(.O (g4393), .I (I7726));
INVX1 gate6416(.O (I10837), .I (g6717));
INVX1 gate6417(.O (g2432), .I (I5513));
INVX1 gate6418(.O (I12293), .I (g7116));
INVX1 gate6419(.O (g10271), .I (I15665));
INVX1 gate6420(.O (I12638), .I (g7708));
INVX1 gate6421(.O (g11447), .I (I17390));
INVX1 gate6422(.O (I13741), .I (g8296));
INVX1 gate6423(.O (I15162), .I (g9958));
INVX1 gate6424(.O (g4549), .I (I7956));
INVX1 gate6425(.O (I17555), .I (g11503));
INVX1 gate6426(.O (I6898), .I (g2964));
INVX1 gate6427(.O (I12265), .I (g7211));
INVX1 gate6428(.O (g11162), .I (g10950));
INVX1 gate6429(.O (g7754), .I (I12427));
INVX1 gate6430(.O (g10461), .I (I15974));
INVX1 gate6431(.O (g5191), .I (g4640));
INVX1 gate6432(.O (g8156), .I (I13051));
INVX1 gate6433(.O (I9248), .I (g4954));
INVX1 gate6434(.O (g3747), .I (g3015));
INVX1 gate6435(.O (I11094), .I (g6657));
INVX1 gate6436(.O (g1973), .I (g466));
INVX1 gate6437(.O (g5391), .I (I8827));
INVX1 gate6438(.O (g8356), .I (I13448));
INVX1 gate6439(.O (g10342), .I (I15792));
INVX1 gate6440(.O (g3398), .I (g2896));
INVX1 gate6441(.O (g6214), .I (g5446));
INVX1 gate6442(.O (g7273), .I (g6365));
INVX1 gate6443(.O (I5020), .I (g1176));
INVX1 gate6444(.O (I6510), .I (g3267));
INVX1 gate6445(.O (g9993), .I (I15193));
INVX1 gate6446(.O (g10145), .I (I15437));
INVX1 gate6447(.O (g10031), .I (I15229));
INVX1 gate6448(.O (g6110), .I (I9783));
INVX1 gate6449(.O (g5637), .I (I9074));
INVX1 gate6450(.O (g6310), .I (I10189));
INVX1 gate6451(.O (g11629), .I (I17701));
INVX1 gate6452(.O (g9822), .I (I14967));
INVX1 gate6453(.O (g10199), .I (g10172));
INVX1 gate6454(.O (g11451), .I (I17410));
INVX1 gate6455(.O (g11472), .I (I17453));
INVX1 gate6456(.O (g7044), .I (I11217));
INVX1 gate6457(.O (g10887), .I (I16623));
INVX1 gate6458(.O (g2912), .I (I6085));
INVX1 gate6459(.O (I13735), .I (g8293));
INVX1 gate6460(.O (g1969), .I (g456));
INVX1 gate6461(.O (g4121), .I (I7264));
INVX1 gate6462(.O (g5107), .I (g4459));
INVX1 gate6463(.O (g8704), .I (g8667));
INVX1 gate6464(.O (g4321), .I (g3863));
INVX1 gate6465(.O (g2157), .I (g1703));
INVX1 gate6466(.O (g11628), .I (I17698));
INVX1 gate6467(.O (g10198), .I (I15568));
INVX1 gate6468(.O (I7131), .I (g2640));
INVX1 gate6469(.O (I7006), .I (g2912));
INVX1 gate6470(.O (g7983), .I (I12793));
INVX1 gate6471(.O (I10201), .I (g5998));
INVX1 gate6472(.O (g5223), .I (g4640));
INVX1 gate6473(.O (I11695), .I (g7052));
INVX1 gate6474(.O (g10528), .I (g10464));
INVX1 gate6475(.O (g10696), .I (g10621));
INVX1 gate6476(.O (g4232), .I (I7487));
INVX1 gate6477(.O (I12835), .I (g7660));
INVX1 gate6478(.O (I13695), .I (g8363));
INVX1 gate6479(.O (g10330), .I (I15778));
INVX1 gate6480(.O (g5858), .I (I9475));
INVX1 gate6481(.O (g10393), .I (g10317));
INVX1 gate6482(.O (I10075), .I (g5724));
INVX1 gate6483(.O (I7766), .I (g3770));
INVX1 gate6484(.O (g8954), .I (I14315));
INVX1 gate6485(.O (I16540), .I (g10722));
INVX1 gate6486(.O (g6236), .I (I9981));
INVX1 gate6487(.O (I6694), .I (g2749));
INVX1 gate6488(.O (g7543), .I (I11961));
INVX1 gate6489(.O (I12586), .I (g7561));
INVX1 gate6490(.O (g11071), .I (g10913));
INVX1 gate6491(.O (g8363), .I (I13469));
INVX1 gate6492(.O (I7487), .I (g3371));
INVX1 gate6493(.O (I8237), .I (g4295));
INVX1 gate6494(.O (g5416), .I (I8851));
INVX1 gate6495(.O (I14494), .I (g8887));
INVX1 gate6496(.O (g3119), .I (I6347));
INVX1 gate6497(.O (g10132), .I (g10063));
INVX1 gate6498(.O (I17519), .I (g11484));
INVX1 gate6499(.O (g10869), .I (I16577));
INVX1 gate6500(.O (I6088), .I (g2235));
INVX1 gate6501(.O (I17176), .I (g11286));
INVX1 gate6502(.O (I17185), .I (g11311));
INVX1 gate6503(.O (I10623), .I (g6002));
INVX1 gate6504(.O (I12442), .I (g7672));
INVX1 gate6505(.O (I17675), .I (g11606));
INVX1 gate6506(.O (I17092), .I (g11217));
INVX1 gate6507(.O (I16203), .I (g10454));
INVX1 gate6508(.O (g4519), .I (I7920));
INVX1 gate6509(.O (g5251), .I (g4640));
INVX1 gate6510(.O (g6590), .I (g5949));
INVX1 gate6511(.O (g6877), .I (I10963));
INVX1 gate6512(.O (I4777), .I (g18));
INVX1 gate6513(.O (g10868), .I (I16574));
INVX1 gate6514(.O (g5811), .I (I9415));
INVX1 gate6515(.O (g5642), .I (I9087));
INVX1 gate6516(.O (g3352), .I (I6538));
INVX1 gate6517(.O (I9783), .I (g5395));
INVX1 gate6518(.O (g2626), .I (g2000));
INVX1 gate6519(.O (g7534), .I (I11942));
INVX1 gate6520(.O (g7729), .I (I12372));
INVX1 gate6521(.O (g7961), .I (g7664));
INVX1 gate6522(.O (g5047), .I (g4354));
INVX1 gate6523(.O (I13457), .I (g8184));
INVX1 gate6524(.O (I10984), .I (g6757));
INVX1 gate6525(.O (g9895), .I (I15088));
INVX1 gate6526(.O (g6657), .I (I10620));
INVX1 gate6527(.O (g10161), .I (I15479));
INVX1 gate6528(.O (g4552), .I (g3880));
INVX1 gate6529(.O (g4606), .I (g3829));
INVX1 gate6530(.O (I15858), .I (g10336));
INVX1 gate6531(.O (g8568), .I (I13797));
INVX1 gate6532(.O (I8089), .I (g3545));
INVX1 gate6533(.O (I10352), .I (g6216));
INVX1 gate6534(.O (g6556), .I (g5747));
INVX1 gate6535(.O (I14352), .I (g8946));
INVX1 gate6536(.O (g7927), .I (g7500));
INVX1 gate6537(.O (I10822), .I (g6584));
INVX1 gate6538(.O (g5874), .I (I9491));
INVX1 gate6539(.O (I9001), .I (g4762));
INVX1 gate6540(.O (g10259), .I (g10141));
INVX1 gate6541(.O (I14418), .I (g8941));
INVX1 gate6542(.O (g10708), .I (I16387));
INVX1 gate6543(.O (I16739), .I (g10856));
INVX1 gate6544(.O (I12430), .I (g7649));
INVX1 gate6545(.O (g3186), .I (I6373));
INVX1 gate6546(.O (g5654), .I (I9123));
INVX1 gate6547(.O (I12493), .I (g7650));
INVX1 gate6548(.O (g10471), .I (g10378));
INVX1 gate6549(.O (g7414), .I (I11794));
INVX1 gate6550(.O (I9293), .I (g5486));
INVX1 gate6551(.O (g3386), .I (g3144));
INVX1 gate6552(.O (g10087), .I (I15314));
INVX1 gate6553(.O (g8357), .I (I13451));
INVX1 gate6554(.O (I9129), .I (g4892));
INVX1 gate6555(.O (g7946), .I (g7416));
INVX1 gate6556(.O (g10258), .I (g10198));
INVX1 gate6557(.O (g3975), .I (g3121));
INVX1 gate6558(.O (I7173), .I (g2644));
INVX1 gate6559(.O (I9329), .I (g5504));
INVX1 gate6560(.O (I5973), .I (g2247));
INVX1 gate6561(.O (g4586), .I (g4089));
INVX1 gate6562(.O (g11394), .I (I17225));
INVX1 gate6563(.O (g6464), .I (I10398));
INVX1 gate6564(.O (g7903), .I (g7446));
INVX1 gate6565(.O (g2683), .I (g2037));
INVX1 gate6566(.O (I11689), .I (g7044));
INVX1 gate6567(.O (I6870), .I (g2852));
INVX1 gate6568(.O (g3274), .I (I6454));
INVX1 gate6569(.O (g3426), .I (g3121));
INVX1 gate6570(.O (g5880), .I (g5361));
INVX1 gate6571(.O (I12035), .I (g6930));
INVX1 gate6572(.O (I13280), .I (g8250));
INVX1 gate6573(.O (g2778), .I (g2276));
INVX1 gate6574(.O (g10244), .I (g10131));
INVX1 gate6575(.O (I9727), .I (g5250));
INVX1 gate6576(.O (I7369), .I (g4051));
INVX1 gate6577(.O (g3370), .I (I6560));
INVX1 gate6578(.O (I10589), .I (g5763));
INVX1 gate6579(.O (I13624), .I (g8320));
INVX1 gate6580(.O (I14194), .I (g8798));
INVX1 gate6581(.O (g11420), .I (I17315));
INVX1 gate6582(.O (g6563), .I (g5783));
INVX1 gate6583(.O (I7920), .I (g3440));
INVX1 gate6584(.O (g5272), .I (I8724));
INVX1 gate6585(.O (g11319), .I (I17116));
INVX1 gate6586(.O (g7036), .I (g6420));
INVX1 gate6587(.O (g9085), .I (g8892));
INVX1 gate6588(.O (g10069), .I (I15296));
INVX1 gate6589(.O (I7459), .I (g3720));
INVX1 gate6590(.O (I9221), .I (g5236));
INVX1 gate6591(.O (g4525), .I (g3880));
INVX1 gate6592(.O (g7436), .I (g7227));
INVX1 gate6593(.O (g8626), .I (g8498));
INVX1 gate6594(.O (g6295), .I (I10144));
INVX1 gate6595(.O (I12517), .I (g7737));
INVX1 gate6596(.O (I13102), .I (g7928));
INVX1 gate6597(.O (g6237), .I (I9984));
INVX1 gate6598(.O (g11446), .I (I17387));
INVX1 gate6599(.O (g10774), .I (I16458));
INVX1 gate6600(.O (I17438), .I (g11444));
INVX1 gate6601(.O (I10477), .I (g6049));
INVX1 gate6602(.O (I16366), .I (g10591));
INVX1 gate6603(.O (g5417), .I (I8854));
INVX1 gate6604(.O (g2075), .I (I4883));
INVX1 gate6605(.O (I14477), .I (g8943));
INVX1 gate6606(.O (g10879), .I (I16607));
INVX1 gate6607(.O (I16632), .I (g10861));
INVX1 gate6608(.O (g11059), .I (g10974));
INVX1 gate6609(.O (g6844), .I (I10904));
INVX1 gate6610(.O (g7335), .I (I11653));
INVX1 gate6611(.O (g2475), .I (g192));
INVX1 gate6612(.O (I14119), .I (g8779));
INVX1 gate6613(.O (g1988), .I (g766));
INVX1 gate6614(.O (g3544), .I (g3164));
INVX1 gate6615(.O (g2949), .I (I6150));
INVX1 gate6616(.O (g7288), .I (I11540));
INVX1 gate6617(.O (g11540), .I (g11519));
INVX1 gate6618(.O (g5982), .I (I9598));
INVX1 gate6619(.O (g10878), .I (I16604));
INVX1 gate6620(.O (I7793), .I (g3783));
INVX1 gate6621(.O (I10864), .I (g6634));
INVX1 gate6622(.O (g3636), .I (I6815));
INVX1 gate6623(.O (g5629), .I (I9065));
INVX1 gate6624(.O (I9953), .I (g5484));
INVX1 gate6625(.O (g6089), .I (g4977));
INVX1 gate6626(.O (I12193), .I (g7270));
INVX1 gate6627(.O (g10171), .I (I15507));
INVX1 gate6628(.O (g6731), .I (g6001));
INVX1 gate6629(.O (I9068), .I (g4768));
INVX1 gate6630(.O (g7805), .I (I12580));
INVX1 gate6631(.O (I5655), .I (g557));
INVX1 gate6632(.O (g7916), .I (g7651));
INVX1 gate6633(.O (g11203), .I (g11112));
INVX1 gate6634(.O (g5542), .I (I8967));
INVX1 gate6635(.O (g7022), .I (g6389));
INVX1 gate6636(.O (g3306), .I (I6477));
INVX1 gate6637(.O (g2998), .I (g2462));
INVX1 gate6638(.O (g2646), .I (g1992));
INVX1 gate6639(.O (g4158), .I (g3304));
INVX1 gate6640(.O (g7422), .I (I11810));
INVX1 gate6641(.O (g7749), .I (I12412));
INVX1 gate6642(.O (I6065), .I (g2226));
INVX1 gate6643(.O (g6557), .I (g5748));
INVX1 gate6644(.O (I12165), .I (g6882));
INVX1 gate6645(.O (I12523), .I (g7421));
INVX1 gate6646(.O (g10792), .I (I16492));
INVX1 gate6647(.O (g11044), .I (I16793));
INVX1 gate6648(.O (g3790), .I (g3228));
INVX1 gate6649(.O (I15281), .I (g10025));
INVX1 gate6650(.O (g2084), .I (I4900));
INVX1 gate6651(.O (g2603), .I (I5710));
INVX1 gate6652(.O (I8967), .I (g4482));
INVX1 gate6653(.O (g6705), .I (I10682));
INVX1 gate6654(.O (g2039), .I (g1781));
INVX1 gate6655(.O (I9677), .I (g5190));
INVX1 gate6656(.O (g3387), .I (I6587));
INVX1 gate6657(.O (I10305), .I (g6180));
INVX1 gate6658(.O (g5800), .I (I9402));
INVX1 gate6659(.O (I5410), .I (g901));
INVX1 gate6660(.O (g3461), .I (I6671));
INVX1 gate6661(.O (I15377), .I (g10104));
INVX1 gate6662(.O (g6242), .I (I9995));
INVX1 gate6663(.O (g2850), .I (I5976));
INVX1 gate6664(.O (g9431), .I (g9085));
INVX1 gate6665(.O (g7798), .I (I12559));
INVX1 gate6666(.O (g11301), .I (I17084));
INVX1 gate6667(.O (g10459), .I (I15968));
INVX1 gate6668(.O (g9812), .I (g9490));
INVX1 gate6669(.O (g3756), .I (g3015));
INVX1 gate6670(.O (g4587), .I (g3829));
INVX1 gate6671(.O (I12475), .I (g7545));
INVX1 gate6672(.O (g11377), .I (I17202));
INVX1 gate6673(.O (I9866), .I (g5274));
INVX1 gate6674(.O (g6948), .I (I11088));
INVX1 gate6675(.O (g3622), .I (I6757));
INVX1 gate6676(.O (g9958), .I (I15157));
INVX1 gate6677(.O (g7560), .I (I12012));
INVX1 gate6678(.O (g4275), .I (g3664));
INVX1 gate6679(.O (g4311), .I (g4130));
INVX1 gate6680(.O (g10458), .I (I15965));
INVX1 gate6681(.O (g8782), .I (I14083));
INVX1 gate6682(.O (g3427), .I (g3144));
INVX1 gate6683(.O (I15562), .I (g10098));
INVX1 gate6684(.O (I9349), .I (g5515));
INVX1 gate6685(.O (g6955), .I (I11103));
INVX1 gate6686(.O (I10036), .I (g5701));
INVX1 gate6687(.O (g4615), .I (I8024));
INVX1 gate6688(.O (g5213), .I (g4640));
INVX1 gate6689(.O (g11645), .I (I17739));
INVX1 gate6690(.O (I10177), .I (g6103));
INVX1 gate6691(.O (I10560), .I (g5887));
INVX1 gate6692(.O (I11456), .I (g6440));
INVX1 gate6693(.O (I14101), .I (g8774));
INVX1 gate6694(.O (I9848), .I (g5557));
INVX1 gate6695(.O (I15290), .I (g9984));
INVX1 gate6696(.O (g6254), .I (I10021));
INVX1 gate6697(.O (g8475), .I (g8314));
INVX1 gate6698(.O (g4174), .I (I7339));
INVX1 gate6699(.O (g6814), .I (I10852));
INVX1 gate6700(.O (g9765), .I (I14910));
INVX1 gate6701(.O (I17636), .I (g11577));
INVX1 gate6702(.O (I15698), .I (g10235));
INVX1 gate6703(.O (g10545), .I (I16200));
INVX1 gate6704(.O (g2919), .I (I6102));
INVX1 gate6705(.O (g7037), .I (I11198));
INVX1 gate6706(.O (g10079), .I (I15305));
INVX1 gate6707(.O (g10444), .I (g10325));
INVX1 gate6708(.O (I9699), .I (g5426));
INVX1 gate6709(.O (g6150), .I (I9869));
INVX1 gate6710(.O (I14642), .I (g9088));
INVX1 gate6711(.O (g7437), .I (I11829));
INVX1 gate6712(.O (I16784), .I (g10895));
INVX1 gate6713(.O (I5667), .I (g566));
INVX1 gate6714(.O (I6395), .I (g2334));
INVX1 gate6715(.O (I6891), .I (g2962));
INVX1 gate6716(.O (g8292), .I (I13230));
INVX1 gate6717(.O (g2952), .I (g2455));
INVX1 gate6718(.O (I16956), .I (g11096));
INVX1 gate6719(.O (g3345), .I (I6531));
INVX1 gate6720(.O (I16376), .I (g10596));
INVX1 gate6721(.O (I13314), .I (g8260));
INVX1 gate6722(.O (g4284), .I (g3664));
INVX1 gate6723(.O (g7579), .I (I12053));
INVX1 gate6724(.O (g8526), .I (I13735));
INVX1 gate6725(.O (g10598), .I (I16273));
INVX1 gate6726(.O (g3763), .I (I6968));
INVX1 gate6727(.O (I10733), .I (g6099));
INVX1 gate6728(.O (g4545), .I (I7952));
INVX1 gate6729(.O (I11076), .I (g6649));
INVX1 gate6730(.O (I11085), .I (g6433));
INVX1 gate6731(.O (g3391), .I (g2896));
INVX1 gate6732(.O (g9733), .I (I14876));
INVX1 gate6733(.O (I15427), .I (g10088));
INVX1 gate6734(.O (I16095), .I (g10401));
INVX1 gate6735(.O (g4180), .I (I7357));
INVX1 gate6736(.O (g5490), .I (I8911));
INVX1 gate6737(.O (g9270), .I (I14485));
INVX1 gate6738(.O (g4380), .I (I7701));
INVX1 gate6739(.O (g11427), .I (I17334));
INVX1 gate6740(.O (g5166), .I (g4682));
INVX1 gate6741(.O (I11596), .I (g6831));
INVX1 gate6742(.O (g4591), .I (g3829));
INVX1 gate6743(.O (I15632), .I (g10184));
INVX1 gate6744(.O (g11366), .I (I17191));
INVX1 gate6745(.O (g3637), .I (I6818));
INVX1 gate6746(.O (I7216), .I (g2952));
INVX1 gate6747(.O (g7752), .I (I12421));
INVX1 gate6748(.O (g11632), .I (I17710));
INVX1 gate6749(.O (g8484), .I (g8336));
INVX1 gate6750(.O (I16181), .I (g10491));
INVX1 gate6751(.O (I10630), .I (g5889));
INVX1 gate6752(.O (g8439), .I (I13615));
INVX1 gate6753(.O (g2004), .I (I4820));
INVX1 gate6754(.O (I10693), .I (g6068));
INVX1 gate6755(.O (g6836), .I (I10888));
INVX1 gate6756(.O (I12372), .I (g7137));
INVX1 gate6757(.O (g7917), .I (g7497));
INVX1 gate6758(.O (g2986), .I (I6220));
INVX1 gate6759(.O (g3307), .I (I6480));
INVX1 gate6760(.O (g9473), .I (g9103));
INVX1 gate6761(.O (I7671), .I (g3351));
INVX1 gate6762(.O (g2647), .I (g1993));
INVX1 gate6763(.O (g10159), .I (I15473));
INVX1 gate6764(.O (g4420), .I (I7766));
INVX1 gate6765(.O (g10125), .I (I15377));
INVX1 gate6766(.O (g10532), .I (g10473));
INVX1 gate6767(.O (g10901), .I (g10802));
INVX1 gate6768(.O (I10009), .I (g5542));
INVX1 gate6769(.O (g5649), .I (I9108));
INVX1 gate6770(.O (g3359), .I (I6543));
INVX1 gate6771(.O (I15403), .I (g10069));
INVX1 gate6772(.O (g1965), .I (g119));
INVX1 gate6773(.O (g4507), .I (g3546));
INVX1 gate6774(.O (g5348), .I (I8815));
INVX1 gate6775(.O (g6967), .I (I11119));
INVX1 gate6776(.O (I5555), .I (g110));
INVX1 gate6777(.O (I11269), .I (g6545));
INVX1 gate6778(.O (g9980), .I (I15181));
INVX1 gate6779(.O (g2764), .I (I5850));
INVX1 gate6780(.O (I8462), .I (g4475));
INVX1 gate6781(.O (g11403), .I (I17252));
INVX1 gate6782(.O (g10158), .I (I15470));
INVX1 gate6783(.O (g11547), .I (g11519));
INVX1 gate6784(.O (g7042), .I (I11211));
INVX1 gate6785(.O (I11773), .I (g7257));
INVX1 gate6786(.O (g10783), .I (I16479));
INVX1 gate6787(.O (g4794), .I (I8164));
INVX1 gate6788(.O (I11942), .I (g6909));
INVX1 gate6789(.O (I13773), .I (g8384));
INVX1 gate6790(.O (I5792), .I (g2080));
INVX1 gate6791(.O (g7442), .I (g7237));
INVX1 gate6792(.O (g8702), .I (g8664));
INVX1 gate6793(.O (I13341), .I (g8210));
INVX1 gate6794(.O (I12790), .I (g7618));
INVX1 gate6795(.O (g7786), .I (I12523));
INVX1 gate6796(.O (g2503), .I (g1872));
INVX1 gate6797(.O (g3757), .I (I6952));
INVX1 gate6798(.O (I9352), .I (g4944));
INVX1 gate6799(.O (I17312), .I (g11392));
INVX1 gate6800(.O (g10353), .I (I15823));
INVX1 gate6801(.O (g3416), .I (g3144));
INVX1 gate6802(.O (g6993), .I (I11135));
INVX1 gate6803(.O (I11180), .I (g6506));
INVX1 gate6804(.O (I16190), .I (g10493));
INVX1 gate6805(.O (I14485), .I (g8883));
INVX1 gate6806(.O (g7364), .I (I11740));
INVX1 gate6807(.O (I6815), .I (g2755));
INVX1 gate6808(.O (I9717), .I (g5426));
INVX1 gate6809(.O (I15551), .I (g10080));
INVX1 gate6810(.O (I14555), .I (g9009));
INVX1 gate6811(.O (g3522), .I (g3164));
INVX1 gate6812(.O (g8952), .I (I14309));
INVX1 gate6813(.O (g11572), .I (g11561));
INVX1 gate6814(.O (I11734), .I (g7024));
INVX1 gate6815(.O (g8276), .I (I13200));
INVX1 gate6816(.O (g3811), .I (I7029));
INVX1 gate6817(.O (g2224), .I (g695));
INVX1 gate6818(.O (I6097), .I (g2391));
INVX1 gate6819(.O (g5063), .I (g4363));
INVX1 gate6820(.O (I10914), .I (g6728));
INVX1 gate6821(.O (g7454), .I (g7148));
INVX1 gate6822(.O (I6726), .I (g3306));
INVX1 gate6823(.O (I14570), .I (g9028));
INVX1 gate6824(.O (I9893), .I (g5557));
INVX1 gate6825(.O (I13335), .I (g8206));
INVX1 gate6826(.O (g7770), .I (I12475));
INVX1 gate6827(.O (I14914), .I (g9533));
INVX1 gate6828(.O (g4515), .I (I7916));
INVX1 gate6829(.O (g4204), .I (I7429));
INVX1 gate6830(.O (I15127), .I (g9919));
INVX1 gate6831(.O (I16546), .I (g10724));
INVX1 gate6832(.O (g8561), .I (I13776));
INVX1 gate6833(.O (g2320), .I (g18));
INVX1 gate6834(.O (I10907), .I (g6705));
INVX1 gate6835(.O (g7725), .I (I12360));
INVX1 gate6836(.O (I8842), .I (g4556));
INVX1 gate6837(.O (g7532), .I (I11932));
INVX1 gate6838(.O (I7308), .I (g3070));
INVX1 gate6839(.O (g3874), .I (g2920));
INVX1 gate6840(.O (I8192), .I (g3566));
INVX1 gate6841(.O (I12208), .I (g7124));
INVX1 gate6842(.O (I8298), .I (g4437));
INVX1 gate6843(.O (I8085), .I (g3664));
INVX1 gate6844(.O (I13965), .I (g8451));
INVX1 gate6845(.O (g8004), .I (I12838));
INVX1 gate6846(.O (g6921), .I (I11037));
INVX1 gate6847(.O (g8986), .I (I14379));
INVX1 gate6848(.O (I5494), .I (g1690));
INVX1 gate6849(.O (I13131), .I (g7979));
INVX1 gate6850(.O (I14239), .I (g8803));
INVX1 gate6851(.O (I15956), .I (g10402));
INVX1 gate6852(.O (g2617), .I (g1997));
INVX1 gate6853(.O (g2906), .I (I6071));
INVX1 gate6854(.O (I14567), .I (g9027));
INVX1 gate6855(.O (g2789), .I (g2276));
INVX1 gate6856(.O (g5619), .I (g4840));
INVX1 gate6857(.O (g5167), .I (g4682));
INVX1 gate6858(.O (I15980), .I (g10414));
AN2X1 gate6859(.O (g11103), .I1 (g2250), .I2 (g10937));
AN2X1 gate6860(.O (g9900), .I1 (g9845), .I2 (g8327));
AN2X1 gate6861(.O (g11095), .I1 (g845), .I2 (g10950));
AN2X1 gate6862(.O (g3880), .I1 (g3186), .I2 (g2023));
AN2X1 gate6863(.O (g4973), .I1 (g1645), .I2 (g4467));
AN2X1 gate6864(.O (g7389), .I1 (g7001), .I2 (g3880));
AN2X1 gate6865(.O (g7888), .I1 (g7465), .I2 (g7025));
AN2X1 gate6866(.O (g4969), .I1 (g1642), .I2 (g4463));
AN2X1 gate6867(.O (g8224), .I1 (g1882), .I2 (g7887));
AN2X1 gate6868(.O (g2892), .I1 (g1980), .I2 (g1976));
AN2X1 gate6869(.O (g5686), .I1 (g158), .I2 (g5361));
AN2X1 gate6870(.O (g10308), .I1 (g10217), .I2 (g9085));
AN2X1 gate6871(.O (g4123), .I1 (g2695), .I2 (g3037));
AN2X1 gate6872(.O (g8120), .I1 (g1909), .I2 (g7944));
AN2X1 gate6873(.O (g6788), .I1 (g287), .I2 (g5876));
AN2X1 gate6874(.O (g5598), .I1 (g778), .I2 (g4824));
AN2X1 gate6875(.O (g9694), .I1 (g278), .I2 (g9432));
AN2X1 gate6876(.O (g10495), .I1 (g10431), .I2 (g3971));
AN2X1 gate6877(.O (g2945), .I1 (g2411), .I2 (g1684));
AN2X1 gate6878(.O (g11190), .I1 (g5623), .I2 (g11065));
AN2X1 gate6879(.O (g8789), .I1 (g8639), .I2 (g8719));
AN2X1 gate6880(.O (g9852), .I1 (g9728), .I2 (g9563));
AN2X1 gate6881(.O (g5625), .I1 (g1053), .I2 (g4399));
AN2X1 gate6882(.O (g4875), .I1 (g995), .I2 (g3914));
AN2X1 gate6883(.O (g9701), .I1 (g1574), .I2 (g9474));
AN2X1 gate6884(.O (g7138), .I1 (g6055), .I2 (g6707));
AN2X1 gate6885(.O (g10752), .I1 (g10692), .I2 (g3586));
AN2X1 gate6886(.O (g11211), .I1 (g11058), .I2 (g5534));
AN2X1 gate6887(.O (g11024), .I1 (g435), .I2 (g10974));
AN2X1 gate6888(.O (g8547), .I1 (g8307), .I2 (g7693));
AN2X1 gate6889(.O (g10669), .I1 (g10577), .I2 (g9429));
AN2X1 gate6890(.O (g7707), .I1 (g691), .I2 (g7206));
AN2X1 gate6891(.O (g4884), .I1 (g3813), .I2 (g2971));
AN2X1 gate6892(.O (g4839), .I1 (g225), .I2 (g3946));
AN2X1 gate6893(.O (g9870), .I1 (g1561), .I2 (g9816));
AN2X1 gate6894(.O (g6640), .I1 (g5281), .I2 (g5801));
AN2X1 gate6895(.O (g9650), .I1 (g2797), .I2 (g9240));
AN2X1 gate6896(.O (g5687), .I1 (g139), .I2 (g5361));
AN2X1 gate6897(.O (g7957), .I1 (g2885), .I2 (g7527));
AN2X1 gate6898(.O (g3512), .I1 (g2050), .I2 (g2971));
AN2X1 gate6899(.O (g8244), .I1 (g7847), .I2 (g4336));
AN2X1 gate6900(.O (g7449), .I1 (g6868), .I2 (g4355));
AN2X1 gate6901(.O (g4235), .I1 (g1011), .I2 (g3914));
AN2X1 gate6902(.O (g4343), .I1 (g345), .I2 (g3586));
AN2X1 gate6903(.O (g11296), .I1 (g5482), .I2 (g11241));
AN2X1 gate6904(.O (g9594), .I1 (g1), .I2 (g9292));
AN2X1 gate6905(.O (g6829), .I1 (g213), .I2 (g6596));
AN2X1 gate6906(.O (g4334), .I1 (g1160), .I2 (g3703));
AN2X1 gate6907(.O (g9943), .I1 (g9923), .I2 (g9367));
AN2X1 gate6908(.O (g5525), .I1 (g1721), .I2 (g4292));
AN2X1 gate6909(.O (g4548), .I1 (g440), .I2 (g3990));
AN3X1 gate6910(.O (g8876), .I1 (g8105), .I2 (g6764), .I3 (g8858));
AN2X1 gate6911(.O (g6733), .I1 (g5678), .I2 (g4324));
AN2X1 gate6912(.O (g4804), .I1 (g476), .I2 (g3458));
AN2X1 gate6913(.O (g10705), .I1 (g10564), .I2 (g4840));
AN2X1 gate6914(.O (g9934), .I1 (g9913), .I2 (g9624));
AN2X1 gate6915(.O (g6225), .I1 (g566), .I2 (g5082));
AN2X1 gate6916(.O (g6324), .I1 (g1240), .I2 (g5949));
AN2X1 gate6917(.O (g10686), .I1 (g10612), .I2 (g3863));
AN2X1 gate6918(.O (g6540), .I1 (g1223), .I2 (g6072));
AN2X1 gate6919(.O (g8663), .I1 (g8538), .I2 (g4013));
AN2X1 gate6920(.O (g11581), .I1 (g1308), .I2 (g11539));
AN2X1 gate6921(.O (g6206), .I1 (g560), .I2 (g5068));
AN2X1 gate6922(.O (g4518), .I1 (g452), .I2 (g3975));
AN2X1 gate6923(.O (g3989), .I1 (g248), .I2 (g3164));
AN2X1 gate6924(.O (g7730), .I1 (g7260), .I2 (g2347));
AN2X1 gate6925(.O (g5174), .I1 (g1235), .I2 (g4681));
AN2X1 gate6926(.O (g7504), .I1 (g7148), .I2 (g2847));
AN2X1 gate6927(.O (g7185), .I1 (g1887), .I2 (g6724));
AN2X1 gate6928(.O (g2563), .I1 (I5689), .I2 (I5690));
AN2X1 gate6929(.O (g7881), .I1 (g7612), .I2 (g3810));
AN2X1 gate6930(.O (g11070), .I1 (g2008), .I2 (g10913));
AN2X1 gate6931(.O (g9859), .I1 (g9736), .I2 (g9573));
AN3X1 gate6932(.O (g8877), .I1 (g8103), .I2 (g6764), .I3 (g8858));
AN2X1 gate6933(.O (g11590), .I1 (g2274), .I2 (g11561));
AN2X1 gate6934(.O (g6199), .I1 (g557), .I2 (g5062));
AN2X1 gate6935(.O (g9266), .I1 (g8932), .I2 (g3398));
AN2X1 gate6936(.O (g5545), .I1 (g1730), .I2 (g4321));
AN2X1 gate6937(.O (g5180), .I1 (g4541), .I2 (g4533));
AN2X1 gate6938(.O (g5591), .I1 (g1615), .I2 (g4514));
AN2X1 gate6939(.O (g8556), .I1 (g8412), .I2 (g8029));
AN2X1 gate6940(.O (g11094), .I1 (g374), .I2 (g10883));
AN2X1 gate6941(.O (g5853), .I1 (g5044), .I2 (g1927));
AN2X1 gate6942(.O (g6245), .I1 (g575), .I2 (g5098));
AN2X1 gate6943(.O (g4360), .I1 (g1861), .I2 (g3748));
AN3X1 gate6944(.O (g8930), .I1 (g8100), .I2 (g6368), .I3 (g8828));
AN2X1 gate6945(.O (g5507), .I1 (g4310), .I2 (g3528));
AN2X1 gate6946(.O (g11150), .I1 (g3087), .I2 (g10913));
AN2X1 gate6947(.O (g8464), .I1 (g8302), .I2 (g7416));
AN2X1 gate6948(.O (g9692), .I1 (g272), .I2 (g9432));
AN2X1 gate6949(.O (g4996), .I1 (g1428), .I2 (g4682));
AN2X1 gate6950(.O (g7131), .I1 (g6044), .I2 (g6700));
AN2X1 gate6951(.O (g11019), .I1 (g421), .I2 (g10974));
AN2X1 gate6952(.O (g9960), .I1 (g9951), .I2 (g9536));
AN2X1 gate6953(.O (g11196), .I1 (g4912), .I2 (g11068));
AN2X1 gate6954(.O (g11018), .I1 (g7286), .I2 (g10974));
AN2X1 gate6955(.O (g6819), .I1 (g243), .I2 (g6596));
AN2X1 gate6956(.O (g10595), .I1 (g10550), .I2 (g4347));
AN2X1 gate6957(.O (g10494), .I1 (g10433), .I2 (g3945));
AN2X1 gate6958(.O (g10623), .I1 (g10544), .I2 (g4536));
AN2X1 gate6959(.O (g4878), .I1 (g1868), .I2 (g3531));
AN2X1 gate6960(.O (g5204), .I1 (g4838), .I2 (g2126));
AN2X1 gate6961(.O (g8844), .I1 (g8609), .I2 (g8709));
AN2X1 gate6962(.O (g6701), .I1 (g6185), .I2 (g4228));
AN2X1 gate6963(.O (g10782), .I1 (g10725), .I2 (g5146));
AN2X1 gate6964(.O (g5100), .I1 (g1791), .I2 (g4606));
AN2X1 gate6965(.O (g4882), .I1 (g1089), .I2 (g3638));
AN2X1 gate6966(.O (g8731), .I1 (g8622), .I2 (g7918));
AN2X1 gate6967(.O (g6215), .I1 (g1504), .I2 (g5128));
AN2X1 gate6968(.O (g6886), .I1 (g1932), .I2 (g6420));
AN2X1 gate6969(.O (g3586), .I1 (g3323), .I2 (g2191));
AN2X1 gate6970(.O (g8557), .I1 (g8415), .I2 (g8033));
AN3X1 gate6971(.O (g8966), .I1 (g8081), .I2 (g6778), .I3 (g8849));
AN2X1 gate6972(.O (g8071), .I1 (g691), .I2 (g7826));
AN2X1 gate6973(.O (g11597), .I1 (g11576), .I2 (g5446));
AN2X1 gate6974(.O (g9828), .I1 (g9722), .I2 (g9785));
AN2X1 gate6975(.O (g2918), .I1 (g2411), .I2 (g1672));
AN2X1 gate6976(.O (g9830), .I1 (g9725), .I2 (g9785));
AN3X1 gate6977(.O (g8955), .I1 (g8110), .I2 (g6368), .I3 (g8828));
AN2X1 gate6978(.O (g9592), .I1 (g4), .I2 (g9292));
AN2X1 gate6979(.O (g5123), .I1 (g1618), .I2 (g4669));
AN2X1 gate6980(.O (g7059), .I1 (g6078), .I2 (g6714));
AN2X1 gate6981(.O (g8254), .I1 (g2773), .I2 (g7909));
AN2X1 gate6982(.O (g7459), .I1 (g7148), .I2 (g2814));
AN2X1 gate6983(.O (g11102), .I1 (g861), .I2 (g10950));
AN2X1 gate6984(.O (g7718), .I1 (g709), .I2 (g7221));
AN2X1 gate6985(.O (g7535), .I1 (g7148), .I2 (g2874));
AN2X1 gate6986(.O (g9703), .I1 (g1577), .I2 (g9474));
AN2X1 gate6987(.O (g5528), .I1 (g4322), .I2 (g3537));
AN2X1 gate6988(.O (g5151), .I1 (g4478), .I2 (g2733));
AN2X1 gate6989(.O (g9932), .I1 (g9911), .I2 (g9624));
AN2X1 gate6990(.O (g5530), .I1 (g1636), .I2 (g4305));
AN2X1 gate6991(.O (g3506), .I1 (g986), .I2 (g2760));
AN2X1 gate6992(.O (g8769), .I1 (g8629), .I2 (g5151));
AN2X1 gate6993(.O (g6887), .I1 (g6187), .I2 (g6566));
AN2X1 gate6994(.O (g6228), .I1 (g5605), .I2 (g713));
AN2X1 gate6995(.O (g6322), .I1 (g1275), .I2 (g5949));
AN2X1 gate6996(.O (g3111), .I1 (I6337), .I2 (I6338));
AN3X1 gate6997(.O (g8967), .I1 (g8085), .I2 (g6778), .I3 (g8849));
AN2X1 gate6998(.O (g5010), .I1 (g1458), .I2 (g4640));
AN2X1 gate6999(.O (g3275), .I1 (g115), .I2 (g2356));
AN2X1 gate7000(.O (g10809), .I1 (g4811), .I2 (g10754));
AN2X1 gate7001(.O (g2895), .I1 (g2411), .I2 (g1678));
AN2X1 gate7002(.O (g7721), .I1 (g736), .I2 (g7237));
AN2X1 gate7003(.O (g9866), .I1 (g1549), .I2 (g9802));
AN2X1 gate7004(.O (g9716), .I1 (g1534), .I2 (g9490));
AN2X1 gate7005(.O (g10808), .I1 (g10744), .I2 (g3829));
AN2X1 gate7006(.O (g3374), .I1 (g1231), .I2 (g3047));
AN2X1 gate7007(.O (g4492), .I1 (g1786), .I2 (g3685));
AN2X1 gate7008(.O (g8822), .I1 (g8614), .I2 (g8752));
AN2X1 gate7009(.O (g10560), .I1 (g10487), .I2 (g4575));
AN3X1 gate7010(.O (g11456), .I1 (g3765), .I2 (g3517), .I3 (g11422));
AN2X1 gate7011(.O (g9848), .I1 (g9724), .I2 (g9557));
AN2X1 gate7012(.O (g4714), .I1 (g646), .I2 (g3333));
AN2X1 gate7013(.O (g6550), .I1 (g1231), .I2 (g6089));
AN2X1 gate7014(.O (g5172), .I1 (g4555), .I2 (g4549));
AN2X1 gate7015(.O (g10642), .I1 (g10612), .I2 (g3829));
AN2X1 gate7016(.O (g3284), .I1 (g2531), .I2 (g677));
AN2X1 gate7017(.O (g9699), .I1 (g284), .I2 (g9432));
AN2X1 gate7018(.O (g9855), .I1 (g302), .I2 (g9772));
AN2X1 gate7019(.O (g5618), .I1 (g1630), .I2 (g4551));
AN2X1 gate7020(.O (g6891), .I1 (g1950), .I2 (g6435));
AN2X1 gate7021(.O (g7940), .I1 (g7620), .I2 (g4013));
AN2X1 gate7022(.O (g11085), .I1 (g312), .I2 (g10897));
AN2X1 gate7023(.O (g4736), .I1 (g396), .I2 (g3379));
AN2X1 gate7024(.O (g4968), .I1 (g1432), .I2 (g4682));
AN2X1 gate7025(.O (g8837), .I1 (g8646), .I2 (g8697));
AN2X1 gate7026(.O (g9644), .I1 (g1182), .I2 (g9125));
AN2X1 gate7027(.O (g5804), .I1 (g1546), .I2 (g5261));
AN2X1 gate7028(.O (g8462), .I1 (g8300), .I2 (g7406));
AN4X1 gate7029(.O (I6330), .I1 (g2549), .I2 (g2556), .I3 (g2562), .I4 (g2570));
AN2X1 gate7030(.O (g11156), .I1 (g333), .I2 (g10934));
AN2X1 gate7031(.O (g6342), .I1 (g293), .I2 (g5886));
AN2X1 gate7032(.O (g9867), .I1 (g1552), .I2 (g9807));
AN2X1 gate7033(.O (g9717), .I1 (g1537), .I2 (g9490));
AN2X1 gate7034(.O (g4871), .I1 (g1864), .I2 (g3523));
AN2X1 gate7035(.O (g10454), .I1 (g10435), .I2 (g3411));
AN2X1 gate7036(.O (g4722), .I1 (g426), .I2 (g3353));
AN2X1 gate7037(.O (g7741), .I1 (g6961), .I2 (g3880));
AN2X1 gate7038(.O (g4500), .I1 (g1357), .I2 (g3941));
AN2X1 gate7039(.O (g9386), .I1 (g1327), .I2 (g9151));
AN2X1 gate7040(.O (g8842), .I1 (g8607), .I2 (g8707));
AN2X1 gate7041(.O (g9599), .I1 (g8), .I2 (g9292));
AN2X1 gate7042(.O (g9274), .I1 (g8974), .I2 (g5708));
AN2X1 gate7043(.O (g5518), .I1 (g4317), .I2 (g3532));
AN2X1 gate7044(.O (g9614), .I1 (g1197), .I2 (g9111));
AN2X1 gate7045(.O (g4838), .I1 (g3275), .I2 (g4122));
AN2X1 gate7046(.O (g9125), .I1 (g8966), .I2 (g6674));
AN2X1 gate7047(.O (g7217), .I1 (g4610), .I2 (g6432));
AN2X1 gate7048(.O (g11557), .I1 (g2707), .I2 (g11519));
AN2X1 gate7049(.O (g2911), .I1 (g2411), .I2 (g1675));
AN2X1 gate7050(.O (g11210), .I1 (g11078), .I2 (g4515));
AN2X1 gate7051(.O (g7466), .I1 (g7148), .I2 (g2821));
AN2X1 gate7052(.O (g9939), .I1 (g9918), .I2 (g9367));
AN2X1 gate7053(.O (g11279), .I1 (g4939), .I2 (g11200));
AN3X1 gate7054(.O (g10518), .I1 (g10513), .I2 (g10440), .I3 (I16145));
AN2X1 gate7055(.O (g4477), .I1 (g1129), .I2 (g3878));
AN2X1 gate7056(.O (g8708), .I1 (g7605), .I2 (g8592));
AN2X1 gate7057(.O (g7055), .I1 (g5900), .I2 (g6579));
AN2X1 gate7058(.O (g5264), .I1 (g1095), .I2 (g4763));
AN2X1 gate7059(.O (g6329), .I1 (g1265), .I2 (g5949));
AN2X1 gate7060(.O (g6828), .I1 (g1377), .I2 (g6596));
AN2X1 gate7061(.O (g8176), .I1 (g5299), .I2 (g7853));
AN2X1 gate7062(.O (g6830), .I1 (g1380), .I2 (g6596));
AN2X1 gate7063(.O (g8005), .I1 (g7510), .I2 (g6871));
AN2X1 gate7064(.O (g4099), .I1 (g770), .I2 (g3281));
AN2X1 gate7065(.O (g11601), .I1 (g1351), .I2 (g11574));
AN2X1 gate7066(.O (g11187), .I1 (g5597), .I2 (g11061));
AN2X1 gate7067(.O (g6746), .I1 (g6228), .I2 (g6166));
AN2X1 gate7068(.O (g6221), .I1 (g782), .I2 (g5598));
AN2X1 gate7069(.O (g8765), .I1 (g8630), .I2 (g5151));
AN2X1 gate7070(.O (g9622), .I1 (g1200), .I2 (g9111));
AN2X1 gate7071(.O (g11143), .I1 (g10923), .I2 (g4567));
AN2X1 gate7072(.O (g9904), .I1 (g9886), .I2 (g9676));
AN2X1 gate7073(.O (g8733), .I1 (g8625), .I2 (g7920));
AN3X1 gate7074(.O (g8974), .I1 (g8094), .I2 (g6368), .I3 (g8858));
AN2X1 gate7075(.O (g6624), .I1 (g348), .I2 (g6171));
AN2X1 gate7076(.O (g11169), .I1 (g530), .I2 (g11112));
AN2X1 gate7077(.O (g8073), .I1 (g709), .I2 (g7826));
AN2X1 gate7078(.O (g9841), .I1 (g9706), .I2 (g9512));
AN2X1 gate7079(.O (g5882), .I1 (g5592), .I2 (g3829));
AN2X1 gate7080(.O (g8796), .I1 (g8645), .I2 (g8725));
AN2X1 gate7081(.O (g11168), .I1 (g534), .I2 (g11112));
AN2X1 gate7082(.O (g4269), .I1 (g1015), .I2 (g3914));
AN2X1 gate7083(.O (g5271), .I1 (g727), .I2 (g4772));
AN2X1 gate7084(.O (g10348), .I1 (g10272), .I2 (g3705));
AN2X1 gate7085(.O (g5611), .I1 (g1047), .I2 (g4382));
AN2X1 gate7086(.O (g8069), .I1 (g673), .I2 (g7826));
AN2X1 gate7087(.O (g9695), .I1 (g1567), .I2 (g9474));
AN2X1 gate7088(.O (g10304), .I1 (g10211), .I2 (g9079));
AN2X1 gate7089(.O (g8469), .I1 (g8305), .I2 (g7422));
AN2X1 gate7090(.O (g4712), .I1 (g1071), .I2 (g3638));
AN2X1 gate7091(.O (g6576), .I1 (g5762), .I2 (g5503));
AN2X1 gate7092(.O (g10622), .I1 (g10543), .I2 (g4525));
AN2X1 gate7093(.O (g11015), .I1 (g5217), .I2 (g10827));
AN2X1 gate7094(.O (g5674), .I1 (g148), .I2 (g5361));
AN2X1 gate7095(.O (g9359), .I1 (g1308), .I2 (g9173));
AN2X1 gate7096(.O (g9223), .I1 (g6454), .I2 (g8960));
AN2X1 gate7097(.O (g11556), .I1 (g2701), .I2 (g11519));
AN2X1 gate7098(.O (g9858), .I1 (g1595), .I2 (g9774));
AN2X1 gate7099(.O (g5541), .I1 (g4331), .I2 (g3582));
AN2X1 gate7100(.O (g4534), .I1 (g363), .I2 (g3586));
AN2X1 gate7101(.O (g6198), .I1 (g1499), .I2 (g5128));
AN2X1 gate7102(.O (g6747), .I1 (g2214), .I2 (g5897));
AN2X1 gate7103(.O (g6699), .I1 (g6177), .I2 (g4221));
AN2X1 gate7104(.O (g6855), .I1 (g1964), .I2 (g6392));
AN2X1 gate7105(.O (g3804), .I1 (g3098), .I2 (g2203));
AN2X1 gate7106(.O (g5680), .I1 (g153), .I2 (g5361));
AN2X1 gate7107(.O (g9642), .I1 (g2654), .I2 (g9240));
AN2X1 gate7108(.O (g5744), .I1 (g1528), .I2 (g5191));
AN2X1 gate7109(.O (g10333), .I1 (g10262), .I2 (g3307));
AN2X1 gate7110(.O (g8399), .I1 (g6094), .I2 (g8229));
AN2X1 gate7111(.O (g9447), .I1 (g1762), .I2 (g9030));
AN2X1 gate7112(.O (g4903), .I1 (g1849), .I2 (g4243));
AN2X1 gate7113(.O (g11178), .I1 (g516), .I2 (g11112));
AN2X1 gate7114(.O (g8510), .I1 (g8414), .I2 (g7972));
AN2X1 gate7115(.O (g8245), .I1 (g7850), .I2 (g4339));
AN2X1 gate7116(.O (g6319), .I1 (g1296), .I2 (g5949));
AN2X1 gate7117(.O (g11186), .I1 (g5594), .I2 (g11059));
AN2X1 gate7118(.O (g3908), .I1 (g186), .I2 (g3164));
AN2X1 gate7119(.O (g2951), .I1 (g2411), .I2 (g1681));
AN2X1 gate7120(.O (g6352), .I1 (g278), .I2 (g5894));
AN2X1 gate7121(.O (g9595), .I1 (g901), .I2 (g9205));
AN2X1 gate7122(.O (g4831), .I1 (g810), .I2 (g4109));
AN2X1 gate7123(.O (g5492), .I1 (g1654), .I2 (g4263));
AN2X1 gate7124(.O (g9272), .I1 (g8934), .I2 (g3424));
AN2X1 gate7125(.O (g10312), .I1 (g10220), .I2 (g9094));
AN2X1 gate7126(.O (g6186), .I1 (g546), .I2 (g5042));
AN2X1 gate7127(.O (g9612), .I1 (g2652), .I2 (g9240));
AN2X1 gate7128(.O (g9417), .I1 (g1738), .I2 (g9052));
AN2X1 gate7129(.O (g9935), .I1 (g9914), .I2 (g9624));
AN2X1 gate7130(.O (g8701), .I1 (g7597), .I2 (g8582));
AN2X1 gate7131(.O (g10745), .I1 (g10658), .I2 (g3586));
AN2X1 gate7132(.O (g11216), .I1 (g956), .I2 (g11162));
AN2X1 gate7133(.O (g9328), .I1 (g8971), .I2 (g5708));
AN2X1 gate7134(.O (g11587), .I1 (g1327), .I2 (g11546));
AN2X1 gate7135(.O (g6821), .I1 (g237), .I2 (g6596));
AN2X1 gate7136(.O (g6325), .I1 (g1245), .I2 (g5949));
AN2X1 gate7137(.O (g4560), .I1 (g431), .I2 (g4002));
AN2X1 gate7138(.O (g7368), .I1 (g6980), .I2 (g3880));
AN2X1 gate7139(.O (g6083), .I1 (g552), .I2 (g5619));
AN2X1 gate7140(.O (g6544), .I1 (g1227), .I2 (g6081));
AN2X1 gate7141(.O (g5476), .I1 (g1615), .I2 (g4237));
AN2X1 gate7142(.O (g7743), .I1 (g6967), .I2 (g3880));
AN2X1 gate7143(.O (g4869), .I1 (g1083), .I2 (g3638));
AN2X1 gate7144(.O (g5722), .I1 (g1598), .I2 (g5144));
AN2X1 gate7145(.O (g6790), .I1 (g5813), .I2 (g4398));
AN2X1 gate7146(.O (g8408), .I1 (g704), .I2 (g8139));
AN2X1 gate7147(.O (g10761), .I1 (g10700), .I2 (g10699));
AN2X1 gate7148(.O (g7734), .I1 (g6944), .I2 (g3880));
AN2X1 gate7149(.O (g8136), .I1 (g7926), .I2 (g7045));
AN2X1 gate7150(.O (g6187), .I1 (g5569), .I2 (g2340));
AN2X1 gate7151(.O (g4752), .I1 (g401), .I2 (g3385));
AN2X1 gate7152(.O (g9902), .I1 (g9894), .I2 (g9392));
AN2X1 gate7153(.O (g8768), .I1 (g8623), .I2 (g5151));
AN2X1 gate7154(.O (g5500), .I1 (g1657), .I2 (g4272));
AN2X1 gate7155(.O (g2496), .I1 (g374), .I2 (g369));
AN2X1 gate7156(.O (g6756), .I1 (g3010), .I2 (g5877));
AN3X1 gate7157(.O (g8972), .I1 (g8085), .I2 (g6764), .I3 (g8858));
AN2X1 gate7158(.O (g6622), .I1 (g336), .I2 (g6165));
AN2X1 gate7159(.O (g11639), .I1 (g11612), .I2 (g7897));
AN2X1 gate7160(.O (g9366), .I1 (g1311), .I2 (g9173));
AN2X1 gate7161(.O (g11230), .I1 (g471), .I2 (g11062));
AN2X1 gate7162(.O (g10328), .I1 (g10252), .I2 (g3307));
AN2X1 gate7163(.O (g5024), .I1 (g1284), .I2 (g4513));
AN2X1 gate7164(.O (g4364), .I1 (g1215), .I2 (g3756));
AN2X1 gate7165(.O (g9649), .I1 (g916), .I2 (g9205));
AN2X1 gate7166(.O (g5795), .I1 (g1543), .I2 (g5251));
AN2X1 gate7167(.O (g5737), .I1 (g1524), .I2 (g5183));
AN2X1 gate7168(.O (g6841), .I1 (g1400), .I2 (g6596));
AN2X1 gate7169(.O (g4054), .I1 (g1753), .I2 (g2793));
AN2X1 gate7170(.O (g6345), .I1 (g5823), .I2 (g4426));
AN2X1 gate7171(.O (g11391), .I1 (g11275), .I2 (g7912));
AN2X1 gate7172(.O (g9851), .I1 (g296), .I2 (g9770));
AN2X1 gate7173(.O (g6763), .I1 (g5802), .I2 (g4381));
AN2X1 gate7174(.O (g4770), .I1 (g416), .I2 (g3415));
AN3X1 gate7175(.O (I16142), .I1 (g10511), .I2 (g10509), .I3 (g10507));
AN2X1 gate7176(.O (g9698), .I1 (g1571), .I2 (g9474));
AN2X1 gate7177(.O (g4725), .I1 (g1032), .I2 (g3914));
AN2X1 gate7178(.O (g5477), .I1 (g1887), .I2 (g4241));
AN2X1 gate7179(.O (g9964), .I1 (g9954), .I2 (g9536));
AN2X1 gate7180(.O (g5523), .I1 (g1663), .I2 (g4290));
AN2X1 gate7181(.O (g4553), .I1 (g435), .I2 (g3995));
AN2X1 gate7182(.O (g8550), .I1 (g8402), .I2 (g8011));
AN2X1 gate7183(.O (g8845), .I1 (g8611), .I2 (g8711));
AN2X1 gate7184(.O (g2081), .I1 (g932), .I2 (g928));
AN2X1 gate7185(.O (g6359), .I1 (g281), .I2 (g5898));
AN2X1 gate7186(.O (g11586), .I1 (g1324), .I2 (g11545));
AN2X1 gate7187(.O (g11007), .I1 (g5147), .I2 (g10827));
AN2X1 gate7188(.O (g5104), .I1 (g1796), .I2 (g4608));
AN2X1 gate7189(.O (g5099), .I1 (g4821), .I2 (g3829));
AN2X1 gate7190(.O (g6757), .I1 (g2221), .I2 (g5919));
AN2X1 gate7191(.O (g5499), .I1 (g1627), .I2 (g4270));
AN2X1 gate7192(.O (g4389), .I1 (g3529), .I2 (g3092));
AN2X1 gate7193(.O (g6416), .I1 (g3497), .I2 (g5774));
AN2X1 gate7194(.O (g9720), .I1 (g1546), .I2 (g9490));
AN2X1 gate7195(.O (g4990), .I1 (g1444), .I2 (g4682));
AN2X1 gate7196(.O (g9619), .I1 (g2772), .I2 (g9010));
AN4X1 gate7197(.O (I6630), .I1 (g2677), .I2 (g2683), .I3 (g2689), .I4 (g2701));
AN2X1 gate7198(.O (g6047), .I1 (g2017), .I2 (g4977));
AN2X1 gate7199(.O (g9652), .I1 (g953), .I2 (g9223));
AN3X1 gate7200(.O (g10515), .I1 (g10505), .I2 (g10469), .I3 (I16142));
AN2X1 gate7201(.O (g9843), .I1 (g9711), .I2 (g9519));
AN2X1 gate7202(.O (g5273), .I1 (g1074), .I2 (g4776));
AN2X1 gate7203(.O (g11465), .I1 (g11434), .I2 (g5446));
AN2X1 gate7204(.O (g5044), .I1 (g4348), .I2 (g1918));
AN2X1 gate7205(.O (g11237), .I1 (g5472), .I2 (g11109));
AN2X1 gate7206(.O (g9834), .I1 (g9731), .I2 (g9785));
AN2X1 gate7207(.O (g6654), .I1 (g363), .I2 (g6214));
AN2X1 gate7208(.O (g5444), .I1 (g1041), .I2 (g4880));
AN2X1 gate7209(.O (g3714), .I1 (g1690), .I2 (g2991));
AN2X1 gate7210(.O (g11340), .I1 (g11285), .I2 (g4424));
AN2X1 gate7211(.O (g9598), .I1 (g2086), .I2 (g9274));
AN2X1 gate7212(.O (g8097), .I1 (g6200), .I2 (g7851));
AN2X1 gate7213(.O (g8726), .I1 (g8608), .I2 (g7913));
AN2X1 gate7214(.O (g6880), .I1 (g4816), .I2 (g6562));
AN2X1 gate7215(.O (g4338), .I1 (g1157), .I2 (g3707));
AN2X1 gate7216(.O (g5543), .I1 (g4874), .I2 (g4312));
AN3X1 gate7217(.O (g8960), .I1 (g8085), .I2 (g6368), .I3 (g8828));
AN2X1 gate7218(.O (g4109), .I1 (g806), .I2 (g3287));
AN2X1 gate7219(.O (g10759), .I1 (g10698), .I2 (g10697));
AN2X1 gate7220(.O (g9938), .I1 (g9917), .I2 (g9367));
AN2X1 gate7221(.O (g10758), .I1 (g10652), .I2 (g4013));
AN2X1 gate7222(.O (g4759), .I1 (g406), .I2 (g3392));
AN2X1 gate7223(.O (g9909), .I1 (g9891), .I2 (g9804));
AN2X1 gate7224(.O (g7127), .I1 (g6663), .I2 (g2241));
AN2X1 gate7225(.O (g11165), .I1 (g476), .I2 (g11112));
AN2X1 gate7226(.O (g6234), .I1 (g2244), .I2 (g5151));
AN2X1 gate7227(.O (g6328), .I1 (g1260), .I2 (g5949));
AN2X1 gate7228(.O (g8401), .I1 (g677), .I2 (g8124));
AN2X1 gate7229(.O (g11006), .I1 (g5125), .I2 (g10827));
AN2X1 gate7230(.O (g4865), .I1 (g1080), .I2 (g3638));
AN2X1 gate7231(.O (g4715), .I1 (g1077), .I2 (g3638));
AN3X1 gate7232(.O (g4604), .I1 (g3056), .I2 (g3753), .I3 (g2325));
AN2X1 gate7233(.O (g5513), .I1 (g1675), .I2 (g4282));
AN2X1 gate7234(.O (g11222), .I1 (g965), .I2 (g11055));
AN2X1 gate7235(.O (g4498), .I1 (g1145), .I2 (g3940));
AN2X1 gate7236(.O (g6554), .I1 (g5075), .I2 (g6183));
AN2X1 gate7237(.O (g7732), .I1 (g6935), .I2 (g3880));
AN2X1 gate7238(.O (g9586), .I1 (g2727), .I2 (g9173));
AN3X1 gate7239(.O (g5178), .I1 (g2047), .I2 (g4401), .I3 (g4104));
AN2X1 gate7240(.O (g4584), .I1 (g3710), .I2 (g2322));
AN2X1 gate7241(.O (g7472), .I1 (g7148), .I2 (g2829));
AN2X1 gate7242(.O (g11253), .I1 (g981), .I2 (g11072));
AN2X1 gate7243(.O (g5182), .I1 (g1240), .I2 (g4713));
AN2X1 gate7244(.O (g9860), .I1 (g1598), .I2 (g9775));
AN2X1 gate7245(.O (g8703), .I1 (g7601), .I2 (g8585));
AN2X1 gate7246(.O (g11600), .I1 (g1346), .I2 (g11573));
AN2X1 gate7247(.O (g9710), .I1 (g1586), .I2 (g9474));
AN2X1 gate7248(.O (g9645), .I1 (g1203), .I2 (g9111));
AN2X1 gate7249(.O (g11236), .I1 (g5469), .I2 (g11108));
AN2X1 gate7250(.O (g4162), .I1 (g3106), .I2 (g2971));
AN2X1 gate7251(.O (g6090), .I1 (g553), .I2 (g5627));
AN2X1 gate7252(.O (g9691), .I1 (g269), .I2 (g9432));
AN2X1 gate7253(.O (g11372), .I1 (g11316), .I2 (g4266));
AN2X1 gate7254(.O (g6823), .I1 (g1368), .I2 (g6596));
AN2X1 gate7255(.O (g11175), .I1 (g501), .I2 (g11112));
AN2X1 gate7256(.O (g8068), .I1 (g664), .I2 (g7826));
AN2X1 gate7257(.O (g9607), .I1 (g12), .I2 (g9274));
AN2X1 gate7258(.O (g9962), .I1 (g9952), .I2 (g9536));
AN2X1 gate7259(.O (g6348), .I1 (g296), .I2 (g5891));
AN2X1 gate7260(.O (g9659), .I1 (g956), .I2 (g9223));
AN2X1 gate7261(.O (g9358), .I1 (g1318), .I2 (g9151));
AN2X1 gate7262(.O (g3104), .I1 (I6316), .I2 (I6317));
AN2X1 gate7263(.O (g4486), .I1 (g1711), .I2 (g3910));
AN2X1 gate7264(.O (g9587), .I1 (g892), .I2 (g8995));
AN2X1 gate7265(.O (g5632), .I1 (g1636), .I2 (g4563));
AN2X1 gate7266(.O (g9111), .I1 (g8965), .I2 (g6674));
AN2X1 gate7267(.O (g4881), .I1 (g991), .I2 (g3914));
AN2X1 gate7268(.O (g11209), .I1 (g11074), .I2 (g9448));
AN2X1 gate7269(.O (g8848), .I1 (g8715), .I2 (g8713));
AN2X1 gate7270(.O (g4070), .I1 (g3263), .I2 (g2330));
AN2X1 gate7271(.O (g6463), .I1 (g5052), .I2 (g6210));
AN2X1 gate7272(.O (g8699), .I1 (g7595), .I2 (g8579));
AN4X1 gate7273(.O (I5689), .I1 (g1419), .I2 (g1424), .I3 (g1428), .I4 (g1432));
AN2X1 gate7274(.O (g7820), .I1 (g1896), .I2 (g7479));
AN2X1 gate7275(.O (g11021), .I1 (g448), .I2 (g10974));
AN2X1 gate7276(.O (g5917), .I1 (g1044), .I2 (g5320));
AN2X1 gate7277(.O (g6619), .I1 (g49), .I2 (g6156));
AN2X1 gate7278(.O (g6318), .I1 (g1300), .I2 (g5949));
AN2X1 gate7279(.O (g6872), .I1 (g1896), .I2 (g6389));
AN2X1 gate7280(.O (g11320), .I1 (g11201), .I2 (g4379));
AN2X1 gate7281(.O (g10514), .I1 (g10489), .I2 (g4580));
AN2X1 gate7282(.O (g4006), .I1 (g201), .I2 (g3228));
AN2X1 gate7283(.O (g9853), .I1 (g299), .I2 (g9771));
AN2X1 gate7284(.O (g11274), .I1 (g4913), .I2 (g11197));
AN2X1 gate7285(.O (g6193), .I1 (g2206), .I2 (g5151));
AN2X1 gate7286(.O (g8119), .I1 (g6239), .I2 (g7890));
AN2X1 gate7287(.O (g9420), .I1 (g1747), .I2 (g9030));
AN2X1 gate7288(.O (g5233), .I1 (g1791), .I2 (g4492));
AN2X1 gate7289(.O (g7581), .I1 (g7092), .I2 (g5420));
AN2X1 gate7290(.O (g6549), .I1 (g5515), .I2 (g6175));
AN2X1 gate7291(.O (g11464), .I1 (g11433), .I2 (g5446));
AN2X1 gate7292(.O (g4801), .I1 (g516), .I2 (g3439));
AN2X1 gate7293(.O (g6834), .I1 (g1365), .I2 (g6596));
AN2X1 gate7294(.O (g4487), .I1 (g1718), .I2 (g3911));
AN2X1 gate7295(.O (g2939), .I1 (g2411), .I2 (g1687));
AN2X1 gate7296(.O (g7060), .I1 (g6739), .I2 (g5521));
AN2X1 gate7297(.O (g5770), .I1 (g4466), .I2 (g5128));
AN2X1 gate7298(.O (g5725), .I1 (g1580), .I2 (g5166));
AN2X1 gate7299(.O (g11641), .I1 (g11615), .I2 (g7901));
AN2X1 gate7300(.O (g2544), .I1 (g1341), .I2 (g1336));
AN2X1 gate7301(.O (g11292), .I1 (g11252), .I2 (g4250));
AN2X1 gate7302(.O (g5532), .I1 (g1681), .I2 (g4307));
AN2X1 gate7303(.O (g11153), .I1 (g3771), .I2 (g10913));
AN2X1 gate7304(.O (g9905), .I1 (g9872), .I2 (g9680));
AN2X1 gate7305(.O (g7739), .I1 (g6957), .I2 (g3880));
AN2X1 gate7306(.O (g6321), .I1 (g1284), .I2 (g5949));
AN2X1 gate7307(.O (g8386), .I1 (g6085), .I2 (g8219));
AN3X1 gate7308(.O (g8975), .I1 (g8089), .I2 (g6764), .I3 (g8858));
AN2X1 gate7309(.O (g2306), .I1 (g1223), .I2 (g1218));
AN2X1 gate7310(.O (g6625), .I1 (g1218), .I2 (g6178));
AN2X1 gate7311(.O (g7937), .I1 (g7606), .I2 (g4013));
AN2X1 gate7312(.O (g10788), .I1 (g8303), .I2 (g10754));
AN2X1 gate7313(.O (g10325), .I1 (g10248), .I2 (g3307));
AN2X1 gate7314(.O (g8170), .I1 (g5270), .I2 (g7853));
AN2X1 gate7315(.O (g5706), .I1 (g1574), .I2 (g5121));
AN2X1 gate7316(.O (g2756), .I1 (g936), .I2 (g2081));
AN2X1 gate7317(.O (g8821), .I1 (g8643), .I2 (g8751));
AN2X1 gate7318(.O (g10946), .I1 (g5225), .I2 (g10827));
AN2X1 gate7319(.O (g4169), .I1 (g2765), .I2 (g3066));
AN2X1 gate7320(.O (g5029), .I1 (g1077), .I2 (g4521));
AN2X1 gate7321(.O (g11164), .I1 (g4889), .I2 (g11112));
AN2X1 gate7322(.O (g4007), .I1 (g2683), .I2 (g2276));
AN2X1 gate7323(.O (g4059), .I1 (g1756), .I2 (g2796));
AN2X1 gate7324(.O (g4868), .I1 (g1027), .I2 (g3914));
AN2X1 gate7325(.O (g5675), .I1 (g131), .I2 (g5361));
AN2X1 gate7326(.O (g4718), .I1 (g650), .I2 (g3343));
AN2X1 gate7327(.O (g10682), .I1 (g10600), .I2 (g3863));
AN2X1 gate7328(.O (g6687), .I1 (g5486), .I2 (g5840));
AN2X1 gate7329(.O (g7704), .I1 (g682), .I2 (g7197));
AN2X1 gate7330(.O (g4582), .I1 (g525), .I2 (g4055));
AN2X1 gate7331(.O (g4261), .I1 (g1019), .I2 (g3914));
AN2X1 gate7332(.O (g3422), .I1 (g225), .I2 (g3228));
AN2X1 gate7333(.O (g5745), .I1 (g1549), .I2 (g5192));
AN2X1 gate7334(.O (g8387), .I1 (g6086), .I2 (g8220));
AN2X1 gate7335(.O (g7954), .I1 (g2874), .I2 (g7512));
AN2X1 gate7336(.O (g11283), .I1 (g4966), .I2 (g11205));
AN2X1 gate7337(.O (g8461), .I1 (g8298), .I2 (g7403));
AN2X1 gate7338(.O (g10760), .I1 (g10695), .I2 (g10691));
AN2X1 gate7339(.O (g11492), .I1 (g11480), .I2 (g4807));
AN3X1 gate7340(.O (g7032), .I1 (g2965), .I2 (g6626), .I3 (g5292));
AN2X1 gate7341(.O (g8756), .I1 (g7431), .I2 (g8674));
AN2X1 gate7342(.O (g9151), .I1 (g8967), .I2 (g6674));
AN2X1 gate7343(.O (g6341), .I1 (g272), .I2 (g5885));
AN2X1 gate7344(.O (g10506), .I1 (g10390), .I2 (g2135));
AN2X1 gate7345(.O (g9648), .I1 (g16), .I2 (g9274));
AN2X1 gate7346(.O (g7453), .I1 (g7148), .I2 (g2809));
AN2X1 gate7347(.O (g6525), .I1 (g5995), .I2 (g3102));
AN2X1 gate7348(.O (g6645), .I1 (g67), .I2 (g6202));
AN2X1 gate7349(.O (g5707), .I1 (g1595), .I2 (g5122));
AN2X1 gate7350(.O (g8046), .I1 (g7548), .I2 (g5128));
AN2X1 gate7351(.O (g11091), .I1 (g833), .I2 (g10950));
AN2X1 gate7352(.O (g11174), .I1 (g496), .I2 (g11112));
AN2X1 gate7353(.O (g9010), .I1 (g6454), .I2 (g8930));
AN2X1 gate7354(.O (g8403), .I1 (g6101), .I2 (g8239));
AN2X1 gate7355(.O (g5201), .I1 (g1250), .I2 (g4721));
AN2X1 gate7356(.O (g8841), .I1 (g8605), .I2 (g8704));
AN2X1 gate7357(.O (g6879), .I1 (g1914), .I2 (g6407));
AN2X1 gate7358(.O (g8763), .I1 (g7440), .I2 (g8680));
AN2X1 gate7359(.O (g4502), .I1 (g2031), .I2 (g3938));
AN2X1 gate7360(.O (g9839), .I1 (g9702), .I2 (g9742));
AN2X1 gate7361(.O (g6358), .I1 (g5841), .I2 (g4441));
AN2X1 gate7362(.O (g5575), .I1 (g1618), .I2 (g4501));
AN2X1 gate7363(.O (g4940), .I1 (g3500), .I2 (g4440));
AN2X1 gate7364(.O (g8107), .I1 (g6226), .I2 (g7882));
AN2X1 gate7365(.O (g10240), .I1 (g10150), .I2 (g9103));
AN2X1 gate7366(.O (g11192), .I1 (g5628), .I2 (g11066));
AN2X1 gate7367(.O (g9618), .I1 (g910), .I2 (g9205));
AN2X1 gate7368(.O (g5539), .I1 (g1684), .I2 (g4314));
AN2X1 gate7369(.O (g8416), .I1 (g731), .I2 (g8151));
AN2X1 gate7370(.O (g9693), .I1 (g275), .I2 (g9432));
AN2X1 gate7371(.O (g11553), .I1 (g2683), .I2 (g11519));
AN2X1 gate7372(.O (g8047), .I1 (g7557), .I2 (g5919));
AN2X1 gate7373(.O (g5268), .I1 (g1098), .I2 (g4769));
AN2X1 gate7374(.O (g9555), .I1 (g9107), .I2 (g3391));
AN2X1 gate7375(.O (g6180), .I1 (g2190), .I2 (g5128));
AN2X1 gate7376(.O (g6832), .I1 (g1383), .I2 (g6596));
AN2X1 gate7377(.O (g10633), .I1 (g10600), .I2 (g3829));
AN2X1 gate7378(.O (g7894), .I1 (g7617), .I2 (g3816));
AN2X1 gate7379(.O (g8654), .I1 (g8529), .I2 (g4013));
AN2X1 gate7380(.O (g9621), .I1 (g1179), .I2 (g9125));
AN2X1 gate7381(.O (g6794), .I1 (g5819), .I2 (g4415));
AN2X1 gate7382(.O (g9313), .I1 (g8876), .I2 (g5708));
AN2X1 gate7383(.O (g4883), .I1 (g248), .I2 (g3946));
AN2X1 gate7384(.O (g3412), .I1 (g219), .I2 (g3228));
AN2X1 gate7385(.O (g7661), .I1 (g7127), .I2 (g2251));
AN3X1 gate7386(.O (g2800), .I1 (g2399), .I2 (g2369), .I3 (g591));
AN2X1 gate7387(.O (g3389), .I1 (g207), .I2 (g3228));
AN2X1 gate7388(.O (g3706), .I1 (g471), .I2 (g3268));
AN2X1 gate7389(.O (g9908), .I1 (g9890), .I2 (g9782));
AN2X1 gate7390(.O (g3429), .I1 (g231), .I2 (g3228));
AN2X1 gate7391(.O (g6628), .I1 (g351), .I2 (g6182));
AN2X1 gate7392(.O (g5470), .I1 (g1044), .I2 (g4222));
AN2X1 gate7393(.O (g7526), .I1 (g7148), .I2 (g2868));
AN2X1 gate7394(.O (g5897), .I1 (g2204), .I2 (g5354));
AN2X1 gate7395(.O (g5025), .I1 (g1482), .I2 (g4640));
AN2X1 gate7396(.O (g6204), .I1 (g3738), .I2 (g4921));
AN2X1 gate7397(.O (g4048), .I1 (g1750), .I2 (g2790));
AN3X1 gate7398(.O (g8935), .I1 (g8106), .I2 (g6778), .I3 (g8849));
AN2X1 gate7399(.O (g3281), .I1 (g766), .I2 (g2525));
AN2X1 gate7400(.O (g9593), .I1 (g898), .I2 (g9205));
AN2X1 gate7401(.O (g4827), .I1 (g213), .I2 (g3946));
AN2X1 gate7402(.O (g10701), .I1 (g10620), .I2 (g10619));
AN2X1 gate7403(.O (g10777), .I1 (g10733), .I2 (g3015));
AN2X1 gate7404(.O (g8130), .I1 (g1936), .I2 (g7952));
AN2X1 gate7405(.O (g9965), .I1 (g9955), .I2 (g9536));
AN2X1 gate7406(.O (g3684), .I1 (g1710), .I2 (g3015));
AN2X1 gate7407(.O (g11213), .I1 (g947), .I2 (g11157));
AN2X1 gate7408(.O (g5006), .I1 (g1462), .I2 (g4640));
AN2X1 gate7409(.O (g9933), .I1 (g9912), .I2 (g9624));
AN2X1 gate7410(.O (g8554), .I1 (g8407), .I2 (g8020));
AN2X1 gate7411(.O (g9641), .I1 (g913), .I2 (g9205));
AN2X1 gate7412(.O (g6123), .I1 (g5630), .I2 (g4311));
AN2X1 gate7413(.O (g6323), .I1 (g1235), .I2 (g5949));
AN2X1 gate7414(.O (g10766), .I1 (g10646), .I2 (g4840));
AN2X1 gate7415(.O (g6666), .I1 (g5301), .I2 (g5818));
AN2X1 gate7416(.O (g4994), .I1 (g1504), .I2 (g4640));
AN2X1 gate7417(.O (g5755), .I1 (g5103), .I2 (g5354));
AN2X1 gate7418(.O (g11592), .I1 (g3717), .I2 (g11561));
AN2X1 gate7419(.O (g6351), .I1 (g6210), .I2 (g5052));
AN2X1 gate7420(.O (g6875), .I1 (g1905), .I2 (g6400));
AN2X1 gate7421(.O (g4816), .I1 (g4070), .I2 (g2336));
AN2X1 gate7422(.O (g9658), .I1 (g947), .I2 (g9240));
AN2X1 gate7423(.O (g6530), .I1 (g6207), .I2 (g3829));
AN2X1 gate7424(.O (g8366), .I1 (g8199), .I2 (g7265));
AN2X1 gate7425(.O (g9835), .I1 (g9735), .I2 (g9785));
AN2X1 gate7426(.O (g6655), .I1 (g5296), .I2 (g5812));
AN3X1 gate7427(.O (g5445), .I1 (g4631), .I2 (g3875), .I3 (g2733));
AN2X1 gate7428(.O (g5173), .I1 (g3094), .I2 (g4676));
AN2X1 gate7429(.O (g7970), .I1 (g7384), .I2 (g7703));
AN2X1 gate7430(.O (g3098), .I1 (g2331), .I2 (g2198));
AN2X1 gate7431(.O (g5491), .I1 (g1624), .I2 (g4262));
AN2X1 gate7432(.O (g9271), .I1 (g6681), .I2 (g8949));
AN2X1 gate7433(.O (g11152), .I1 (g369), .I2 (g10903));
AN2X1 gate7434(.O (g9611), .I1 (g2651), .I2 (g9010));
AN2X1 gate7435(.O (g6410), .I1 (g2804), .I2 (g5759));
AN2X1 gate7436(.O (g10451), .I1 (g10444), .I2 (g3365));
AN2X1 gate7437(.O (g4397), .I1 (g3475), .I2 (g2181));
AN2X1 gate7438(.O (g7224), .I1 (g5398), .I2 (g6441));
AN2X1 gate7439(.O (g5602), .I1 (g1624), .I2 (g4535));
AN2X1 gate7440(.O (g4421), .I1 (g4112), .I2 (g2980));
AN2X1 gate7441(.O (g6884), .I1 (g5569), .I2 (g6564));
AN2X1 gate7442(.O (g6839), .I1 (g1397), .I2 (g6596));
AN2X1 gate7443(.O (g8698), .I1 (g7591), .I2 (g8576));
AN3X1 gate7444(.O (g8964), .I1 (g8255), .I2 (g6368), .I3 (g8849));
AN2X1 gate7445(.O (g8260), .I1 (g2775), .I2 (g7911));
AN2X1 gate7446(.O (g11413), .I1 (g11354), .I2 (g10679));
AN2X1 gate7447(.O (g4950), .I1 (g1415), .I2 (g4682));
AN2X1 gate7448(.O (g5535), .I1 (g4327), .I2 (g3544));
AN2X1 gate7449(.O (g7277), .I1 (g6772), .I2 (g731));
AN2X1 gate7450(.O (g8463), .I1 (g8301), .I2 (g7410));
AN2X1 gate7451(.O (g3268), .I1 (g466), .I2 (g2511));
AN2X1 gate7452(.O (g10785), .I1 (g10728), .I2 (g5177));
AN2X1 gate7453(.O (g6618), .I1 (g658), .I2 (g6016));
AN2X1 gate7454(.O (g6235), .I1 (g569), .I2 (g5089));
AN2X1 gate7455(.O (g10950), .I1 (g10788), .I2 (g6355));
AN2X1 gate7456(.O (g4723), .I1 (g3626), .I2 (g2779));
AN2X1 gate7457(.O (g8720), .I1 (g8601), .I2 (g7905));
AN2X1 gate7458(.O (g6693), .I1 (g5494), .I2 (g5845));
AN2X1 gate7459(.O (g11020), .I1 (g452), .I2 (g10974));
AN2X1 gate7460(.O (g11583), .I1 (g1314), .I2 (g11541));
AN2X1 gate7461(.O (g8118), .I1 (g1900), .I2 (g7941));
AN2X1 gate7462(.O (g8167), .I1 (g5253), .I2 (g7853));
AN2X1 gate7463(.O (g6334), .I1 (g1389), .I2 (g5904));
AN2X1 gate7464(.O (g7892), .I1 (g7616), .I2 (g3815));
AN2X1 gate7465(.O (g8652), .I1 (g8523), .I2 (g4013));
AN2X1 gate7466(.O (g5721), .I1 (g1577), .I2 (g5143));
AN2X1 gate7467(.O (g10367), .I1 (g10362), .I2 (g3375));
AN2X1 gate7468(.O (g9901), .I1 (g9893), .I2 (g9392));
AN2X1 gate7469(.O (g6792), .I1 (g290), .I2 (g5881));
AN2X1 gate7470(.O (g11282), .I1 (g4958), .I2 (g11203));
AN2X1 gate7471(.O (g7945), .I1 (g2847), .I2 (g7473));
AN3X1 gate7472(.O (g8971), .I1 (g8081), .I2 (g6764), .I3 (g8858));
AN2X1 gate7473(.O (g11302), .I1 (g5508), .I2 (g11244));
AN2X1 gate7474(.O (g4585), .I1 (g521), .I2 (g4060));
AN2X1 gate7475(.O (g6621), .I1 (g52), .I2 (g6164));
AN2X1 gate7476(.O (g5502), .I1 (g1932), .I2 (g4275));
AN2X1 gate7477(.O (g11105), .I1 (g3634), .I2 (g10937));
AN2X1 gate7478(.O (g7709), .I1 (g6856), .I2 (g4333));
AN2X1 gate7479(.O (g8598), .I1 (g8471), .I2 (g7432));
AN2X1 gate7480(.O (g7140), .I1 (g6069), .I2 (g6711));
AN2X1 gate7481(.O (g9600), .I1 (g904), .I2 (g9205));
AN2X1 gate7482(.O (g9864), .I1 (g1604), .I2 (g9778));
AN2X1 gate7483(.O (g11640), .I1 (g11613), .I2 (g7900));
AN2X1 gate7484(.O (g5188), .I1 (g4504), .I2 (g4496));
AN2X1 gate7485(.O (g7435), .I1 (g7260), .I2 (g6572));
AN2X1 gate7486(.O (g7876), .I1 (g7609), .I2 (g3790));
AN2X1 gate7487(.O (g5030), .I1 (g1280), .I2 (g4523));
AN2X1 gate7488(.O (g4058), .I1 (g2707), .I2 (g2276));
AN2X1 gate7489(.O (g6776), .I1 (g5809), .I2 (g4390));
AN2X1 gate7490(.O (g4890), .I1 (g630), .I2 (g4739));
AN2X1 gate7491(.O (g2525), .I1 (g762), .I2 (g758));
AN2X1 gate7492(.O (g10301), .I1 (g8892), .I2 (g10223));
AN2X1 gate7493(.O (g4505), .I1 (g354), .I2 (g3586));
AN2X1 gate7494(.O (g9623), .I1 (g17), .I2 (g9274));
AN2X1 gate7495(.O (g10739), .I1 (g10676), .I2 (g3368));
AN2X1 gate7496(.O (g11027), .I1 (g391), .I2 (g10974));
AN2X1 gate7497(.O (g10738), .I1 (g10692), .I2 (g4840));
AN2X1 gate7498(.O (g8687), .I1 (g8558), .I2 (g8036));
AN2X1 gate7499(.O (g6360), .I1 (g302), .I2 (g5899));
AN2X1 gate7500(.O (g9871), .I1 (g1564), .I2 (g9668));
AN2X1 gate7501(.O (g5108), .I1 (g1801), .I2 (g4614));
AN2X1 gate7502(.O (g11248), .I1 (g976), .I2 (g11071));
AN2X1 gate7503(.O (g4992), .I1 (g1407), .I2 (g4682));
AN2X1 gate7504(.O (g11552), .I1 (g2677), .I2 (g11519));
AN2X1 gate7505(.O (g9651), .I1 (g944), .I2 (g9240));
AN2X1 gate7506(.O (g11204), .I1 (g971), .I2 (g11083));
AN2X1 gate7507(.O (g7824), .I1 (g1932), .I2 (g7479));
AN2X1 gate7508(.O (g4480), .I1 (g1133), .I2 (g3905));
AN2X1 gate7509(.O (g6179), .I1 (g5115), .I2 (g5354));
AN2X1 gate7510(.O (g8710), .I1 (g7607), .I2 (g8595));
AN2X1 gate7511(.O (g7590), .I1 (g7102), .I2 (g5425));
AN2X1 gate7512(.O (g9384), .I1 (g968), .I2 (g9223));
AN2X1 gate7513(.O (g3407), .I1 (g2561), .I2 (g3012));
AN2X1 gate7514(.O (g9838), .I1 (g9700), .I2 (g9754));
AN2X1 gate7515(.O (g3718), .I1 (g192), .I2 (g3164));
AN2X1 gate7516(.O (g10661), .I1 (g10594), .I2 (g3015));
AN2X1 gate7517(.O (g11380), .I1 (g11321), .I2 (g4285));
AN3X1 gate7518(.O (g8879), .I1 (g8110), .I2 (g6764), .I3 (g8858));
AN2X1 gate7519(.O (g7930), .I1 (g7621), .I2 (g3110));
AN3X1 gate7520(.O (g8962), .I1 (g8089), .I2 (g6368), .I3 (g8828));
AN2X1 gate7521(.O (g10715), .I1 (g2272), .I2 (g10630));
AN2X1 gate7522(.O (g8659), .I1 (g8535), .I2 (g4013));
AN2X1 gate7523(.O (g3015), .I1 (g2028), .I2 (g2191));
AN2X1 gate7524(.O (g9643), .I1 (g950), .I2 (g9223));
AN2X1 gate7525(.O (g9205), .I1 (g6454), .I2 (g8957));
AN2X1 gate7526(.O (g5538), .I1 (g1669), .I2 (g4313));
AN2X1 gate7527(.O (g4000), .I1 (g1744), .I2 (g2778));
AN2X1 gate7528(.O (g4126), .I1 (g2701), .I2 (g3040));
AN2X1 gate7529(.O (g4400), .I1 (g4088), .I2 (g3829));
AN2X1 gate7530(.O (g2794), .I1 (I5886), .I2 (I5887));
AN2X1 gate7531(.O (g4760), .I1 (g486), .I2 (g3393));
AN2X1 gate7532(.O (g6238), .I1 (g572), .I2 (g5096));
AN2X1 gate7533(.O (g10784), .I1 (g10727), .I2 (g5169));
AN2X1 gate7534(.O (g8174), .I1 (g5284), .I2 (g7853));
AN2X1 gate7535(.O (g6332), .I1 (g1374), .I2 (g5904));
AN2X1 gate7536(.O (g5067), .I1 (g305), .I2 (g4811));
AN2X1 gate7537(.O (g5418), .I1 (g1512), .I2 (g4344));
AN2X1 gate7538(.O (g10297), .I1 (g8892), .I2 (g10211));
AN2X1 gate7539(.O (g6353), .I1 (g299), .I2 (g5895));
AN2X1 gate7540(.O (g11026), .I1 (g386), .I2 (g10974));
AN2X1 gate7541(.O (g11212), .I1 (g944), .I2 (g11155));
AN2X1 gate7542(.O (g6744), .I1 (g4828), .I2 (g6151));
AN2X1 gate7543(.O (g5493), .I1 (g1923), .I2 (g4265));
AN2X1 gate7544(.O (g10671), .I1 (g10578), .I2 (g9431));
AN2X1 gate7545(.O (g4383), .I1 (g2517), .I2 (g3829));
AN2X1 gate7546(.O (g5256), .I1 (g4297), .I2 (g2779));
AN2X1 gate7547(.O (g4220), .I1 (g105), .I2 (g3539));
AN2X1 gate7548(.O (g8380), .I1 (g8252), .I2 (g4240));
AN2X1 gate7549(.O (g7071), .I1 (g5916), .I2 (g6590));
AN2X1 gate7550(.O (g4779), .I1 (g501), .I2 (g3427));
AN2X1 gate7551(.O (g9613), .I1 (g1176), .I2 (g9125));
AN2X1 gate7552(.O (g7705), .I1 (g6853), .I2 (g4328));
AN2X1 gate7553(.O (g9269), .I1 (g8933), .I2 (g3413));
AN2X1 gate7554(.O (g5181), .I1 (g4520), .I2 (g4510));
AN2X1 gate7555(.O (g4977), .I1 (g4567), .I2 (g4807));
AN2X1 gate7556(.O (g7948), .I1 (g2855), .I2 (g7497));
AN2X1 gate7557(.O (g11149), .I1 (g324), .I2 (g10930));
AN2X1 gate7558(.O (g9862), .I1 (g1601), .I2 (g9777));
AN2X1 gate7559(.O (g11387), .I1 (g11284), .I2 (g3629));
AN2X1 gate7560(.O (g7955), .I1 (g2877), .I2 (g7516));
AN2X1 gate7561(.O (g4161), .I1 (g2719), .I2 (g3060));
AN2X1 gate7562(.O (g11148), .I1 (g2321), .I2 (g10913));
AN2X1 gate7563(.O (g9712), .I1 (g1528), .I2 (g9490));
AN2X1 gate7564(.O (g8931), .I1 (g8807), .I2 (g8164));
AN2X1 gate7565(.O (g11097), .I1 (g378), .I2 (g10884));
AN3X1 gate7566(.O (g5421), .I1 (g4631), .I2 (g2733), .I3 (g3819));
AN2X1 gate7567(.O (g11104), .I1 (g2963), .I2 (g10937));
AN2X1 gate7568(.O (g5263), .I1 (g709), .I2 (g4761));
AN2X1 gate7569(.O (g6092), .I1 (g1059), .I2 (g5320));
AN2X1 gate7570(.O (g4999), .I1 (g1499), .I2 (g4640));
AN4X1 gate7571(.O (I6338), .I1 (g2475), .I2 (g2456), .I3 (g2451), .I4 (g2446));
AN3X1 gate7572(.O (g7409), .I1 (g4976), .I2 (g632), .I3 (g6858));
AN2X1 gate7573(.O (g4103), .I1 (g2683), .I2 (g2997));
AN4X1 gate7574(.O (I6309), .I1 (g2446), .I2 (g2451), .I3 (g2456), .I4 (g2475));
AN2X1 gate7575(.O (g6580), .I1 (g1801), .I2 (g5944));
AN2X1 gate7576(.O (g5631), .I1 (g1056), .I2 (g4416));
AN2X1 gate7577(.O (g9414), .I1 (g1730), .I2 (g9052));
AN2X1 gate7578(.O (g9660), .I1 (g1188), .I2 (g9125));
AN2X1 gate7579(.O (g9946), .I1 (g9926), .I2 (g9392));
AN2X1 gate7580(.O (g5257), .I1 (g691), .I2 (g4755));
AN2X1 gate7581(.O (g4732), .I1 (g391), .I2 (g3372));
AN2X1 gate7582(.O (g3108), .I1 (I6330), .I2 (I6331));
AN2X1 gate7583(.O (g4753), .I1 (g481), .I2 (g3386));
AN2X1 gate7584(.O (g9903), .I1 (g9885), .I2 (g9673));
AN2X1 gate7585(.O (g10625), .I1 (g10546), .I2 (g4552));
AN2X1 gate7586(.O (g5605), .I1 (g4828), .I2 (g704));
AN2X1 gate7587(.O (g6623), .I1 (g55), .I2 (g6170));
AN2X1 gate7588(.O (g11228), .I1 (g466), .I2 (g11060));
AN2X1 gate7589(.O (g11011), .I1 (g1968), .I2 (g10809));
AN2X1 gate7590(.O (g6889), .I1 (g1941), .I2 (g6427));
AN2X1 gate7591(.O (g8040), .I1 (g7523), .I2 (g5128));
AN2X1 gate7592(.O (g7822), .I1 (g1914), .I2 (g7479));
AN2X1 gate7593(.O (g8123), .I1 (g1918), .I2 (g7946));
AN2X1 gate7594(.O (g11582), .I1 (g1311), .I2 (g11540));
AN2X1 gate7595(.O (g4316), .I1 (g1965), .I2 (g3400));
AN2X1 gate7596(.O (g10969), .I1 (g3625), .I2 (g10809));
AN2X1 gate7597(.O (g5041), .I1 (g3983), .I2 (g4401));
AN2X1 gate7598(.O (g9335), .I1 (g8975), .I2 (g5708));
AN2X1 gate7599(.O (g9831), .I1 (g9727), .I2 (g9785));
AN2X1 gate7600(.O (g4565), .I1 (g534), .I2 (g4010));
AN2X1 gate7601(.O (g9422), .I1 (g1750), .I2 (g9030));
AN2X1 gate7602(.O (g8648), .I1 (g4588), .I2 (g8511));
AN3X1 gate7603(.O (g8875), .I1 (g8255), .I2 (g6368), .I3 (g8858));
AN2X1 gate7604(.O (g5168), .I1 (g1512), .I2 (g4679));
AN2X1 gate7605(.O (g7895), .I1 (g7503), .I2 (g7036));
AN2X1 gate7606(.O (g8655), .I1 (g8532), .I2 (g4013));
AN2X1 gate7607(.O (g3396), .I1 (g213), .I2 (g3228));
AN2X1 gate7608(.O (g4914), .I1 (g1062), .I2 (g4436));
AN2X1 gate7609(.O (g9947), .I1 (g9927), .I2 (g9392));
AN2X1 gate7610(.O (g5772), .I1 (g1555), .I2 (g5214));
AN2X1 gate7611(.O (g6838), .I1 (g192), .I2 (g6596));
AN2X1 gate7612(.O (g5531), .I1 (g1666), .I2 (g4306));
AN2X1 gate7613(.O (g6795), .I1 (g5036), .I2 (g5878));
AN2X1 gate7614(.O (g10503), .I1 (g10388), .I2 (g2135));
AN2X1 gate7615(.O (g8010), .I1 (g7738), .I2 (g7413));
AN2X1 gate7616(.O (g8410), .I1 (g713), .I2 (g8143));
AN2X1 gate7617(.O (g6231), .I1 (g818), .I2 (g5608));
AN2X1 gate7618(.O (g10581), .I1 (g10531), .I2 (g9453));
AN2X1 gate7619(.O (g10450), .I1 (g10364), .I2 (g3359));
AN2X1 gate7620(.O (g2804), .I1 (g2132), .I2 (g1891));
AN2X1 gate7621(.O (g3418), .I1 (g2379), .I2 (g3012));
AN2X1 gate7622(.O (g4820), .I1 (g186), .I2 (g3946));
AN2X1 gate7623(.O (g9653), .I1 (g1185), .I2 (g9125));
AN2X1 gate7624(.O (g6205), .I1 (g1515), .I2 (g5151));
AN2X1 gate7625(.O (g10818), .I1 (g10730), .I2 (g4545));
AN2X1 gate7626(.O (g8172), .I1 (g5275), .I2 (g7853));
AN2X1 gate7627(.O (g10496), .I1 (g10429), .I2 (g3977));
AN2X1 gate7628(.O (g5074), .I1 (g1771), .I2 (g4587));
AN2X1 gate7629(.O (g9869), .I1 (g1558), .I2 (g9814));
AN2X1 gate7630(.O (g9719), .I1 (g1543), .I2 (g9490));
AN2X1 gate7631(.O (g10741), .I1 (g10635), .I2 (g4013));
AN2X1 gate7632(.O (g3381), .I1 (g940), .I2 (g2756));
AN2X1 gate7633(.O (g5863), .I1 (g5272), .I2 (g2173));
AN2X1 gate7634(.O (g8693), .I1 (g3738), .I2 (g8509));
AN2X1 gate7635(.O (g5480), .I1 (g4279), .I2 (g3519));
AN2X1 gate7636(.O (g4581), .I1 (g3766), .I2 (g3254));
AN2X1 gate7637(.O (g3685), .I1 (g1781), .I2 (g2981));
AN2X1 gate7638(.O (g5569), .I1 (g4816), .I2 (g2338));
AN2X1 gate7639(.O (g8555), .I1 (g8409), .I2 (g8025));
AN2X1 gate7640(.O (g3263), .I1 (g2503), .I2 (g2328));
AN2X1 gate7641(.O (g9364), .I1 (g965), .I2 (g9223));
AN2X1 gate7642(.O (g4784), .I1 (g506), .I2 (g3432));
AN2X1 gate7643(.O (g9454), .I1 (g8994), .I2 (g5708));
AN4X1 gate7644(.O (I6331), .I1 (g2060), .I2 (g2070), .I3 (g2074), .I4 (g2077));
AN2X1 gate7645(.O (g11299), .I1 (g5498), .I2 (g11243));
AN2X1 gate7646(.O (g6983), .I1 (g6592), .I2 (g3105));
AN2X1 gate7647(.O (g7958), .I1 (g736), .I2 (g7697));
AN2X1 gate7648(.O (g4995), .I1 (g1474), .I2 (g4640));
AN2X1 gate7649(.O (g4079), .I1 (g2765), .I2 (g2276));
AN2X1 gate7650(.O (g2264), .I1 (g1771), .I2 (g1766));
AN2X1 gate7651(.O (g2160), .I1 (g745), .I2 (g746));
AN2X1 gate7652(.O (g3257), .I1 (g378), .I2 (g2496));
AN2X1 gate7653(.O (g3101), .I1 (I6309), .I2 (I6310));
AN2X1 gate7654(.O (g5000), .I1 (g1470), .I2 (g4640));
AN2X1 gate7655(.O (g3301), .I1 (g1346), .I2 (g2544));
AN2X1 gate7656(.O (g5126), .I1 (g3076), .I2 (g4638));
AN4X1 gate7657(.O (I5084), .I1 (g1462), .I2 (g1470), .I3 (g1474), .I4 (g1478));
AN2X1 gate7658(.O (g9412), .I1 (g1727), .I2 (g9052));
AN2X1 gate7659(.O (g9389), .I1 (g1330), .I2 (g9151));
AN2X1 gate7660(.O (g2379), .I1 (g744), .I2 (g743));
AN2X1 gate7661(.O (g10706), .I1 (g10567), .I2 (g4840));
AN3X1 gate7662(.O (I16145), .I1 (g10366), .I2 (g10447), .I3 (g10446));
AN2X1 gate7663(.O (g10597), .I1 (g10533), .I2 (g4359));
AN3X1 gate7664(.O (g8965), .I1 (g8110), .I2 (g6778), .I3 (g8849));
AN2X1 gate7665(.O (g5608), .I1 (g814), .I2 (g4831));
AN2X1 gate7666(.O (g5220), .I1 (g1083), .I2 (g4729));
AN2X1 gate7667(.O (g10624), .I1 (g10545), .I2 (g4544));
AN2X1 gate7668(.O (g10300), .I1 (g8892), .I2 (g10220));
AN2X1 gate7669(.O (g5023), .I1 (g1071), .I2 (g4511));
AN2X1 gate7670(.O (g4432), .I1 (g3723), .I2 (g1975));
AN2X1 gate7671(.O (g4053), .I1 (g2701), .I2 (g2276));
AN2X1 gate7672(.O (g8050), .I1 (g7596), .I2 (g5919));
AN2X1 gate7673(.O (g5588), .I1 (g1639), .I2 (g4508));
AN3X1 gate7674(.O (g6679), .I1 (g4631), .I2 (g6074), .I3 (g2733));
AN2X1 gate7675(.O (g9963), .I1 (g9953), .I2 (g9536));
AN2X1 gate7676(.O (g3772), .I1 (g2542), .I2 (g3089));
AN2X1 gate7677(.O (g5051), .I1 (g4432), .I2 (g2834));
AN2X1 gate7678(.O (g6831), .I1 (g207), .I2 (g6596));
AN2X1 gate7679(.O (g2981), .I1 (g1776), .I2 (g2264));
AN2X1 gate7680(.O (g8724), .I1 (g8606), .I2 (g7910));
AN2X1 gate7681(.O (g4157), .I1 (g2713), .I2 (g3055));
AN2X1 gate7682(.O (g9707), .I1 (g1583), .I2 (g9474));
AN3X1 gate7683(.O (g8878), .I1 (g8099), .I2 (g6368), .I3 (g8858));
AN2X1 gate7684(.O (g2132), .I1 (g1872), .I2 (g1882));
AN2X1 gate7685(.O (g10763), .I1 (g10639), .I2 (g4840));
AN3X1 gate7686(.O (g8289), .I1 (g6777), .I2 (g8109), .I3 (g6475));
AN2X1 gate7687(.O (g7898), .I1 (g7511), .I2 (g7041));
AN2X1 gate7688(.O (g11271), .I1 (g5624), .I2 (g11191));
AN2X1 gate7689(.O (g11461), .I1 (g11429), .I2 (g5446));
AN2X1 gate7690(.O (g5732), .I1 (g1604), .I2 (g5176));
AN2X1 gate7691(.O (g11145), .I1 (g315), .I2 (g10927));
AN2X1 gate7692(.O (g11031), .I1 (g411), .I2 (g10974));
AN2X1 gate7693(.O (g9865), .I1 (g1607), .I2 (g9780));
AN2X1 gate7694(.O (g5944), .I1 (g1796), .I2 (g5233));
AN2X1 gate7695(.O (g9715), .I1 (g1531), .I2 (g9490));
AN2X1 gate7696(.O (g9604), .I1 (g1194), .I2 (g9111));
AN2X1 gate7697(.O (g8799), .I1 (g8647), .I2 (g8727));
AN2X1 gate7698(.O (g11198), .I1 (g4919), .I2 (g11069));
AN2X1 gate7699(.O (g6873), .I1 (g3263), .I2 (g6557));
AN2X1 gate7700(.O (g6632), .I1 (g61), .I2 (g6190));
AN2X1 gate7701(.O (g6095), .I1 (g1062), .I2 (g5320));
AN2X1 gate7702(.O (g3863), .I1 (g3323), .I2 (g2728));
AN2X1 gate7703(.O (g9833), .I1 (g9729), .I2 (g9785));
AN2X1 gate7704(.O (g6653), .I1 (g70), .I2 (g6213));
AN2X1 gate7705(.O (g6102), .I1 (g1038), .I2 (g5320));
AN2X1 gate7706(.O (g7819), .I1 (g1887), .I2 (g7479));
AN2X1 gate7707(.O (g11393), .I1 (g11280), .I2 (g7916));
AN2X1 gate7708(.O (g2511), .I1 (g461), .I2 (g456));
AN2X1 gate7709(.O (g7088), .I1 (g2331), .I2 (g6737));
AN2X1 gate7710(.O (g9584), .I1 (g2726), .I2 (g9173));
AN2X1 gate7711(.O (g9896), .I1 (g9883), .I2 (g9624));
AN3X1 gate7712(.O (g8209), .I1 (g4094), .I2 (g3792), .I3 (g7980));
AN2X1 gate7713(.O (g6752), .I1 (g6187), .I2 (g2343));
AN2X1 gate7714(.O (g4778), .I1 (g421), .I2 (g3426));
AN2X1 gate7715(.O (g11161), .I1 (g1969), .I2 (g10937));
AN2X1 gate7716(.O (g9268), .I1 (g6681), .I2 (g8947));
AN2X1 gate7717(.O (g5681), .I1 (g135), .I2 (g5361));
AN2X1 gate7718(.O (g7951), .I1 (g2868), .I2 (g7505));
AN2X1 gate7719(.O (g9419), .I1 (g1744), .I2 (g9030));
AN2X1 gate7720(.O (g10268), .I1 (g10183), .I2 (g3307));
AN2X1 gate7721(.O (g5533), .I1 (g1724), .I2 (g4308));
AN2X1 gate7722(.O (g9052), .I1 (g8936), .I2 (g7192));
AN2X1 gate7723(.O (g6786), .I1 (g178), .I2 (g5919));
AN2X1 gate7724(.O (g10670), .I1 (g10571), .I2 (g9091));
AN2X1 gate7725(.O (g11087), .I1 (g829), .I2 (g10950));
AN2X1 gate7726(.O (g4949), .I1 (g3505), .I2 (g4449));
AN2X1 gate7727(.O (g6364), .I1 (g5851), .I2 (g4454));
AN2X1 gate7728(.O (g7825), .I1 (g1941), .I2 (g7479));
AN2X1 gate7729(.O (g3400), .I1 (g115), .I2 (g3164));
AN2X1 gate7730(.O (g4998), .I1 (g1304), .I2 (g4485));
AN2X1 gate7731(.O (g10667), .I1 (g10576), .I2 (g9427));
AN2X1 gate7732(.O (g7136), .I1 (g6050), .I2 (g6704));
AN2X1 gate7733(.O (g6532), .I1 (g339), .I2 (g6057));
AN2X1 gate7734(.O (g9385), .I1 (g1324), .I2 (g9151));
AN4X1 gate7735(.O (I5690), .I1 (g1436), .I2 (g1440), .I3 (g1444), .I4 (g1448));
AN2X1 gate7736(.O (g4484), .I1 (g1137), .I2 (g3909));
AN2X1 gate7737(.O (g9897), .I1 (g9884), .I2 (g9624));
AN2X1 gate7738(.O (g9425), .I1 (g1753), .I2 (g9030));
AN2X1 gate7739(.O (g3383), .I1 (g186), .I2 (g3228));
AN2X1 gate7740(.O (g5601), .I1 (g1035), .I2 (g4375));
AN2X1 gate7741(.O (g7943), .I1 (g2840), .I2 (g7467));
AN2X1 gate7742(.O (g11171), .I1 (g481), .I2 (g11112));
AN2X1 gate7743(.O (g3423), .I1 (I6630), .I2 (I6631));
AN2X1 gate7744(.O (g7230), .I1 (g6064), .I2 (g6444));
AN2X1 gate7745(.O (g4952), .I1 (g1648), .I2 (g4457));
AN2X1 gate7746(.O (g8736), .I1 (g7439), .I2 (g8635));
AN2X1 gate7747(.O (g6787), .I1 (g266), .I2 (g5875));
AN3X1 gate7748(.O (g8968), .I1 (g8089), .I2 (g6778), .I3 (g8849));
AN2X1 gate7749(.O (g10306), .I1 (g10214), .I2 (g9082));
AN2X1 gate7750(.O (g9331), .I1 (g8972), .I2 (g5708));
AN2X1 gate7751(.O (g11459), .I1 (g11427), .I2 (g5446));
AN2X1 gate7752(.O (g4561), .I1 (g538), .I2 (g4003));
AN2X1 gate7753(.O (g11425), .I1 (g11350), .I2 (g10899));
AN2X1 gate7754(.O (g11458), .I1 (g11426), .I2 (g5446));
AN2X1 gate7755(.O (g5739), .I1 (g1607), .I2 (g5185));
AN2X1 gate7756(.O (g7496), .I1 (g7148), .I2 (g2840));
AN2X1 gate7757(.O (g4986), .I1 (g1411), .I2 (g4682));
AN2X1 gate7758(.O (g11010), .I1 (g5187), .I2 (g10827));
AN2X1 gate7759(.O (g3999), .I1 (g1741), .I2 (g2777));
AN2X1 gate7760(.O (g8175), .I1 (g5291), .I2 (g7853));
AN2X1 gate7761(.O (g8722), .I1 (g8604), .I2 (g7908));
AN2X1 gate7762(.O (g4764), .I1 (g411), .I2 (g3404));
AN2X1 gate7763(.O (g7137), .I1 (g5590), .I2 (g6361));
AN2X1 gate7764(.O (g7891), .I1 (g7471), .I2 (g7028));
AN2X1 gate7765(.O (g8651), .I1 (g8520), .I2 (g4013));
AN2X1 gate7766(.O (g5479), .I1 (g1845), .I2 (g4243));
AN2X1 gate7767(.O (g11599), .I1 (g1341), .I2 (g11572));
AN2X1 gate7768(.O (g6684), .I1 (g5314), .I2 (g5836));
AN2X1 gate7769(.O (g6745), .I1 (g5605), .I2 (g6158));
AN2X1 gate7770(.O (g6639), .I1 (g357), .I2 (g6196));
AN2X1 gate7771(.O (g10937), .I1 (g4822), .I2 (g10822));
AN2X1 gate7772(.O (g3696), .I1 (g1713), .I2 (g3015));
AN2X1 gate7773(.O (g4503), .I1 (g654), .I2 (g3943));
AN2X1 gate7774(.O (g6791), .I1 (g269), .I2 (g5880));
AN2X1 gate7775(.O (g5190), .I1 (g1245), .I2 (g4716));
AN2X1 gate7776(.O (g5390), .I1 (g3220), .I2 (g4819));
AN2X1 gate7777(.O (g8384), .I1 (g8180), .I2 (g3397));
AN2X1 gate7778(.O (g4224), .I1 (g1092), .I2 (g3638));
AN2X1 gate7779(.O (g5501), .I1 (g1672), .I2 (g4273));
AN2X1 gate7780(.O (g9173), .I1 (g8968), .I2 (g6674));
AN2X1 gate7781(.O (g6759), .I1 (g148), .I2 (g5919));
AN2X1 gate7782(.O (g8838), .I1 (g8602), .I2 (g8702));
AN2X1 gate7783(.O (g8024), .I1 (g7394), .I2 (g4337));
AN2X1 gate7784(.O (g10666), .I1 (g10575), .I2 (g9424));
AN2X1 gate7785(.O (g11158), .I1 (g309), .I2 (g10935));
AN2X1 gate7786(.O (g9602), .I1 (g2650), .I2 (g9010));
AN2X1 gate7787(.O (g5704), .I1 (g143), .I2 (g5361));
AN2X1 gate7788(.O (g4617), .I1 (g3275), .I2 (g3879));
AN2X1 gate7789(.O (g11561), .I1 (g11518), .I2 (g3015));
AN2X1 gate7790(.O (g9868), .I1 (g1555), .I2 (g9812));
AN2X1 gate7791(.O (g11295), .I1 (g5475), .I2 (g11239));
AN2X1 gate7792(.O (g11144), .I1 (g305), .I2 (g10926));
AN2X1 gate7793(.O (g9718), .I1 (g1540), .I2 (g9490));
AN2X1 gate7794(.O (g3434), .I1 (g237), .I2 (g3228));
AN2X1 gate7795(.O (g4987), .I1 (g1440), .I2 (g4682));
AN2X1 gate7796(.O (g4771), .I1 (g496), .I2 (g3416));
AN2X1 gate7797(.O (g5250), .I1 (g1270), .I2 (g4748));
AN2X1 gate7798(.O (g6098), .I1 (g1065), .I2 (g5320));
AN2X1 gate7799(.O (g9582), .I1 (g2725), .I2 (g9173));
AN2X1 gate7800(.O (g6833), .I1 (g186), .I2 (g6596));
AN2X1 gate7801(.O (g3533), .I1 (g1981), .I2 (g2892));
AN2X1 gate7802(.O (g4892), .I1 (g632), .I2 (g4739));
AN2X1 gate7803(.O (g8104), .I1 (g6218), .I2 (g7880));
AN2X1 gate7804(.O (g9415), .I1 (g1733), .I2 (g9052));
AN2X1 gate7805(.O (g8499), .I1 (g8377), .I2 (g4737));
AN2X1 gate7806(.O (g9664), .I1 (g1191), .I2 (g9125));
AN2X1 gate7807(.O (g10740), .I1 (g10676), .I2 (g3384));
AN2X1 gate7808(.O (g2534), .I1 (g798), .I2 (g794));
AN2X1 gate7809(.O (g8754), .I1 (g7420), .I2 (g8667));
AN2X1 gate7810(.O (g9721), .I1 (g9413), .I2 (g4785));
AN2X1 gate7811(.O (g6162), .I1 (g3584), .I2 (g5200));
AN2X1 gate7812(.O (g4991), .I1 (g1508), .I2 (g4640));
AN2X1 gate7813(.O (g6362), .I1 (g5846), .I2 (g4450));
AN4X1 gate7814(.O (I6631), .I1 (g2707), .I2 (g2713), .I3 (g2719), .I4 (g2765));
AN2X1 gate7815(.O (g10685), .I1 (g10608), .I2 (g3863));
AN2X1 gate7816(.O (g4340), .I1 (g1153), .I2 (g3715));
AN2X1 gate7817(.O (g11023), .I1 (g440), .I2 (g10974));
AN2X1 gate7818(.O (g8044), .I1 (g7598), .I2 (g5919));
AN2X1 gate7819(.O (g11224), .I1 (g968), .I2 (g11056));
AN2X1 gate7820(.O (g11571), .I1 (g2018), .I2 (g11561));
AN2X1 gate7821(.O (g4959), .I1 (g1520), .I2 (g4682));
AN2X1 gate7822(.O (g10334), .I1 (g10265), .I2 (g3307));
AN2X1 gate7823(.O (g5626), .I1 (g1633), .I2 (g4557));
AN2X1 gate7824(.O (g9940), .I1 (g9920), .I2 (g9367));
AN2X1 gate7825(.O (g4876), .I1 (g1086), .I2 (g3638));
AN2X1 gate7826(.O (g6728), .I1 (g6250), .I2 (g4318));
AN2X1 gate7827(.O (g6730), .I1 (g1872), .I2 (g6128));
AN2X1 gate7828(.O (g9689), .I1 (g263), .I2 (g9432));
AN2X1 gate7829(.O (g10762), .I1 (g10635), .I2 (g4840));
AN2X1 gate7830(.O (g6070), .I1 (g1050), .I2 (g5320));
AN2X1 gate7831(.O (g9428), .I1 (g1756), .I2 (g9030));
AN2X1 gate7832(.O (g9030), .I1 (g8935), .I2 (g7192));
AN2X1 gate7833(.O (g9430), .I1 (g1759), .I2 (g9030));
AN2X1 gate7834(.O (g8927), .I1 (g7872), .I2 (g8807));
AN2X1 gate7835(.O (g7068), .I1 (g5912), .I2 (g6586));
AN2X1 gate7836(.O (g8014), .I1 (g7740), .I2 (g7419));
AN2X1 gate7837(.O (g11392), .I1 (g11278), .I2 (g7914));
AN2X1 gate7838(.O (g5782), .I1 (g1558), .I2 (g5223));
AN2X1 gate7839(.O (g9910), .I1 (g9892), .I2 (g9809));
AN2X1 gate7840(.O (g4824), .I1 (g774), .I2 (g4099));
AN2X1 gate7841(.O (g6331), .I1 (g201), .I2 (g5904));
AN2X1 gate7842(.O (g4236), .I1 (g1098), .I2 (g3638));
AN2X1 gate7843(.O (g11559), .I1 (g2719), .I2 (g11519));
AN2X1 gate7844(.O (g9609), .I1 (g907), .I2 (g9205));
AN2X1 gate7845(.O (g11558), .I1 (g2713), .I2 (g11519));
AN2X1 gate7846(.O (g6087), .I1 (g1056), .I2 (g5320));
AN2X1 gate7847(.O (g4877), .I1 (g243), .I2 (g3946));
AN2X1 gate7848(.O (g5526), .I1 (g1950), .I2 (g4294));
AN2X1 gate7849(.O (g10751), .I1 (g10646), .I2 (g4013));
AN2X1 gate7850(.O (g10772), .I1 (g10655), .I2 (g4840));
AN2X1 gate7851(.O (g8135), .I1 (g1945), .I2 (g7956));
AN2X1 gate7852(.O (g11544), .I1 (g11515), .I2 (g10584));
AN2X1 gate7853(.O (g5084), .I1 (g1776), .I2 (g4591));
AN2X1 gate7854(.O (g8382), .I1 (g6077), .I2 (g8213));
AN2X1 gate7855(.O (g10230), .I1 (g8892), .I2 (g10145));
AN2X1 gate7856(.O (g5484), .I1 (g1896), .I2 (g4256));
AN2X1 gate7857(.O (g7241), .I1 (g6772), .I2 (g6172));
AN2X1 gate7858(.O (g3942), .I1 (g219), .I2 (g3164));
AN2X1 gate7859(.O (g10638), .I1 (g10608), .I2 (g3829));
AN2X1 gate7860(.O (g4064), .I1 (g1759), .I2 (g2799));
AN2X1 gate7861(.O (g9365), .I1 (g1321), .I2 (g9151));
AN2X1 gate7862(.O (g9861), .I1 (g9738), .I2 (g9579));
AN2X1 gate7863(.O (g8749), .I1 (g7604), .I2 (g8660));
AN2X1 gate7864(.O (g11255), .I1 (g456), .I2 (g11075));
AN2X1 gate7865(.O (g11189), .I1 (g5616), .I2 (g11064));
AN2X1 gate7866(.O (g10510), .I1 (g10393), .I2 (g2135));
AN3X1 gate7867(.O (g8947), .I1 (g8056), .I2 (g6368), .I3 (g8828));
AN2X1 gate7868(.O (g2917), .I1 (g2424), .I2 (g1657));
AN2X1 gate7869(.O (g5919), .I1 (g5216), .I2 (g2965));
AN2X1 gate7870(.O (g11188), .I1 (g5604), .I2 (g11063));
AN2X1 gate7871(.O (g9846), .I1 (g287), .I2 (g9764));
AN2X1 gate7872(.O (g7818), .I1 (g1878), .I2 (g7479));
AN2X1 gate7873(.O (g11460), .I1 (g11428), .I2 (g5446));
AN2X1 gate7874(.O (g5276), .I1 (g736), .I2 (g4780));
AN2X1 gate7875(.O (g11030), .I1 (g406), .I2 (g10974));
AN2X1 gate7876(.O (g11093), .I1 (g841), .I2 (g10950));
AN2X1 gate7877(.O (g7893), .I1 (g7478), .I2 (g7031));
AN2X1 gate7878(.O (g8653), .I1 (g8526), .I2 (g4013));
AN2X1 gate7879(.O (g10442), .I1 (g10311), .I2 (g2135));
AN2X1 gate7880(.O (g6535), .I1 (g345), .I2 (g6063));
AN2X1 gate7881(.O (g8102), .I1 (g6209), .I2 (g7878));
AN4X1 gate7882(.O (I5085), .I1 (g1490), .I2 (g1494), .I3 (g1504), .I4 (g1508));
AN2X1 gate7883(.O (g5004), .I1 (g1296), .I2 (g4499));
AN2X1 gate7884(.O (g3912), .I1 (g207), .I2 (g3164));
AN2X1 gate7885(.O (g7186), .I1 (g2503), .I2 (g6403));
AN2X1 gate7886(.O (g4489), .I1 (g348), .I2 (g3586));
AN2X1 gate7887(.O (g9662), .I1 (g2094), .I2 (g9292));
AN2X1 gate7888(.O (g9418), .I1 (g1741), .I2 (g9052));
AN2X1 gate7889(.O (g11218), .I1 (g959), .I2 (g11053));
AN2X1 gate7890(.O (g4471), .I1 (g1121), .I2 (g3862));
AN2X1 gate7891(.O (g10746), .I1 (g10643), .I2 (g4013));
AN2X1 gate7892(.O (g7125), .I1 (g1212), .I2 (g6648));
AN2X1 gate7893(.O (g7821), .I1 (g1905), .I2 (g7479));
AN2X1 gate7894(.O (g6246), .I1 (g178), .I2 (g5361));
AN2X1 gate7895(.O (g9256), .I1 (g6689), .I2 (g8963));
AN2X1 gate7896(.O (g8042), .I1 (g7533), .I2 (g5128));
AN2X1 gate7897(.O (g10237), .I1 (g10145), .I2 (g9100));
AN2X1 gate7898(.O (g7939), .I1 (g2829), .I2 (g7460));
AN2X1 gate7899(.O (g8786), .I1 (g8638), .I2 (g8716));
AN2X1 gate7900(.O (g10684), .I1 (g10604), .I2 (g3863));
AN2X1 gate7901(.O (g11455), .I1 (g11435), .I2 (g5446));
AN2X1 gate7902(.O (g8364), .I1 (g658), .I2 (g8235));
AN3X1 gate7903(.O (g2990), .I1 (g2061), .I2 (g2557), .I3 (g1814));
AN2X1 gate7904(.O (g9847), .I1 (g290), .I2 (g9766));
AN2X1 gate7905(.O (g8054), .I1 (g7584), .I2 (g5919));
AN2X1 gate7906(.O (g5617), .I1 (g1050), .I2 (g4391));
AN2X1 gate7907(.O (g6502), .I1 (g5981), .I2 (g3095));
AN2X1 gate7908(.O (g5789), .I1 (g1561), .I2 (g5232));
AN2X1 gate7909(.O (g4009), .I1 (g1747), .I2 (g2789));
AN2X1 gate7910(.O (g11277), .I1 (g4920), .I2 (g11199));
AN2X1 gate7911(.O (g6940), .I1 (g6472), .I2 (g1945));
AN2X1 gate7912(.O (g7061), .I1 (g790), .I2 (g6760));
AN2X1 gate7913(.O (g11595), .I1 (g1336), .I2 (g11575));
AN2X1 gate7914(.O (g5771), .I1 (g1534), .I2 (g5213));
AN2X1 gate7915(.O (g8553), .I1 (g8405), .I2 (g8015));
AN2X1 gate7916(.O (g4836), .I1 (g643), .I2 (g3520));
AN2X1 gate7917(.O (g5547), .I1 (g1733), .I2 (g4326));
AN2X1 gate7918(.O (g6216), .I1 (g2232), .I2 (g5151));
AN2X1 gate7919(.O (g4967), .I1 (g1515), .I2 (g4682));
AN2X1 gate7920(.O (g6671), .I1 (g342), .I2 (g6227));
AN2X1 gate7921(.O (g7200), .I1 (g3098), .I2 (g6418));
AN2X1 gate7922(.O (g3661), .I1 (g382), .I2 (g3257));
AN2X1 gate7923(.O (g7046), .I1 (g5892), .I2 (g6570));
AN2X1 gate7924(.O (g4229), .I1 (g999), .I2 (g3914));
AN2X1 gate7925(.O (g8389), .I1 (g6091), .I2 (g8225));
AN2X1 gate7926(.O (g6430), .I1 (g5044), .I2 (g5791));
AN2X1 gate7927(.O (g8706), .I1 (g7602), .I2 (g8589));
AN2X1 gate7928(.O (g4993), .I1 (g1448), .I2 (g4682));
AN2X1 gate7929(.O (g6247), .I1 (g127), .I2 (g5361));
AN2X1 gate7930(.O (g9257), .I1 (g6689), .I2 (g8964));
AN2X1 gate7931(.O (g11170), .I1 (g525), .I2 (g11112));
AN2X1 gate7932(.O (g7145), .I1 (g6082), .I2 (g6718));
AN2X1 gate7933(.O (g5738), .I1 (g1586), .I2 (g5184));
AN2X1 gate7934(.O (g6826), .I1 (g225), .I2 (g6596));
AN2X1 gate7935(.O (g7191), .I1 (g6343), .I2 (g4323));
AN2X1 gate7936(.O (g3998), .I1 (g2677), .I2 (g2276));
AN2X1 gate7937(.O (g6741), .I1 (g3284), .I2 (g6141));
AN2X1 gate7938(.O (g5478), .I1 (g1905), .I2 (g4242));
AN2X1 gate7939(.O (g11167), .I1 (g538), .I2 (g11112));
AN2X1 gate7940(.O (g11194), .I1 (g5637), .I2 (g11067));
AN2X1 gate7941(.O (g11589), .I1 (g1333), .I2 (g11548));
AN2X1 gate7942(.O (g6638), .I1 (g64), .I2 (g6195));
AN2X1 gate7943(.O (g4921), .I1 (g2779), .I2 (g4431));
AN2X1 gate7944(.O (g7536), .I1 (g7148), .I2 (g2877));
AN2X1 gate7945(.O (g9585), .I1 (g889), .I2 (g8995));
AN2X1 gate7946(.O (g2957), .I1 (g2424), .I2 (g1663));
AN2X1 gate7947(.O (g11588), .I1 (g1330), .I2 (g11547));
AN2X1 gate7948(.O (g5690), .I1 (g1567), .I2 (g5112));
AN2X1 gate7949(.O (g6883), .I1 (g1923), .I2 (g6413));
AN2X1 gate7950(.O (g4837), .I1 (g1068), .I2 (g3638));
AN3X1 gate7951(.O (g8963), .I1 (g8056), .I2 (g6368), .I3 (g8849));
AN2X1 gate7952(.O (g8791), .I1 (g8641), .I2 (g8721));
AN2X1 gate7953(.O (g6217), .I1 (g563), .I2 (g5073));
AN4X1 gate7954(.O (I6316), .I1 (g2082), .I2 (g2087), .I3 (g2381), .I4 (g2395));
AN2X1 gate7955(.O (g11022), .I1 (g444), .I2 (g10974));
AN2X1 gate7956(.O (g5915), .I1 (g4168), .I2 (g4977));
AN2X1 gate7957(.O (g4788), .I1 (g511), .I2 (g3436));
AN2X1 gate7958(.O (g8759), .I1 (g7437), .I2 (g8677));
AN2X1 gate7959(.O (g5110), .I1 (g1806), .I2 (g4618));
AN2X1 gate7960(.O (g11254), .I1 (g986), .I2 (g11073));
AN2X1 gate7961(.O (g6827), .I1 (g219), .I2 (g6596));
AN3X1 gate7962(.O (g8957), .I1 (g8081), .I2 (g6368), .I3 (g8828));
AN2X1 gate7963(.O (g6333), .I1 (g197), .I2 (g5904));
AN2X1 gate7964(.O (g8049), .I1 (g7567), .I2 (g5919));
AN2X1 gate7965(.O (g4392), .I1 (g3273), .I2 (g3829));
AN2X1 gate7966(.O (g9856), .I1 (g1592), .I2 (g9773));
AN2X1 gate7967(.O (g9411), .I1 (g1724), .I2 (g9052));
AN2X1 gate7968(.O (g5002), .I1 (g1494), .I2 (g4640));
AN2X1 gate7969(.O (g11101), .I1 (g857), .I2 (g10950));
AN2X1 gate7970(.O (g11177), .I1 (g511), .I2 (g11112));
AN2X1 gate7971(.O (g11560), .I1 (g2765), .I2 (g11519));
AN2X1 gate7972(.O (g8098), .I1 (g6201), .I2 (g7852));
AN2X1 gate7973(.O (g3970), .I1 (g225), .I2 (g3164));
AN2X1 gate7974(.O (g4941), .I1 (g1038), .I2 (g4451));
AN2X1 gate7975(.O (g10453), .I1 (g10437), .I2 (g3395));
AN2X1 gate7976(.O (g5877), .I1 (g4921), .I2 (g639));
AN2X1 gate7977(.O (g6662), .I1 (g366), .I2 (g6220));
AN2X1 gate7978(.O (g7935), .I1 (g2821), .I2 (g7454));
AN2X1 gate7979(.O (g6067), .I1 (g1047), .I2 (g5320));
AN4X1 gate7980(.O (I6317), .I1 (g2406), .I2 (g2420), .I3 (g2434), .I4 (g2438));
AN2X1 gate7981(.O (g9863), .I1 (g9740), .I2 (g9576));
AN4X1 gate7982(.O (I5886), .I1 (g174), .I2 (g170), .I3 (g2249), .I4 (g2254));
AN2X1 gate7983(.O (g6994), .I1 (g6758), .I2 (g3829));
AN2X1 gate7984(.O (g9713), .I1 (g1589), .I2 (g9474));
AN2X1 gate7985(.O (g4431), .I1 (g2268), .I2 (g3533));
AN2X1 gate7986(.O (g4252), .I1 (g1007), .I2 (g3914));
AN2X1 gate7987(.O (g11166), .I1 (g542), .I2 (g11112));
AN2X1 gate7988(.O (g7130), .I1 (g6041), .I2 (g6697));
AN2X1 gate7989(.O (g11009), .I1 (g5179), .I2 (g10827));
AN2X1 gate7990(.O (g7542), .I1 (g7148), .I2 (g2885));
AN2X1 gate7991(.O (g8019), .I1 (g7386), .I2 (g4332));
AN2X1 gate7992(.O (g11008), .I1 (g5171), .I2 (g10827));
AN2X1 gate7993(.O (g3516), .I1 (g1209), .I2 (g3015));
AN2X1 gate7994(.O (g8052), .I1 (g7573), .I2 (g5128));
AN2X1 gate7995(.O (g3987), .I1 (g243), .I2 (g3164));
AN2X1 gate7996(.O (g4765), .I1 (g491), .I2 (g3405));
AN2X1 gate7997(.O (g11555), .I1 (g2695), .I2 (g11519));
AN2X1 gate7998(.O (g9857), .I1 (g9734), .I2 (g9569));
AN2X1 gate7999(.O (g8728), .I1 (g8610), .I2 (g7915));
AN2X1 gate8000(.O (g8730), .I1 (g8613), .I2 (g7917));
AN2X1 gate8001(.O (g8185), .I1 (g664), .I2 (g7997));
AN2X1 gate8002(.O (g5194), .I1 (g1610), .I2 (g4717));
AN2X1 gate8003(.O (g8385), .I1 (g6084), .I2 (g8218));
AN2X1 gate8004(.O (g4610), .I1 (g3804), .I2 (g2212));
AN2X1 gate8005(.O (g7902), .I1 (g7661), .I2 (g6587));
AN2X1 gate8006(.O (g4073), .I1 (g3200), .I2 (g3222));
AN2X1 gate8007(.O (g8070), .I1 (g682), .I2 (g7826));
AN2X1 gate8008(.O (g5731), .I1 (g1583), .I2 (g5175));
AN2X1 gate8009(.O (g11238), .I1 (g5474), .I2 (g11110));
AN2X1 gate8010(.O (g4473), .I1 (g1125), .I2 (g3874));
AN2X1 gate8011(.O (g8470), .I1 (g8308), .I2 (g7427));
AN2X1 gate8012(.O (g5489), .I1 (g4287), .I2 (g3521));
AN2X1 gate8013(.O (g3991), .I1 (g1738), .I2 (g2774));
AN4X1 gate8014(.O (I5887), .I1 (g2078), .I2 (g2083), .I3 (g166), .I4 (g2095));
AN2X1 gate8015(.O (g7823), .I1 (g1923), .I2 (g7479));
AN2X1 gate8016(.O (g4069), .I1 (g1762), .I2 (g2802));
AN3X1 gate8017(.O (g11519), .I1 (g1317), .I2 (g3015), .I3 (g11492));
AN2X1 gate8018(.O (g11176), .I1 (g506), .I2 (g11112));
AN2X1 gate8019(.O (g11092), .I1 (g837), .I2 (g10950));
AN2X1 gate8020(.O (g11154), .I1 (g330), .I2 (g10932));
AN2X1 gate8021(.O (g9608), .I1 (g7), .I2 (g9292));
AN2X1 gate8022(.O (g11637), .I1 (g11626), .I2 (g5446));
AN2X1 gate8023(.O (g2091), .I1 (g976), .I2 (g971));
AN2X1 gate8024(.O (g8406), .I1 (g695), .I2 (g8131));
AN2X1 gate8025(.O (g5254), .I1 (g4335), .I2 (g4165));
AN2X1 gate8026(.O (g7260), .I1 (g6752), .I2 (g2345));
AN2X1 gate8027(.O (g5150), .I1 (g1275), .I2 (g4678));
AN2X1 gate8028(.O (g8766), .I1 (g8612), .I2 (g5151));
AN2X1 gate8029(.O (g9588), .I1 (g3272), .I2 (g9173));
AN2X1 gate8030(.O (g8801), .I1 (g8742), .I2 (g8729));
AN2X1 gate8031(.O (g7063), .I1 (g5903), .I2 (g6582));
AN2X1 gate8032(.O (g10303), .I1 (g10208), .I2 (g9076));
AN2X1 gate8033(.O (g5009), .I1 (g1486), .I2 (g4640));
AN2X1 gate8034(.O (g9665), .I1 (g1314), .I2 (g9151));
AN2X1 gate8035(.O (g8748), .I1 (g7670), .I2 (g8656));
AN2X1 gate8036(.O (g11215), .I1 (g953), .I2 (g11160));
AN2X1 gate8037(.O (g10750), .I1 (g10687), .I2 (g3586));
AN3X1 gate8038(.O (g5769), .I1 (g2112), .I2 (g4921), .I3 (g3818));
AN2X1 gate8039(.O (g8755), .I1 (g7426), .I2 (g8671));
AN2X1 gate8040(.O (g6673), .I1 (g5305), .I2 (g5822));
AN2X1 gate8041(.O (g5212), .I1 (g1255), .I2 (g4726));
AN2X1 gate8042(.O (g7720), .I1 (g727), .I2 (g7232));
AN3X1 gate8043(.O (g5918), .I1 (g2965), .I2 (g5292), .I3 (g4609));
AN2X1 gate8044(.O (g8045), .I1 (g7547), .I2 (g5128));
AN2X1 gate8045(.O (g8173), .I1 (g7971), .I2 (g3112));
AN2X1 gate8046(.O (g11349), .I1 (g11288), .I2 (g7964));
AN2X1 gate8047(.O (g7843), .I1 (g7599), .I2 (g5919));
AN2X1 gate8048(.O (g9696), .I1 (g281), .I2 (g9432));
AN2X1 gate8049(.O (g6772), .I1 (g6228), .I2 (g722));
AN2X1 gate8050(.O (g6058), .I1 (g1035), .I2 (g5320));
AN2X1 gate8051(.O (g6531), .I1 (g79), .I2 (g6056));
AN2X1 gate8052(.O (g6743), .I1 (g4106), .I2 (g6146));
AN2X1 gate8053(.O (g6890), .I1 (g6752), .I2 (g6568));
AN2X1 gate8054(.O (g7549), .I1 (g7269), .I2 (g3829));
AN2X1 gate8055(.O (g8169), .I1 (g5265), .I2 (g7853));
AN2X1 gate8056(.O (g11304), .I1 (g5520), .I2 (g11245));
AN2X1 gate8057(.O (g9944), .I1 (g9924), .I2 (g9392));
AN2X1 gate8058(.O (g9240), .I1 (g6454), .I2 (g8962));
AN2X1 gate8059(.O (g8059), .I1 (g7592), .I2 (g5919));
AN2X1 gate8060(.O (g8718), .I1 (g8600), .I2 (g7903));
AN2X1 gate8061(.O (g8767), .I1 (g8616), .I2 (g5151));
AN2X1 gate8062(.O (g9316), .I1 (g8877), .I2 (g5708));
AN2X1 gate8063(.O (g7625), .I1 (g673), .I2 (g7085));
AN2X1 gate8064(.O (g8793), .I1 (g8644), .I2 (g8723));
AN2X1 gate8065(.O (g2940), .I1 (g2424), .I2 (g1654));
AN2X1 gate8066(.O (g4114), .I1 (g1351), .I2 (g3301));
AN2X1 gate8067(.O (g11636), .I1 (g11624), .I2 (g7936));
AN2X1 gate8068(.O (g10949), .I1 (g2947), .I2 (g10809));
AN2X1 gate8069(.O (g4870), .I1 (g237), .I2 (g3946));
AN2X1 gate8070(.O (g3563), .I1 (g3275), .I2 (g2126));
AN2X1 gate8071(.O (g10948), .I1 (g2223), .I2 (g10809));
AN2X1 gate8072(.O (g8246), .I1 (g7846), .I2 (g7442));
AN2X1 gate8073(.O (g5788), .I1 (g1540), .I2 (g5231));
AN2X1 gate8074(.O (g4008), .I1 (g2689), .I2 (g2276));
AN2X1 gate8075(.O (g9596), .I1 (g2649), .I2 (g9010));
AN2X1 gate8076(.O (g5249), .I1 (g1089), .I2 (g4747));
AN2X1 gate8077(.O (g11585), .I1 (g1321), .I2 (g11543));
AN2X1 gate8078(.O (g3089), .I1 (g2054), .I2 (g2050));
AN2X1 gate8079(.O (g4972), .I1 (g1436), .I2 (g4682));
AN2X1 gate8080(.O (g11554), .I1 (g2689), .I2 (g11519));
AN2X1 gate8081(.O (g7586), .I1 (g7096), .I2 (g5423));
AN2X1 gate8082(.O (g10673), .I1 (g10580), .I2 (g9450));
AN3X1 gate8083(.O (g4806), .I1 (g3215), .I2 (g3992), .I3 (g2493));
AN2X1 gate8084(.O (g5485), .I1 (g1914), .I2 (g4257));
AN2X1 gate8085(.O (g9936), .I1 (g9915), .I2 (g9624));
AN2X1 gate8086(.O (g2910), .I1 (g2424), .I2 (g1660));
AN2X1 gate8087(.O (g9317), .I1 (g6109), .I2 (g8875));
AN2X1 gate8088(.O (g10933), .I1 (g10853), .I2 (g3982));
AN2X1 gate8089(.O (g8388), .I1 (g8177), .I2 (g7689));
AN2X1 gate8090(.O (g4465), .I1 (g1117), .I2 (g3828));
AN2X1 gate8091(.O (g7141), .I1 (g6073), .I2 (g6716));
AN2X1 gate8092(.O (g10508), .I1 (g10391), .I2 (g2135));
AN2X1 gate8093(.O (g4230), .I1 (g1095), .I2 (g3638));
AN2X1 gate8094(.O (g10634), .I1 (g10604), .I2 (g3829));
AN2X1 gate8095(.O (g9601), .I1 (g922), .I2 (g9192));
AN2X1 gate8096(.O (g6126), .I1 (g5639), .I2 (g4319));
AN2X1 gate8097(.O (g6326), .I1 (g1250), .I2 (g5949));
AN2X1 gate8098(.O (g7710), .I1 (g700), .I2 (g7214));
AN2X1 gate8099(.O (g8028), .I1 (g7375), .I2 (g7436));
AN2X1 gate8100(.O (g6760), .I1 (g786), .I2 (g6221));
AN2X1 gate8101(.O (g5640), .I1 (g1059), .I2 (g4427));
AN2X1 gate8102(.O (g5031), .I1 (g1478), .I2 (g4640));
AN2X1 gate8103(.O (g4550), .I1 (g342), .I2 (g3586));
AN2X1 gate8104(.O (g7879), .I1 (g7610), .I2 (g3798));
AN2X1 gate8105(.O (g7962), .I1 (g7730), .I2 (g6712));
AN2X1 gate8106(.O (g9597), .I1 (g1170), .I2 (g9125));
AN2X1 gate8107(.O (g10452), .I1 (g10439), .I2 (g3388));
AN2X1 gate8108(.O (g4891), .I1 (g631), .I2 (g4739));
AN2X1 gate8109(.O (g5005), .I1 (g1490), .I2 (g4640));
AN2X1 gate8110(.O (g6423), .I1 (g4348), .I2 (g5784));
AN2X1 gate8111(.O (g8108), .I1 (g1891), .I2 (g7938));
AN3X1 gate8112(.O (g4807), .I1 (g3015), .I2 (g1289), .I3 (g3937));
AN2X1 gate8113(.O (g5911), .I1 (g3322), .I2 (g4977));
AN2X1 gate8114(.O (g9937), .I1 (g9916), .I2 (g9624));
AN2X1 gate8115(.O (g9840), .I1 (g9704), .I2 (g9747));
AN2X1 gate8116(.O (g10780), .I1 (g10723), .I2 (g5124));
AN2X1 gate8117(.O (g8217), .I1 (g1872), .I2 (g7883));
AN2X1 gate8118(.O (g11013), .I1 (g5209), .I2 (g10827));
AN2X1 gate8119(.O (g9390), .I1 (g1333), .I2 (g9151));
AN2X1 gate8120(.O (g11214), .I1 (g950), .I2 (g11159));
AN2X1 gate8121(.O (g6327), .I1 (g1255), .I2 (g5949));
AN2X1 gate8122(.O (g4342), .I1 (g1149), .I2 (g3719));
AN2X1 gate8123(.O (g5796), .I1 (g1564), .I2 (g5252));
AN2X1 gate8124(.O (g5473), .I1 (g4268), .I2 (g3518));
AN2X1 gate8125(.O (g6346), .I1 (g5038), .I2 (g5883));
AN2X1 gate8126(.O (g6633), .I1 (g354), .I2 (g6191));
AN2X1 gate8127(.O (g11005), .I1 (g5119), .I2 (g10827));
AN2X1 gate8128(.O (g8365), .I1 (g668), .I2 (g8240));
AN2X1 gate8129(.O (g8048), .I1 (g7558), .I2 (g5919));
AN2X1 gate8130(.O (g4481), .I1 (g1713), .I2 (g3906));
AN2X1 gate8131(.O (g4097), .I1 (g2677), .I2 (g2989));
AN2X1 gate8132(.O (g8055), .I1 (g7588), .I2 (g5128));
AN2X1 gate8133(.O (g4497), .I1 (g351), .I2 (g3586));
AN2X1 gate8134(.O (g9942), .I1 (g9922), .I2 (g9367));
AN2X1 gate8135(.O (g6696), .I1 (g5504), .I2 (g5850));
AN3X1 gate8136(.O (g10731), .I1 (g5118), .I2 (g1850), .I3 (g10665));
AN2X1 gate8137(.O (g8827), .I1 (g8552), .I2 (g8696));
AN2X1 gate8138(.O (g5540), .I1 (g1727), .I2 (g4315));
AN2X1 gate8139(.O (g4960), .I1 (g1403), .I2 (g4682));
AN2X1 gate8140(.O (g8846), .I1 (g8615), .I2 (g8712));
AN2X1 gate8141(.O (g6508), .I1 (g5983), .I2 (g3096));
AN2X1 gate8142(.O (g6240), .I1 (g182), .I2 (g5361));
AN2X1 gate8143(.O (g7931), .I1 (g2809), .I2 (g7446));
AN2X1 gate8144(.O (g5287), .I1 (g3876), .I2 (g4782));
AN2X1 gate8145(.O (g6472), .I1 (g5853), .I2 (g1936));
AN2X1 gate8146(.O (g11100), .I1 (g853), .I2 (g10950));
AN2X1 gate8147(.O (g11235), .I1 (g5443), .I2 (g11107));
AN2X1 gate8148(.O (g5199), .I1 (g1068), .I2 (g4719));
AN2X1 gate8149(.O (g6316), .I1 (g1270), .I2 (g5949));
AN2X1 gate8150(.O (g7515), .I1 (g7148), .I2 (g2855));
AN2X1 gate8151(.O (g10583), .I1 (g10518), .I2 (g10515));
AN2X1 gate8152(.O (g5781), .I1 (g1537), .I2 (g5222));
AN2X1 gate8153(.O (g8018), .I1 (g7742), .I2 (g7425));
AN2X1 gate8154(.O (g4401), .I1 (g2971), .I2 (g3772));
AN3X1 gate8155(.O (g8994), .I1 (g8110), .I2 (g6778), .I3 (g8925));
AN2X1 gate8156(.O (g2950), .I1 (g2424), .I2 (g1666));
AN2X1 gate8157(.O (g5510), .I1 (g1630), .I2 (g4280));
AN2X1 gate8158(.O (g6347), .I1 (g275), .I2 (g5890));
AN2X1 gate8159(.O (g9357), .I1 (g962), .I2 (g9223));
AN2X1 gate8160(.O (g4828), .I1 (g4106), .I2 (g695));
AN2X1 gate8161(.O (g11407), .I1 (g11339), .I2 (g5949));
AN2X1 gate8162(.O (g4727), .I1 (g386), .I2 (g3364));
AN2X1 gate8163(.O (g10357), .I1 (g10278), .I2 (g2462));
AN2X1 gate8164(.O (g10743), .I1 (g10639), .I2 (g4013));
AN2X1 gate8165(.O (g5259), .I1 (g627), .I2 (g4739));
AN2X1 gate8166(.O (g5694), .I1 (g162), .I2 (g5361));
AN2X1 gate8167(.O (g10769), .I1 (g10652), .I2 (g4840));
AN2X1 gate8168(.O (g11584), .I1 (g1318), .I2 (g11542));
AN2X1 gate8169(.O (g4932), .I1 (g1065), .I2 (g4442));
AN2X1 gate8170(.O (g10768), .I1 (g10649), .I2 (g4840));
AN2X1 gate8171(.O (g6820), .I1 (g1362), .I2 (g6596));
AN2X1 gate8172(.O (g4068), .I1 (g2719), .I2 (g2276));
AN2X1 gate8173(.O (g6317), .I1 (g1304), .I2 (g5949));
AN2X1 gate8174(.O (g5215), .I1 (g4276), .I2 (g3400));
AN2X1 gate8175(.O (g4576), .I1 (g530), .I2 (g4049));
AN2X1 gate8176(.O (g4866), .I1 (g231), .I2 (g3946));
AN2X1 gate8177(.O (g6775), .I1 (g822), .I2 (g6231));
AN2X1 gate8178(.O (g3829), .I1 (g2028), .I2 (g2728));
AN2X1 gate8179(.O (g10662), .I1 (g8892), .I2 (g10571));
AN2X1 gate8180(.O (g8101), .I1 (g6208), .I2 (g7877));
AN2X1 gate8181(.O (g5825), .I1 (g3204), .I2 (g5318));
AN4X1 gate8182(.O (I6310), .I1 (g2396), .I2 (g2407), .I3 (g2421), .I4 (g2435));
AN2X1 gate8183(.O (g7884), .I1 (g7457), .I2 (g7022));
AN2X1 gate8184(.O (g5008), .I1 (g1292), .I2 (g4507));
AN2X1 gate8185(.O (g3974), .I1 (g231), .I2 (g3164));
AN2X1 gate8186(.O (g9949), .I1 (g9929), .I2 (g9392));
AN2X1 gate8187(.O (g2531), .I1 (g658), .I2 (g668));
AN2X1 gate8188(.O (g9292), .I1 (g8878), .I2 (g5708));
AN2X1 gate8189(.O (g10778), .I1 (g1027), .I2 (g10729));
AN2X1 gate8190(.O (g8041), .I1 (g7524), .I2 (g5128));
AN2X1 gate8191(.O (g6079), .I1 (g1053), .I2 (g5320));
AN2X1 gate8192(.O (g7235), .I1 (g6663), .I2 (g6447));
AN2X1 gate8193(.O (g9603), .I1 (g1173), .I2 (g9125));
AN2X1 gate8194(.O (g6840), .I1 (g248), .I2 (g6596));
AN2X1 gate8195(.O (g9850), .I1 (g9726), .I2 (g9560));
AN2X1 gate8196(.O (g7988), .I1 (g1878), .I2 (g7379));
AN2X1 gate8197(.O (g5228), .I1 (g1086), .I2 (g4734));
AN2X1 gate8198(.O (g7134), .I1 (g5587), .I2 (g6354));
AN2X1 gate8199(.O (g5934), .I1 (g5215), .I2 (g1965));
AN2X1 gate8200(.O (g5230), .I1 (g1265), .I2 (g4735));
AN2X1 gate8201(.O (g8168), .I1 (g5262), .I2 (g7853));
AN2X1 gate8202(.O (g9583), .I1 (g886), .I2 (g8995));
AN2X1 gate8203(.O (g10672), .I1 (g10579), .I2 (g9449));
AN2X1 gate8204(.O (g3287), .I1 (g802), .I2 (g2534));
AN2X1 gate8205(.O (g8772), .I1 (g8627), .I2 (g5151));
AN2X1 gate8206(.O (g4893), .I1 (g635), .I2 (g4739));
AN2X1 gate8207(.O (g10331), .I1 (g10256), .I2 (g3307));
AN2X1 gate8208(.O (g8505), .I1 (g8309), .I2 (g4789));
AN2X1 gate8209(.O (g10449), .I1 (g10420), .I2 (g3345));
AN2X1 gate8210(.O (g11273), .I1 (g5638), .I2 (g11195));
AN2X1 gate8211(.O (g8734), .I1 (g8626), .I2 (g7923));
AN2X1 gate8212(.O (g5913), .I1 (g1041), .I2 (g5320));
AN2X1 gate8213(.O (g10448), .I1 (g10421), .I2 (g3335));
AN2X1 gate8214(.O (g6163), .I1 (g4572), .I2 (g5354));
AN2X1 gate8215(.O (g6363), .I1 (g284), .I2 (g5901));
AN2X1 gate8216(.O (g7202), .I1 (g6349), .I2 (g4329));
AN2X1 gate8217(.O (g11463), .I1 (g11432), .I2 (g5446));
AN2X1 gate8218(.O (g8074), .I1 (g718), .I2 (g7826));
AN2X1 gate8219(.O (g4325), .I1 (g1166), .I2 (g3682));
AN2X1 gate8220(.O (g8474), .I1 (g8383), .I2 (g5285));
AN2X1 gate8221(.O (g11234), .I1 (g5424), .I2 (g11106));
AN2X1 gate8222(.O (g5266), .I1 (g718), .I2 (g4766));
AN2X1 gate8223(.O (g4483), .I1 (g336), .I2 (g3586));
AN2X1 gate8224(.O (g5248), .I1 (g673), .I2 (g4738));
AN2X1 gate8225(.O (g11514), .I1 (g11491), .I2 (g5151));
AN2X1 gate8226(.O (g5255), .I1 (g682), .I2 (g4754));
AN2X1 gate8227(.O (g4106), .I1 (g3284), .I2 (g686));
AN2X1 gate8228(.O (g2760), .I1 (g981), .I2 (g2091));
AN2X1 gate8229(.O (g5097), .I1 (g1786), .I2 (g4603));
AN2X1 gate8230(.O (g5726), .I1 (g1601), .I2 (g5167));
AN2X1 gate8231(.O (g5497), .I1 (g4296), .I2 (g3522));
AN2X1 gate8232(.O (g5354), .I1 (g2733), .I2 (g4460));
AN2X1 gate8233(.O (g7933), .I1 (g2814), .I2 (g7450));
AN2X1 gate8234(.O (g9617), .I1 (g9), .I2 (g9274));
AN2X1 gate8235(.O (g9906), .I1 (g9873), .I2 (g9683));
AN2X1 gate8236(.O (g11012), .I1 (g5196), .I2 (g10827));
AN2X1 gate8237(.O (g7050), .I1 (g5896), .I2 (g6575));
AN2X1 gate8238(.O (g10971), .I1 (g10849), .I2 (g3161));
AN2X1 gate8239(.O (g4904), .I1 (g1850), .I2 (g4243));
AN2X1 gate8240(.O (g10369), .I1 (g10361), .I2 (g3382));
AN2X1 gate8241(.O (g8400), .I1 (g6097), .I2 (g8234));
AN2X1 gate8242(.O (g4345), .I1 (g1169), .I2 (g3730));
AN2X1 gate8243(.O (g2161), .I1 (I5084), .I2 (I5085));
AN2X1 gate8244(.O (g5001), .I1 (g1300), .I2 (g4491));
AN2X1 gate8245(.O (g9945), .I1 (g9925), .I2 (g9392));
AN2X1 gate8246(.O (g7271), .I1 (g5028), .I2 (g6499));
AN2X1 gate8247(.O (g9709), .I1 (g1524), .I2 (g9490));
AN2X1 gate8248(.O (g4223), .I1 (g1003), .I2 (g3914));
AN2X1 gate8249(.O (g10716), .I1 (g10497), .I2 (g10675));
AN2X1 gate8250(.O (g11291), .I1 (g11247), .I2 (g4233));
AN2X1 gate8251(.O (g6661), .I1 (g73), .I2 (g6219));
AN2X1 gate8252(.O (g11173), .I1 (g491), .I2 (g11112));
AN2X1 gate8253(.O (g6075), .I1 (g549), .I2 (g5613));
AN2X1 gate8254(.O (g8023), .I1 (g7367), .I2 (g7430));
AN2X1 gate8255(.O (g9907), .I1 (g9888), .I2 (g9686));
AN2X1 gate8256(.O (g10582), .I1 (g10532), .I2 (g9473));
AN2X1 gate8257(.O (g5746), .I1 (g1589), .I2 (g5193));
AN2X1 gate8258(.O (g5221), .I1 (g1260), .I2 (g4730));
AN2X1 gate8259(.O (g9959), .I1 (g9950), .I2 (g9536));
AN2X1 gate8260(.O (g7674), .I1 (g7004), .I2 (g3880));
AN2X1 gate8261(.O (g9690), .I1 (g266), .I2 (g9432));
AN2X1 gate8262(.O (g6627), .I1 (g58), .I2 (g6181));
AN2X1 gate8263(.O (g5703), .I1 (g174), .I2 (g5361));
AN2X1 gate8264(.O (g4522), .I1 (g360), .I2 (g3586));
AN2X1 gate8265(.O (g4115), .I1 (g2689), .I2 (g3009));
AN2X1 gate8266(.O (g7541), .I1 (g7075), .I2 (g3109));
AN2X1 gate8267(.O (g10627), .I1 (g10548), .I2 (g4564));
AN2X1 gate8268(.O (g4047), .I1 (g2695), .I2 (g2276));
AN2X1 gate8269(.O (g6526), .I1 (g76), .I2 (g6052));
AN2X1 gate8270(.O (g2944), .I1 (g2424), .I2 (g1669));
AN2X1 gate8271(.O (g6646), .I1 (g360), .I2 (g6203));
AN2X1 gate8272(.O (g7132), .I1 (g6048), .I2 (g6702));
AN2X1 gate8273(.O (g11029), .I1 (g401), .I2 (g10974));
AN2X1 gate8274(.O (g8051), .I1 (g7572), .I2 (g5128));
AN2X1 gate8275(.O (g8127), .I1 (g1927), .I2 (g7949));
AN2X1 gate8276(.O (g7209), .I1 (g3804), .I2 (g6425));
AN2X1 gate8277(.O (g11028), .I1 (g396), .I2 (g10974));
AN2X1 gate8278(.O (g6439), .I1 (g4479), .I2 (g5919));
AN2X1 gate8279(.O (g10742), .I1 (g10655), .I2 (g3586));
AN2X1 gate8280(.O (g9110), .I1 (g8880), .I2 (g4790));
AN2X1 gate8281(.O (g10681), .I1 (g10567), .I2 (g3586));
AN2X1 gate8282(.O (g4537), .I1 (g444), .I2 (g3988));
AN2X1 gate8283(.O (g9663), .I1 (g959), .I2 (g9223));
AN2X1 gate8284(.O (g5349), .I1 (g2126), .I2 (g4617));
AN2X1 gate8285(.O (g8732), .I1 (g8624), .I2 (g7919));
AN2X1 gate8286(.O (g3807), .I1 (g3003), .I2 (g3062));
AN2X1 gate8287(.O (g8753), .I1 (g7414), .I2 (g8664));
AN2X1 gate8288(.O (g5848), .I1 (g3860), .I2 (g5519));
AN2X1 gate8289(.O (g8508), .I1 (g8411), .I2 (g7967));
AN2X1 gate8290(.O (g8072), .I1 (g700), .I2 (g7826));
AN2X1 gate8291(.O (g5699), .I1 (g1592), .I2 (g5117));
AN2X1 gate8292(.O (g11240), .I1 (g5481), .I2 (g11111));
AN2X1 gate8293(.O (g5398), .I1 (g4610), .I2 (g2224));
AN2X1 gate8294(.O (g6616), .I1 (g6105), .I2 (g3246));
AN2X1 gate8295(.O (g10690), .I1 (g10616), .I2 (g3863));
AN2X1 gate8296(.O (g8043), .I1 (g7582), .I2 (g5128));
AN2X1 gate8297(.O (g9590), .I1 (g895), .I2 (g8995));
AN2X1 gate8298(.O (g4128), .I1 (g1976), .I2 (g2779));
AN2X1 gate8299(.O (g6404), .I1 (g2132), .I2 (g5748));
AN2X1 gate8300(.O (g6647), .I1 (g5288), .I2 (g5808));
AN2X1 gate8301(.O (g10504), .I1 (g10389), .I2 (g2135));
AN2X1 gate8302(.O (g9657), .I1 (g919), .I2 (g9205));
AN2X1 gate8303(.O (g4542), .I1 (g366), .I2 (g3586));
AN2X1 gate8304(.O (g4330), .I1 (g1163), .I2 (g3693));
AN2X1 gate8305(.O (g3497), .I1 (g2804), .I2 (g1900));
AN2X1 gate8306(.O (g5524), .I1 (g1678), .I2 (g4291));
AN2X1 gate8307(.O (g8147), .I1 (g2955), .I2 (g7961));
AN2X1 gate8308(.O (g4554), .I1 (g542), .I2 (g3996));
AN2X1 gate8309(.O (g9899), .I1 (g9889), .I2 (g9367));
AN2X1 gate8310(.O (g5258), .I1 (g700), .I2 (g4756));
AN2X1 gate8311(.O (g7736), .I1 (g6951), .I2 (g3880));
AN2X1 gate8312(.O (g6224), .I1 (g1520), .I2 (g5151));
AN2X1 gate8313(.O (g10626), .I1 (g10547), .I2 (g4558));
AN2X1 gate8314(.O (g6320), .I1 (g1292), .I2 (g5949));
AN2X1 gate8315(.O (g7623), .I1 (g664), .I2 (g7079));
AN2X1 gate8316(.O (g10299), .I1 (g8892), .I2 (g10217));
AN2X1 gate8317(.O (g7889), .I1 (g7615), .I2 (g3814));
AN2X1 gate8318(.O (g10298), .I1 (g8892), .I2 (g10214));
AN2X1 gate8319(.O (g8413), .I1 (g722), .I2 (g8146));
AN2X1 gate8320(.O (g3979), .I1 (g237), .I2 (g3164));
AN2X1 gate8321(.O (g4902), .I1 (g1848), .I2 (g4243));
AN2X1 gate8322(.O (g5211), .I1 (g1080), .I2 (g4724));
AN2X1 gate8323(.O (g4512), .I1 (g357), .I2 (g3586));
AN2X1 gate8324(.O (g7722), .I1 (g7127), .I2 (g6449));
AN2X1 gate8325(.O (g9844), .I1 (g9714), .I2 (g9522));
AN2X1 gate8326(.O (g4490), .I1 (g1141), .I2 (g3913));
AN2X1 gate8327(.O (g4823), .I1 (g207), .I2 (g3946));
AN2X1 gate8328(.O (g6516), .I1 (g5993), .I2 (g3097));
AN2X1 gate8329(.O (g5026), .I1 (g1453), .I2 (g4640));
AN2X1 gate8330(.O (g8820), .I1 (g8705), .I2 (g5422));
AN2X1 gate8331(.O (g10737), .I1 (g10687), .I2 (g4840));
AN3X1 gate8332(.O (g8936), .I1 (g8115), .I2 (g6778), .I3 (g8849));
AN2X1 gate8333(.O (g10232), .I1 (g8892), .I2 (g10150));
AN2X1 gate8334(.O (g6771), .I1 (g263), .I2 (g5866));
AN2X1 gate8335(.O (g5170), .I1 (g1811), .I2 (g4680));
AN2X1 gate8336(.O (g8117), .I1 (g6236), .I2 (g7886));
AN2X1 gate8337(.O (g4529), .I1 (g448), .I2 (g3980));
AN2X1 gate8338(.O (g4348), .I1 (g3497), .I2 (g1909));
AN2X1 gate8339(.O (g9966), .I1 (g9956), .I2 (g9536));
AN2X1 gate8340(.O (g5280), .I1 (g4593), .I2 (g3052));
AN2X1 gate8341(.O (g7139), .I1 (g6060), .I2 (g6709));
AN2X1 gate8342(.O (g11099), .I1 (g382), .I2 (g10885));
AN2X1 gate8343(.O (g6892), .I1 (g6472), .I2 (g5805));
AN2X1 gate8344(.O (g9705), .I1 (g1580), .I2 (g9474));
AN2X1 gate8345(.O (g10512), .I1 (g10395), .I2 (g2135));
AN2X1 gate8346(.O (g11098), .I1 (g849), .I2 (g10950));
AN2X1 gate8347(.O (g8775), .I1 (g8628), .I2 (g5151));
AN2X1 gate8348(.O (g5083), .I1 (g3709), .I2 (g4586));
AN2X1 gate8349(.O (g5544), .I1 (g1687), .I2 (g4320));
AN2X1 gate8350(.O (g11272), .I1 (g5629), .I2 (g11193));
AN2X1 gate8351(.O (g5483), .I1 (g1621), .I2 (g4254));
AN2X1 gate8352(.O (g9948), .I1 (g9928), .I2 (g9392));
AN2X1 gate8353(.O (g4063), .I1 (g2713), .I2 (g2276));
AN2X1 gate8354(.O (g11462), .I1 (g11431), .I2 (g5446));
AN2X1 gate8355(.O (g6738), .I1 (g2531), .I2 (g6137));
AN2X1 gate8356(.O (g8060), .I1 (g7593), .I2 (g5919));
AN2X1 gate8357(.O (g6244), .I1 (g2255), .I2 (g5151));
AN2X1 gate8358(.O (g11032), .I1 (g416), .I2 (g10974));
AN2X1 gate8359(.O (g10445), .I1 (g10315), .I2 (g2135));
AN2X1 gate8360(.O (g9150), .I1 (g8882), .I2 (g4805));
AN2X1 gate8361(.O (g10316), .I1 (g10223), .I2 (g9097));
AN2X1 gate8362(.O (g5756), .I1 (g1531), .I2 (g5202));
AN2X1 gate8363(.O (g4720), .I1 (g1023), .I2 (g3914));
AN2X1 gate8364(.O (g9409), .I1 (g1721), .I2 (g9052));
AN2X1 gate8365(.O (g8995), .I1 (g6454), .I2 (g8929));
AN2X1 gate8366(.O (g6876), .I1 (g4070), .I2 (g6560));
AN2X1 gate8367(.O (g4989), .I1 (g1424), .I2 (g4682));
AN2X1 gate8368(.O (g9836), .I1 (g9737), .I2 (g9785));
AN3X1 gate8369(.O (g6656), .I1 (g2733), .I2 (g6061), .I3 (g4631));
AN2X1 gate8370(.O (g5514), .I1 (g1941), .I2 (g4284));
AN2X1 gate8371(.O (g8390), .I1 (g8268), .I2 (g6465));
AN2X1 gate8372(.O (g5003), .I1 (g1466), .I2 (g4640));
AN2X1 gate8373(.O (g9967), .I1 (g9957), .I2 (g9536));
AN2X1 gate8374(.O (g5145), .I1 (g1639), .I2 (g4673));
AN2X1 gate8375(.O (g4834), .I1 (g219), .I2 (g3946));
AN2X1 gate8376(.O (g4971), .I1 (g1419), .I2 (g4682));
AN2X1 gate8377(.O (g10753), .I1 (g10649), .I2 (g4013));
AN2X1 gate8378(.O (g5695), .I1 (g166), .I2 (g5361));
AN2X1 gate8379(.O (g7613), .I1 (g6940), .I2 (g5984));
AN2X1 gate8380(.O (g10736), .I1 (g10658), .I2 (g4840));
AN2X1 gate8381(.O (g11220), .I1 (g962), .I2 (g11054));
AN2X1 gate8382(.O (g7444), .I1 (g7277), .I2 (g5827));
AN2X1 gate8383(.O (g5536), .I1 (g4867), .I2 (g4298));
AN2X1 gate8384(.O (g6663), .I1 (g6064), .I2 (g2237));
AN2X1 gate8385(.O (g4670), .I1 (g192), .I2 (g3946));
AN2X1 gate8386(.O (g6824), .I1 (g1371), .I2 (g6596));
AN2X1 gate8387(.O (g4253), .I1 (g1074), .I2 (g3638));
AN2X1 gate8388(.O (g8250), .I1 (g2771), .I2 (g7907));
AN2X1 gate8389(.O (g8163), .I1 (g7960), .I2 (g3737));
AN2X1 gate8390(.O (g10764), .I1 (g10643), .I2 (g4840));
AN2X1 gate8391(.O (g5757), .I1 (g1552), .I2 (g5203));
AN2X1 gate8392(.O (g10365), .I1 (g10319), .I2 (g2135));
AN2X1 gate8393(.O (g8032), .I1 (g7385), .I2 (g7438));
AN2X1 gate8394(.O (g11591), .I1 (g2988), .I2 (g11561));
AN2X1 gate8395(.O (g8053), .I1 (g7583), .I2 (g5919));
AN2X1 gate8396(.O (g11147), .I1 (g321), .I2 (g10929));
AN2X1 gate8397(.O (g5522), .I1 (g1633), .I2 (g4289));
AN2X1 gate8398(.O (g5115), .I1 (g1394), .I2 (g4572));
AN2X1 gate8399(.O (g9837), .I1 (g9697), .I2 (g9751));
AN2X1 gate8400(.O (g9620), .I1 (g2653), .I2 (g9240));
AN2X1 gate8401(.O (g11151), .I1 (g327), .I2 (g10931));
AN2X1 gate8402(.O (g11172), .I1 (g486), .I2 (g11112));
AN2X1 gate8403(.O (g7885), .I1 (g7614), .I2 (g3812));
AN2X1 gate8404(.O (g6064), .I1 (g5398), .I2 (g2230));
AN3X1 gate8405(.O (g8929), .I1 (g8095), .I2 (g6368), .I3 (g8828));
AN2X1 gate8406(.O (g5595), .I1 (g1621), .I2 (g4524));
AN2X1 gate8407(.O (g5537), .I1 (g4143), .I2 (g4299));
AN2X1 gate8408(.O (g9842), .I1 (g9708), .I2 (g9516));
AN2X1 gate8409(.O (g4141), .I1 (g2707), .I2 (g3051));
AN2X1 gate8410(.O (g4341), .I1 (g339), .I2 (g3586));
AN2X1 gate8411(.O (g9192), .I1 (g6454), .I2 (g8955));
AN2X1 gate8412(.O (g7679), .I1 (g1950), .I2 (g6863));
AN2X1 gate8413(.O (g7378), .I1 (g6990), .I2 (g3880));
AN2X1 gate8414(.O (g5612), .I1 (g1627), .I2 (g4543));
AN2X1 gate8415(.O (g3939), .I1 (g213), .I2 (g3164));
AN2X1 gate8416(.O (g7135), .I1 (g869), .I2 (g6355));
AN2X1 gate8417(.O (g10970), .I1 (g10852), .I2 (g3390));
AN2X1 gate8418(.O (g11025), .I1 (g426), .I2 (g10974));
AN2X1 gate8419(.O (g9854), .I1 (g9730), .I2 (g9566));
AN2X1 gate8420(.O (g7182), .I1 (g1878), .I2 (g6720));
AN2X1 gate8421(.O (g9941), .I1 (g9921), .I2 (g9367));
AN2X1 gate8422(.O (g6194), .I1 (g554), .I2 (g5043));
AN2X1 gate8423(.O (g5128), .I1 (g4474), .I2 (g2733));
AN2X1 gate8424(.O (g4962), .I1 (g1651), .I2 (g4461));
AN2X1 gate8425(.O (g4358), .I1 (g1209), .I2 (g3747));
AN2X1 gate8426(.O (g8683), .I1 (g4803), .I2 (g8549));
AN2X1 gate8427(.O (g4506), .I1 (g1113), .I2 (g3944));
AN2X1 gate8428(.O (g6471), .I1 (g5224), .I2 (g6014));
AN2X1 gate8429(.O (g8778), .I1 (g8688), .I2 (g2317));
AN2X1 gate8430(.O (g11281), .I1 (g4948), .I2 (g11202));
AN2X1 gate8431(.O (g8735), .I1 (g7600), .I2 (g8632));
AN2X1 gate8432(.O (g11146), .I1 (g318), .I2 (g10928));
AN2X1 gate8433(.O (g3904), .I1 (g2948), .I2 (g2779));
AN2X1 gate8434(.O (g8075), .I1 (g727), .I2 (g7826));
AN2X1 gate8435(.O (g9829), .I1 (g9723), .I2 (g9785));
AN3X1 gate8436(.O (g8949), .I1 (g8255), .I2 (g6368), .I3 (g8828));
AN2X1 gate8437(.O (g7632), .I1 (g7184), .I2 (g5574));
AN2X1 gate8438(.O (g11290), .I1 (g11246), .I2 (g4226));
AN2X1 gate8439(.O (g6350), .I1 (g5837), .I2 (g4435));
AN2X1 gate8440(.O (g10599), .I1 (g10534), .I2 (g4365));
AN2X1 gate8441(.O (g5902), .I1 (g2555), .I2 (g4977));
AN4X1 gate8442(.O (I6337), .I1 (g201), .I2 (g2421), .I3 (g2407), .I4 (g2396));
AN2X1 gate8443(.O (g2276), .I1 (g1765), .I2 (g1610));
AN2X1 gate8444(.O (g6438), .I1 (g5853), .I2 (g5797));
AN2X1 gate8445(.O (g5512), .I1 (g1660), .I2 (g4281));
AN2X1 gate8446(.O (g5090), .I1 (g1781), .I2 (g4592));
AN2X1 gate8447(.O (g7719), .I1 (g718), .I2 (g7227));
AN2X1 gate8448(.O (g2561), .I1 (g742), .I2 (g741));
AN2X1 gate8449(.O (g3695), .I1 (g1712), .I2 (g3015));
AN2X1 gate8450(.O (g8603), .I1 (g3983), .I2 (g8548));
AN2X1 gate8451(.O (g8039), .I1 (g7587), .I2 (g5128));
AN2X1 gate8452(.O (g9610), .I1 (g925), .I2 (g9192));
AN2X1 gate8453(.O (g3536), .I1 (g2390), .I2 (g3103));
AN2X1 gate8454(.O (g5529), .I1 (g4129), .I2 (g4288));
AN2X1 gate8455(.O (g5148), .I1 (g3088), .I2 (g4671));
AN2X1 gate8456(.O (g9124), .I1 (g8881), .I2 (g4802));
AN2X1 gate8457(.O (g9324), .I1 (g8879), .I2 (g5708));
AN2X1 gate8458(.O (g4559), .I1 (g2034), .I2 (g3829));
AN2X1 gate8459(.O (g10561), .I1 (g10549), .I2 (g4583));
AN2X1 gate8460(.O (g5698), .I1 (g1571), .I2 (g5116));
AN2X1 gate8461(.O (g11226), .I1 (g461), .I2 (g11057));
AN2X1 gate8462(.O (g10295), .I1 (g8892), .I2 (g10208));
AN2X1 gate8463(.O (g5260), .I1 (g1092), .I2 (g4758));
AN2X1 gate8464(.O (g10680), .I1 (g10564), .I2 (g3586));
AN2X1 gate8465(.O (g6822), .I1 (g231), .I2 (g6596));
AN2X1 gate8466(.O (g4905), .I1 (g1853), .I2 (g4243));
AN2X1 gate8467(.O (g11551), .I1 (g11538), .I2 (g4013));
AN2X1 gate8468(.O (g3047), .I1 (g1227), .I2 (g2306));
AN2X1 gate8469(.O (g9849), .I1 (g293), .I2 (g9768));
AN2X1 gate8470(.O (g5279), .I1 (g1766), .I2 (g4783));
AN2X1 gate8471(.O (g8404), .I1 (g686), .I2 (g8129));
AN2X1 gate8472(.O (g5720), .I1 (g170), .I2 (g5361));
AN2X1 gate8473(.O (g5318), .I1 (g4401), .I2 (g1857));
AN2X1 gate8474(.O (g8764), .I1 (g7443), .I2 (g8684));
AN2X1 gate8475(.O (g11376), .I1 (g11318), .I2 (g4277));
AN2X1 gate8476(.O (g11297), .I1 (g5490), .I2 (g11242));
AN2X1 gate8477(.O (g9898), .I1 (g9887), .I2 (g9367));
OR2X1 gate8478(.O (g6895), .I1 (g6776), .I2 (g4875));
OR2X1 gate8479(.O (g7189), .I1 (g6632), .I2 (g6053));
OR2X1 gate8480(.O (g9510), .I1 (g9125), .I2 (g9111));
OR2X1 gate8481(.O (g7297), .I1 (g7132), .I2 (g6323));
OR2X1 gate8482(.O (g9088), .I1 (g8927), .I2 (g8381));
OR2X1 gate8483(.O (g9923), .I1 (g9865), .I2 (g9707));
OR2X1 gate8484(.O (g6485), .I1 (g5848), .I2 (g5067));
OR2X1 gate8485(.O (g8771), .I1 (g5483), .I2 (g8652));
OR2X1 gate8486(.O (g5813), .I1 (g5617), .I2 (g4869));
OR2X1 gate8487(.O (g7963), .I1 (g7687), .I2 (g7182));
OR2X1 gate8488(.O (g10643), .I1 (g10624), .I2 (g7736));
OR3X1 gate8489(.O (g9886), .I1 (g9607), .I2 (g9592), .I3 (g9759));
OR3X1 gate8490(.O (g9951), .I1 (g9902), .I2 (g9899), .I3 (g9803));
OR2X1 gate8491(.O (g11625), .I1 (g6535), .I2 (g11597));
OR2X1 gate8492(.O (g8945), .I1 (g8801), .I2 (g8710));
OR2X1 gate8493(.O (g10489), .I1 (g4961), .I2 (g10367));
OR2X1 gate8494(.O (g10559), .I1 (g4141), .I2 (g10512));
OR2X1 gate8495(.O (g10558), .I1 (g4126), .I2 (g10510));
OR2X1 gate8496(.O (g11338), .I1 (g11283), .I2 (g11178));
OR2X1 gate8497(.O (g8435), .I1 (g8403), .I2 (g8075));
OR2X1 gate8498(.O (g10544), .I1 (g5511), .I2 (g10495));
OR2X1 gate8499(.O (g6911), .I1 (g6342), .I2 (g5681));
OR2X1 gate8500(.O (g10865), .I1 (g5538), .I2 (g10752));
OR2X1 gate8501(.O (g3698), .I1 (g3121), .I2 (g2480));
OR2X1 gate8502(.O (g8214), .I1 (g7472), .I2 (g8004));
OR2X1 gate8503(.O (g6124), .I1 (g5181), .I2 (g5188));
OR2X1 gate8504(.O (g6469), .I1 (g5698), .I2 (g4959));
OR2X1 gate8505(.O (g5587), .I1 (g4714), .I2 (g3904));
OR2X1 gate8506(.O (g6177), .I1 (g5444), .I2 (g4712));
OR3X1 gate8507(.O (I14585), .I1 (g8995), .I2 (g9205), .I3 (g9192));
OR2X1 gate8508(.O (g9891), .I1 (g9741), .I2 (g9760));
OR2X1 gate8509(.O (g9913), .I1 (g9849), .I2 (g9691));
OR4X1 gate8510(.O (I5600), .I1 (g496), .I2 (g491), .I3 (g486), .I4 (g481));
OR2X1 gate8511(.O (g11257), .I1 (g11234), .I2 (g11019));
OR2X1 gate8512(.O (g8236), .I1 (g7526), .I2 (g8001));
OR2X1 gate8513(.O (g7385), .I1 (g7235), .I2 (g6746));
OR2X1 gate8514(.O (g6898), .I1 (g6790), .I2 (g4881));
OR2X1 gate8515(.O (g6900), .I1 (g6787), .I2 (g6246));
OR2X1 gate8516(.O (g4264), .I1 (g4048), .I2 (g4053));
OR3X1 gate8517(.O (g9726), .I1 (g9411), .I2 (g9420), .I3 (g9489));
OR2X1 gate8518(.O (g6088), .I1 (g5260), .I2 (g4522));
OR2X1 gate8519(.O (g6923), .I1 (g6353), .I2 (g5695));
OR2X1 gate8520(.O (g8194), .I1 (g5168), .I2 (g7940));
OR3X1 gate8521(.O (g9676), .I1 (g9454), .I2 (g9292), .I3 (g9274));
OR2X1 gate8522(.O (g11256), .I1 (g11186), .I2 (g11018));
OR2X1 gate8523(.O (g3860), .I1 (g3107), .I2 (g2167));
OR2X1 gate8524(.O (g11280), .I1 (g11254), .I2 (g11153));
OR4X1 gate8525(.O (g9727), .I1 (g9650), .I2 (g9663), .I3 (g9362), .I4 (I14866));
OR2X1 gate8526(.O (g4997), .I1 (g4581), .I2 (g4584));
OR2X1 gate8527(.O (g11624), .I1 (g11595), .I2 (g11571));
OR2X1 gate8528(.O (g11300), .I1 (g11213), .I2 (g11091));
OR2X1 gate8529(.O (g4238), .I1 (g3999), .I2 (g4007));
OR2X1 gate8530(.O (g8814), .I1 (g7945), .I2 (g8728));
OR2X1 gate8531(.O (g10401), .I1 (g9317), .I2 (g10291));
OR2X1 gate8532(.O (g8773), .I1 (g5491), .I2 (g8653));
OR2X1 gate8533(.O (g11231), .I1 (g11156), .I2 (g11013));
OR2X1 gate8534(.O (g10864), .I1 (g5532), .I2 (g10751));
OR2X1 gate8535(.O (g9624), .I1 (g9316), .I2 (g9313));
OR3X1 gate8536(.O (g9953), .I1 (g9945), .I2 (g9939), .I3 (g9669));
OR2X1 gate8537(.O (g6122), .I1 (g5172), .I2 (g5180));
OR2X1 gate8538(.O (g6465), .I1 (g5825), .I2 (g5041));
OR2X1 gate8539(.O (g6934), .I1 (g6363), .I2 (g5720));
OR2X1 gate8540(.O (g7664), .I1 (g6855), .I2 (g4084));
OR2X1 gate8541(.O (g7246), .I1 (g6465), .I2 (g6003));
OR2X1 gate8542(.O (g7203), .I1 (g6640), .I2 (g6058));
OR2X1 gate8543(.O (g6096), .I1 (g5268), .I2 (g4542));
OR2X1 gate8544(.O (g9747), .I1 (g9173), .I2 (g9509));
OR2X1 gate8545(.O (g11314), .I1 (g11224), .I2 (g11102));
OR2X1 gate8546(.O (g10733), .I1 (g5227), .I2 (g10674));
OR2X1 gate8547(.O (g8921), .I1 (g8827), .I2 (g8748));
OR4X1 gate8548(.O (I15054), .I1 (g7853), .I2 (g9782), .I3 (g9624), .I4 (g9785));
OR2X1 gate8549(.O (g11269), .I1 (g11196), .I2 (g11031));
OR2X1 gate8550(.O (g5555), .I1 (g4389), .I2 (g4397));
OR2X1 gate8551(.O (g11268), .I1 (g11194), .I2 (g11030));
OR2X1 gate8552(.O (g10485), .I1 (g9317), .I2 (g10376));
OR2X1 gate8553(.O (g10555), .I1 (g4103), .I2 (g10504));
OR2X1 gate8554(.O (g6481), .I1 (g5722), .I2 (g4972));
OR2X1 gate8555(.O (g10712), .I1 (g10662), .I2 (g9531));
OR2X1 gate8556(.O (g11335), .I1 (g11279), .I2 (g11175));
OR2X1 gate8557(.O (g8249), .I1 (g8018), .I2 (g7710));
OR2X1 gate8558(.O (g7638), .I1 (g7265), .I2 (g6488));
OR2X1 gate8559(.O (g10567), .I1 (g10514), .I2 (g7378));
OR2X1 gate8560(.O (g11487), .I1 (g6662), .I2 (g11464));
OR4X1 gate8561(.O (I15210), .I1 (g9839), .I2 (g9964), .I3 (g9852), .I4 (g9882));
OR4X1 gate8562(.O (I5805), .I1 (g2102), .I2 (g2099), .I3 (g2096), .I4 (g2088));
OR2X1 gate8563(.O (g8941), .I1 (g8796), .I2 (g8706));
OR2X1 gate8564(.O (g11443), .I1 (g7130), .I2 (g11407));
OR2X1 gate8565(.O (g4231), .I1 (g3991), .I2 (g3998));
OR2X1 gate8566(.O (g11278), .I1 (g11253), .I2 (g11150));
OR4X1 gate8567(.O (I15039), .I1 (g7853), .I2 (g9809), .I3 (g9624), .I4 (g9785));
OR2X1 gate8568(.O (g11286), .I1 (g10670), .I2 (g11209));
OR2X1 gate8569(.O (g8431), .I1 (g8387), .I2 (g8071));
OR2X1 gate8570(.O (g7133), .I1 (g6616), .I2 (g3067));
OR2X1 gate8571(.O (g11306), .I1 (g11216), .I2 (g11095));
OR2X1 gate8572(.O (g8252), .I1 (g7988), .I2 (g7679));
OR2X1 gate8573(.O (g8812), .I1 (g7939), .I2 (g8724));
OR2X1 gate8574(.O (g7846), .I1 (g7722), .I2 (g7241));
OR2X1 gate8575(.O (g3875), .I1 (g3275), .I2 (g12));
OR2X1 gate8576(.O (g5996), .I1 (g5473), .I2 (g3908));
OR2X1 gate8577(.O (g6592), .I1 (g5100), .I2 (g5882));
OR2X1 gate8578(.O (g8286), .I1 (g8107), .I2 (g7823));
OR2X1 gate8579(.O (g10501), .I1 (g4161), .I2 (g10445));
OR2X1 gate8580(.O (g10728), .I1 (g4973), .I2 (g10642));
OR2X1 gate8581(.O (g8270), .I1 (g7894), .I2 (g3434));
OR2X1 gate8582(.O (g7290), .I1 (g7046), .I2 (g6316));
OR2X1 gate8583(.O (g6068), .I1 (g5220), .I2 (g4497));
OR2X1 gate8584(.O (g6468), .I1 (g5690), .I2 (g4950));
OR2X1 gate8585(.O (g11217), .I1 (g11144), .I2 (g11005));
OR2X1 gate8586(.O (g11478), .I1 (g6532), .I2 (g11455));
OR4X1 gate8587(.O (g9536), .I1 (g9335), .I2 (g9331), .I3 (g9328), .I4 (g9324));
OR2X1 gate8588(.O (g5981), .I1 (g5074), .I2 (g4383));
OR2X1 gate8589(.O (g11486), .I1 (g6654), .I2 (g11463));
OR2X1 gate8590(.O (g8377), .I1 (g8185), .I2 (g7958));
OR2X1 gate8591(.O (g8206), .I1 (g7459), .I2 (g8007));
OR2X1 gate8592(.O (g11580), .I1 (g11413), .I2 (g11544));
OR2X1 gate8593(.O (g8287), .I1 (g8117), .I2 (g7824));
OR2X1 gate8594(.O (g11223), .I1 (g11147), .I2 (g11008));
OR2X1 gate8595(.O (g9522), .I1 (g9173), .I2 (g9125));
OR2X1 gate8596(.O (g8199), .I1 (g7902), .I2 (g7444));
OR2X1 gate8597(.O (g5802), .I1 (g5601), .I2 (g4837));
OR2X1 gate8598(.O (g11321), .I1 (g11230), .I2 (g11105));
OR2X1 gate8599(.O (g6524), .I1 (g5746), .I2 (g4996));
OR2X1 gate8600(.O (g10664), .I1 (g10240), .I2 (g10582));
OR2X1 gate8601(.O (g7257), .I1 (g6701), .I2 (g4725));
OR2X1 gate8602(.O (g7301), .I1 (g7140), .I2 (g6327));
OR2X1 gate8603(.O (g10484), .I1 (g9317), .I2 (g10400));
OR2X1 gate8604(.O (g10554), .I1 (g4097), .I2 (g10503));
OR2X1 gate8605(.O (g8259), .I1 (g8028), .I2 (g7719));
OR2X1 gate8606(.O (g11334), .I1 (g11277), .I2 (g11174));
OR2X1 gate8607(.O (g8819), .I1 (g7957), .I2 (g8734));
OR2X1 gate8608(.O (g8923), .I1 (g8846), .I2 (g8763));
OR2X1 gate8609(.O (g8488), .I1 (g3664), .I2 (g8390));
OR2X1 gate8610(.O (g7441), .I1 (g7271), .I2 (g6789));
OR2X1 gate8611(.O (g6026), .I1 (g5507), .I2 (g3970));
OR2X1 gate8612(.O (g10799), .I1 (g6225), .I2 (g10769));
OR2X1 gate8613(.O (g10798), .I1 (g6217), .I2 (g10768));
OR2X1 gate8614(.O (g10805), .I1 (g10759), .I2 (g10760));
OR2X1 gate8615(.O (g10732), .I1 (g4358), .I2 (g10661));
OR2X1 gate8616(.O (g6061), .I1 (g5204), .I2 (g4));
OR2X1 gate8617(.O (g9512), .I1 (g9151), .I2 (g9125));
OR2X1 gate8618(.O (g10013), .I1 (I15214), .I2 (I15215));
OR2X1 gate8619(.O (g8806), .I1 (g7931), .I2 (g8718));
OR2X1 gate8620(.O (g8943), .I1 (g8837), .I2 (g8749));
OR2X1 gate8621(.O (g11293), .I1 (g11211), .I2 (g10818));
OR2X1 gate8622(.O (g11265), .I1 (g11189), .I2 (g11027));
OR2X1 gate8623(.O (g8887), .I1 (g8842), .I2 (g8755));
OR2X1 gate8624(.O (g5838), .I1 (g5612), .I2 (g4866));
OR2X1 gate8625(.O (g6514), .I1 (g5738), .I2 (g4992));
OR2X1 gate8626(.O (g8322), .I1 (g8136), .I2 (g6891));
OR2X1 gate8627(.O (g8230), .I1 (g7515), .I2 (g7991));
OR2X1 gate8628(.O (g5809), .I1 (g5611), .I2 (g4865));
OR2X1 gate8629(.O (g8433), .I1 (g8399), .I2 (g8073));
OR2X1 gate8630(.O (g11579), .I1 (g5123), .I2 (g11551));
OR2X1 gate8631(.O (g10771), .I1 (g5533), .I2 (g10684));
OR2X1 gate8632(.O (g11615), .I1 (g11601), .I2 (g11592));
OR2X1 gate8633(.O (g9367), .I1 (g9335), .I2 (g9331));
OR3X1 gate8634(.O (g9872), .I1 (g9617), .I2 (g9594), .I3 (g9750));
OR2X1 gate8635(.O (g6522), .I1 (g5744), .I2 (g4994));
OR2X1 gate8636(.O (g8266), .I1 (g7885), .I2 (g3412));
OR2X1 gate8637(.O (g10414), .I1 (g10300), .I2 (g9534));
OR2X1 gate8638(.O (g11275), .I1 (g11248), .I2 (g11148));
OR2X1 gate8639(.O (g11430), .I1 (g11387), .I2 (g4006));
OR2X1 gate8640(.O (g8248), .I1 (g8014), .I2 (g7707));
OR3X1 gate8641(.O (g9686), .I1 (g9454), .I2 (g9292), .I3 (g9274));
OR2X1 gate8642(.O (g8815), .I1 (g7948), .I2 (g8730));
OR2X1 gate8643(.O (g7183), .I1 (g6623), .I2 (g6046));
OR2X1 gate8644(.O (g5983), .I1 (g5084), .I2 (g4392));
OR2X1 gate8645(.O (g8154), .I1 (g7891), .I2 (g6879));
OR2X1 gate8646(.O (g6537), .I1 (g5781), .I2 (g5005));
OR2X1 gate8647(.O (g4309), .I1 (g4069), .I2 (g4079));
OR2X1 gate8648(.O (g10725), .I1 (g4962), .I2 (g10634));
OR2X1 gate8649(.O (g6243), .I1 (g5537), .I2 (g4774));
OR4X1 gate8650(.O (I6351), .I1 (g2405), .I2 (g2389), .I3 (g2380), .I4 (g2372));
OR3X1 gate8651(.O (g9519), .I1 (g9173), .I2 (g9151), .I3 (g9125));
OR2X1 gate8652(.O (g9740), .I1 (g9418), .I2 (g9505));
OR2X1 gate8653(.O (g8267), .I1 (g7889), .I2 (g3422));
OR3X1 gate8654(.O (g10744), .I1 (g10600), .I2 (g10668), .I3 (I16427));
OR2X1 gate8655(.O (g6542), .I1 (g5789), .I2 (g5010));
OR2X1 gate8656(.O (g7303), .I1 (g7145), .I2 (g6329));
OR2X1 gate8657(.O (g10652), .I1 (g10627), .I2 (g7743));
OR2X1 gate8658(.O (g5036), .I1 (g4871), .I2 (g4162));
OR2X1 gate8659(.O (g7240), .I1 (g6687), .I2 (g6095));
OR2X1 gate8660(.O (g8221), .I1 (g7496), .I2 (g7993));
OR2X1 gate8661(.O (g6902), .I1 (g6794), .I2 (g4223));
OR3X1 gate8662(.O (I14776), .I1 (g8995), .I2 (g9205), .I3 (g9192));
OR2X1 gate8663(.O (g10500), .I1 (g4157), .I2 (g10442));
OR2X1 gate8664(.O (g4052), .I1 (g2862), .I2 (g2515));
OR4X1 gate8665(.O (I14858), .I1 (g9585), .I2 (g9595), .I3 (g9610), .I4 (g9602));
OR2X1 gate8666(.O (g6529), .I1 (g5757), .I2 (g5000));
OR2X1 gate8667(.O (g11264), .I1 (g11188), .I2 (g11026));
OR4X1 gate8668(.O (I15209), .I1 (g8169), .I2 (g9905), .I3 (g9934), .I4 (g9830));
OR2X1 gate8669(.O (g8241), .I1 (g7536), .I2 (g7989));
OR2X1 gate8670(.O (g10795), .I1 (g6199), .I2 (g10764));
OR2X1 gate8671(.O (g11607), .I1 (g11586), .I2 (g11557));
OR2X1 gate8672(.O (g8644), .I1 (g8123), .I2 (g8464));
OR3X1 gate8673(.O (g4682), .I1 (g3563), .I2 (g3348), .I3 (g1570));
OR2X1 gate8674(.O (g8818), .I1 (g7955), .I2 (g8733));
OR2X1 gate8675(.O (g2984), .I1 (g2528), .I2 (g2522));
OR2X1 gate8676(.O (g9931), .I1 (g8931), .I2 (g9900));
OR2X1 gate8677(.O (g3414), .I1 (g2911), .I2 (g2917));
OR2X1 gate8678(.O (g9515), .I1 (g9173), .I2 (g9151));
OR2X1 gate8679(.O (g10724), .I1 (g10312), .I2 (g10672));
OR2X1 gate8680(.O (g7294), .I1 (g7068), .I2 (g6320));
OR2X1 gate8681(.O (g5189), .I1 (g4345), .I2 (g3496));
OR2X1 gate8682(.O (g8614), .I1 (g8365), .I2 (g8510));
OR2X1 gate8683(.O (g3513), .I1 (g3118), .I2 (g2180));
OR2X1 gate8684(.O (g6909), .I1 (g6346), .I2 (g5684));
OR4X1 gate8685(.O (I5571), .I1 (g396), .I2 (g391), .I3 (g386), .I4 (g426));
OR2X1 gate8686(.O (g4283), .I1 (g4059), .I2 (g4063));
OR2X1 gate8687(.O (g8939), .I1 (g8791), .I2 (g8701));
OR2X1 gate8688(.O (g2514), .I1 (I5599), .I2 (I5600));
OR2X1 gate8689(.O (g11327), .I1 (g11297), .I2 (g11167));
OR2X1 gate8690(.O (g8187), .I1 (g7542), .I2 (g7998));
OR2X1 gate8691(.O (g11606), .I1 (g11585), .I2 (g11556));
OR2X1 gate8692(.O (g11303), .I1 (g11214), .I2 (g11092));
OR2X1 gate8693(.O (g5309), .I1 (g3664), .I2 (g4401));
OR3X1 gate8694(.O (g9528), .I1 (g9151), .I2 (g9125), .I3 (g9111));
OR2X1 gate8695(.O (g8200), .I1 (g7535), .I2 (g8008));
OR3X1 gate8696(.O (g2522), .I1 (g833), .I2 (g829), .I3 (I5629));
OR4X1 gate8697(.O (g2315), .I1 (g1163), .I2 (g1166), .I3 (g1113), .I4 (I5363));
OR2X1 gate8698(.O (g6506), .I1 (g5731), .I2 (g4989));
OR2X1 gate8699(.O (g10649), .I1 (g10626), .I2 (g7741));
OR2X1 gate8700(.O (g8159), .I1 (g7895), .I2 (g6886));
OR2X1 gate8701(.O (g7626), .I1 (g7060), .I2 (g5267));
OR2X1 gate8702(.O (g10770), .I1 (g5525), .I2 (g10682));
OR2X1 gate8703(.O (g9566), .I1 (g9052), .I2 (g9030));
OR2X1 gate8704(.O (g11483), .I1 (g6633), .I2 (g11460));
OR2X1 gate8705(.O (g8811), .I1 (g7935), .I2 (g8722));
OR3X1 gate8706(.O (g8642), .I1 (g5236), .I2 (g5205), .I3 (g8465));
OR2X1 gate8707(.O (g6545), .I1 (g5795), .I2 (g5025));
OR2X1 gate8708(.O (g10767), .I1 (g5500), .I2 (g10681));
OR2X1 gate8709(.O (g11326), .I1 (g11296), .I2 (g11166));
OR2X1 gate8710(.O (g10898), .I1 (g4220), .I2 (g10777));
OR2X1 gate8711(.O (g11252), .I1 (g11099), .I2 (g10969));
OR2X1 gate8712(.O (g10719), .I1 (g10303), .I2 (g10666));
OR2X1 gate8713(.O (g4609), .I1 (g3400), .I2 (g119));
OR2X1 gate8714(.O (g6507), .I1 (g5732), .I2 (g4990));
OR2X1 gate8715(.O (g10718), .I1 (g6238), .I2 (g10706));
OR2X1 gate8716(.O (g10521), .I1 (I16148), .I2 (I16149));
OR2X1 gate8717(.O (g7075), .I1 (g5104), .I2 (g6530));
OR2X1 gate8718(.O (g7292), .I1 (g7055), .I2 (g6318));
OR2X1 gate8719(.O (g10861), .I1 (g5523), .I2 (g10745));
OR2X1 gate8720(.O (g8417), .I1 (g8246), .I2 (g7721));
OR2X1 gate8721(.O (g6515), .I1 (g5739), .I2 (g4993));
OR4X1 gate8722(.O (I14855), .I1 (g9583), .I2 (g9593), .I3 (g9601), .I4 (g9596));
OR4X1 gate8723(.O (I15205), .I1 (g9838), .I2 (g9963), .I3 (g9850), .I4 (g9878));
OR4X1 gate8724(.O (I15051), .I1 (g7853), .I2 (g9673), .I3 (g9624), .I4 (g9785));
OR3X1 gate8725(.O (g9724), .I1 (g9409), .I2 (g9419), .I3 (g9615));
OR2X1 gate8726(.O (g6528), .I1 (g5756), .I2 (g4999));
OR2X1 gate8727(.O (g8823), .I1 (g8778), .I2 (g8693));
OR2X1 gate8728(.O (g7503), .I1 (g6887), .I2 (g6430));
OR2X1 gate8729(.O (g8148), .I1 (g7884), .I2 (g6872));
OR2X1 gate8730(.O (g8649), .I1 (g8499), .I2 (g4519));
OR2X1 gate8731(.O (g3584), .I1 (g2863), .I2 (g2516));
OR2X1 gate8732(.O (g10776), .I1 (g5544), .I2 (g10758));
OR3X1 gate8733(.O (g9680), .I1 (g9454), .I2 (g9292), .I3 (g9274));
OR2X1 gate8734(.O (g10859), .I1 (g5512), .I2 (g10742));
OR3X1 gate8735(.O (I14866), .I1 (g9590), .I2 (g9609), .I3 (g9619));
OR2X1 gate8736(.O (g7299), .I1 (g7138), .I2 (g6325));
OR2X1 gate8737(.O (g10858), .I1 (g5501), .I2 (g10741));
OR2X1 gate8738(.O (g8193), .I1 (g5145), .I2 (g7937));
OR3X1 gate8739(.O (g9511), .I1 (g9151), .I2 (g9125), .I3 (g9111));
OR2X1 gate8740(.O (g7738), .I1 (g7200), .I2 (g6738));
OR2X1 gate8741(.O (g7244), .I1 (g6699), .I2 (g4720));
OR2X1 gate8742(.O (g3425), .I1 (g2895), .I2 (g2910));
OR2X1 gate8743(.O (g7478), .I1 (g6884), .I2 (g6423));
OR3X1 gate8744(.O (g9714), .I1 (g9664), .I2 (g9366), .I3 (g9654));
OR2X1 gate8745(.O (g10025), .I1 (I15224), .I2 (I15225));
OR2X1 gate8746(.O (g6908), .I1 (g6345), .I2 (g4229));
OR2X1 gate8747(.O (g5028), .I1 (g4836), .I2 (g4128));
OR2X1 gate8748(.O (g8253), .I1 (g8023), .I2 (g7718));
OR2X1 gate8749(.O (g8938), .I1 (g8789), .I2 (g8699));
OR2X1 gate8750(.O (g8813), .I1 (g7943), .I2 (g8726));
OR2X1 gate8751(.O (g9736), .I1 (g9430), .I2 (g9416));
OR2X1 gate8752(.O (g9968), .I1 (I15171), .I2 (I15172));
OR2X1 gate8753(.O (g8552), .I1 (g8217), .I2 (g8388));
OR2X1 gate8754(.O (g5910), .I1 (g5023), .I2 (g4341));
OR2X1 gate8755(.O (g11249), .I1 (g6162), .I2 (g11143));
OR2X1 gate8756(.O (g11482), .I1 (g6628), .I2 (g11459));
OR4X1 gate8757(.O (g9722), .I1 (g9612), .I2 (g9643), .I3 (g9410), .I4 (I14855));
OR4X1 gate8758(.O (I15204), .I1 (g8168), .I2 (g9904), .I3 (g9933), .I4 (g9829));
OR2X1 gate8759(.O (g7236), .I1 (g6684), .I2 (g6092));
OR3X1 gate8760(.O (I14596), .I1 (g8995), .I2 (g9205), .I3 (g9192));
OR2X1 gate8761(.O (g8645), .I1 (g8127), .I2 (g8469));
OR2X1 gate8762(.O (g11647), .I1 (g6622), .I2 (g11637));
OR2X1 gate8763(.O (g6777), .I1 (g5691), .I2 (g5052));
OR3X1 gate8764(.O (g9737), .I1 (g9657), .I2 (g9658), .I3 (g9655));
OR4X1 gate8765(.O (I16149), .I1 (g10472), .I2 (g10470), .I3 (g10468), .I4 (g10467));
OR2X1 gate8766(.O (g11233), .I1 (g11085), .I2 (g10946));
OR2X1 gate8767(.O (g8607), .I1 (g8406), .I2 (g8554));
OR4X1 gate8768(.O (I16148), .I1 (g10386), .I2 (g10384), .I3 (g10476), .I4 (g10474));
OR2X1 gate8769(.O (g8158), .I1 (g7893), .I2 (g6883));
OR2X1 gate8770(.O (g5846), .I1 (g4932), .I2 (g4236));
OR2X1 gate8771(.O (g5396), .I1 (g4481), .I2 (g3684));
OR2X1 gate8772(.O (g5803), .I1 (g5575), .I2 (g4820));
OR2X1 gate8773(.O (g11331), .I1 (g11272), .I2 (g11171));
OR2X1 gate8774(.O (g7295), .I1 (g7071), .I2 (g6321));
OR2X1 gate8775(.O (g6541), .I1 (g5788), .I2 (g5009));
OR2X1 gate8776(.O (g8615), .I1 (g8413), .I2 (g8557));
OR2X1 gate8777(.O (g9742), .I1 (g9173), .I2 (g9528));
OR2X1 gate8778(.O (g9926), .I1 (g9868), .I2 (g9715));
OR2X1 gate8779(.O (g9754), .I1 (g9173), .I2 (g9511));
OR2X1 gate8780(.O (g8284), .I1 (g8102), .I2 (g7821));
OR2X1 gate8781(.O (g2204), .I1 (g1393), .I2 (g1394));
OR2X1 gate8782(.O (g7471), .I1 (g6880), .I2 (g6416));
OR2X1 gate8783(.O (g7242), .I1 (g6693), .I2 (g6098));
OR2X1 gate8784(.O (g5847), .I1 (g5626), .I2 (g4877));
OR2X1 gate8785(.O (g6901), .I1 (g6788), .I2 (g6247));
OR2X1 gate8786(.O (g8559), .I1 (g8380), .I2 (g4731));
OR3X1 gate8787(.O (g9729), .I1 (g9618), .I2 (g9357), .I3 (g9656));
OR2X1 gate8788(.O (g10860), .I1 (g5513), .I2 (g10743));
OR2X1 gate8789(.O (g9927), .I1 (g9869), .I2 (g9716));
OR2X1 gate8790(.O (g10497), .I1 (g5052), .I2 (g10396));
OR4X1 gate8791(.O (g9885), .I1 (g9739), .I2 (g9598), .I3 (g9662), .I4 (g9746));
OR4X1 gate8792(.O (g2528), .I1 (g861), .I2 (g857), .I3 (g853), .I4 (g849));
OR2X1 gate8793(.O (g11229), .I1 (g11154), .I2 (g11012));
OR2X1 gate8794(.O (g8973), .I1 (g8821), .I2 (g8735));
OR2X1 gate8795(.O (g10658), .I1 (g10595), .I2 (g7674));
OR2X1 gate8796(.O (g10339), .I1 (g10232), .I2 (g9556));
OR4X1 gate8797(.O (I5363), .I1 (g1149), .I2 (g1153), .I3 (g1157), .I4 (g1160));
OR2X1 gate8798(.O (g11310), .I1 (g11220), .I2 (g11100));
OR2X1 gate8799(.O (g6500), .I1 (g5725), .I2 (g4986));
OR2X1 gate8800(.O (g10855), .I1 (g6075), .I2 (g10736));
OR2X1 gate8801(.O (g9916), .I1 (g9855), .I2 (g9694));
OR2X1 gate8802(.O (g10411), .I1 (g10299), .I2 (g9529));
OR2X1 gate8803(.O (g11603), .I1 (g11582), .I2 (g11553));
OR4X1 gate8804(.O (I5357), .I1 (g1265), .I2 (g1260), .I3 (g1255), .I4 (g1250));
OR2X1 gate8805(.O (g9560), .I1 (g9052), .I2 (g9030));
OR2X1 gate8806(.O (g6672), .I1 (g5941), .I2 (g5259));
OR3X1 gate8807(.O (g9873), .I1 (g9623), .I2 (g9599), .I3 (g9758));
OR2X1 gate8808(.O (g6523), .I1 (g5745), .I2 (g4995));
OR2X1 gate8809(.O (g10707), .I1 (g5545), .I2 (g10686));
OR4X1 gate8810(.O (I5626), .I1 (g521), .I2 (g525), .I3 (g530), .I4 (g534));
OR2X1 gate8811(.O (g9579), .I1 (g9052), .I2 (g9030));
OR2X1 gate8812(.O (g7298), .I1 (g7136), .I2 (g6324));
OR2X1 gate8813(.O (g6551), .I1 (g5804), .I2 (g5031));
OR2X1 gate8814(.O (g6099), .I1 (g5273), .I2 (g4550));
OR2X1 gate8815(.O (g8282), .I1 (g8101), .I2 (g7819));
OR2X1 gate8816(.O (g9917), .I1 (g9856), .I2 (g9695));
OR4X1 gate8817(.O (I15057), .I1 (g7853), .I2 (g9680), .I3 (g9624), .I4 (g9785));
OR2X1 gate8818(.O (g7219), .I1 (g6661), .I2 (g6076));
OR2X1 gate8819(.O (g10019), .I1 (I15219), .I2 (I15220));
OR2X1 gate8820(.O (g5857), .I1 (g5418), .I2 (g4670));
OR4X1 gate8821(.O (g9725), .I1 (g9642), .I2 (g9659), .I3 (g9616), .I4 (I14862));
OR2X1 gate8822(.O (g11298), .I1 (g11212), .I2 (g11087));
OR2X1 gate8823(.O (g10402), .I1 (g10295), .I2 (g9554));
OR4X1 gate8824(.O (g2521), .I1 (g538), .I2 (g542), .I3 (g476), .I4 (I5626));
OR3X1 gate8825(.O (I14751), .I1 (g8995), .I2 (g9205), .I3 (g9192));
OR2X1 gate8826(.O (g10866), .I1 (g5539), .I2 (g10753));
OR2X1 gate8827(.O (g6534), .I1 (g5772), .I2 (g5003));
OR2X1 gate8828(.O (g11232), .I1 (g11158), .I2 (g11015));
OR3X1 gate8829(.O (g9706), .I1 (g9644), .I2 (g9386), .I3 (g9591));
OR2X1 gate8830(.O (g10001), .I1 (I15204), .I2 (I15205));
OR2X1 gate8831(.O (g8776), .I1 (g5510), .I2 (g8655));
OR2X1 gate8832(.O (g7225), .I1 (g6666), .I2 (g6079));
OR3X1 gate8833(.O (g9888), .I1 (g9648), .I2 (g9608), .I3 (g9757));
OR2X1 gate8834(.O (g11261), .I1 (g11238), .I2 (g11023));
OR3X1 gate8835(.O (g9956), .I1 (g9948), .I2 (g9942), .I3 (g9815));
OR2X1 gate8836(.O (g10923), .I1 (g10778), .I2 (g10715));
OR2X1 gate8837(.O (g8264), .I1 (g7879), .I2 (g3389));
OR2X1 gate8838(.O (g6513), .I1 (g5737), .I2 (g4991));
OR3X1 gate8839(.O (I14835), .I1 (g9621), .I2 (g9645), .I3 (g9588));
OR2X1 gate8840(.O (g8641), .I1 (g8120), .I2 (g8463));
OR3X1 gate8841(.O (g5361), .I1 (g4316), .I2 (g4093), .I3 (g126));
OR2X1 gate8842(.O (g11316), .I1 (g11226), .I2 (g11103));
OR4X1 gate8843(.O (I16161), .I1 (g10479), .I2 (g10478), .I3 (g10477), .I4 (g10475));
OR2X1 gate8844(.O (g6916), .I1 (g6348), .I2 (g5687));
OR2X1 gate8845(.O (g8777), .I1 (g5522), .I2 (g8659));
OR4X1 gate8846(.O (g2353), .I1 (g1403), .I2 (g1407), .I3 (g1411), .I4 (g1415));
OR2X1 gate8847(.O (g7510), .I1 (g7186), .I2 (g6730));
OR3X1 gate8848(.O (g9957), .I1 (g9949), .I2 (g9943), .I3 (g9776));
OR2X1 gate8849(.O (g2744), .I1 (I5804), .I2 (I5805));
OR2X1 gate8850(.O (g7245), .I1 (g6696), .I2 (g6102));
OR2X1 gate8851(.O (g7291), .I1 (g7050), .I2 (g6317));
OR2X1 gate8852(.O (g8611), .I1 (g8410), .I2 (g8556));
OR4X1 gate8853(.O (I15199), .I1 (g8167), .I2 (g9903), .I3 (g9932), .I4 (g9828));
OR2X1 gate8854(.O (g10550), .I1 (g4942), .I2 (g10450));
OR2X1 gate8855(.O (g11330), .I1 (g11304), .I2 (g11170));
OR2X1 gate8856(.O (g10721), .I1 (g10306), .I2 (g10669));
OR2X1 gate8857(.O (g8153), .I1 (g7888), .I2 (g6875));
OR2X1 gate8858(.O (g10773), .I1 (g5540), .I2 (g10685));
OR2X1 gate8859(.O (g3688), .I1 (g3144), .I2 (g2454));
OR4X1 gate8860(.O (I15225), .I1 (g9842), .I2 (g9967), .I3 (g9859), .I4 (g9881));
OR2X1 gate8861(.O (g6042), .I1 (g5535), .I2 (g3987));
OR2X1 gate8862(.O (g10655), .I1 (g10561), .I2 (g7389));
OR2X1 gate8863(.O (g11259), .I1 (g11236), .I2 (g11021));
OR2X1 gate8864(.O (g11225), .I1 (g11149), .I2 (g11009));
OR2X1 gate8865(.O (g5914), .I1 (g5029), .I2 (g4343));
OR2X1 gate8866(.O (g11258), .I1 (g11235), .I2 (g11020));
OR2X1 gate8867(.O (g6054), .I1 (g5199), .I2 (g4483));
OR3X1 gate8868(.O (g9728), .I1 (g9412), .I2 (g9422), .I3 (g9426));
OR3X1 gate8869(.O (g9730), .I1 (g9414), .I2 (g9425), .I3 (g9423));
OR2X1 gate8870(.O (g5820), .I1 (g5595), .I2 (g4834));
OR3X1 gate8871(.O (g8574), .I1 (g5679), .I2 (g7853), .I3 (g8465));
OR2X1 gate8872(.O (g11602), .I1 (g11581), .I2 (g11552));
OR2X1 gate8873(.O (g10502), .I1 (g4169), .I2 (g10365));
OR2X1 gate8874(.O (g10557), .I1 (g4123), .I2 (g10508));
OR4X1 gate8875(.O (I15171), .I1 (g8175), .I2 (g9909), .I3 (g9896), .I4 (g9835));
OR2X1 gate8876(.O (g11337), .I1 (g11282), .I2 (g11177));
OR2X1 gate8877(.O (g7465), .I1 (g6876), .I2 (g6410));
OR2X1 gate8878(.O (g8262), .I1 (g7970), .I2 (g7625));
OR2X1 gate8879(.O (g8889), .I1 (g8844), .I2 (g8756));
OR2X1 gate8880(.O (g7096), .I1 (g6544), .I2 (g5911));
OR2X1 gate8881(.O (g5995), .I1 (g5097), .I2 (g5099));
OR2X1 gate8882(.O (g8285), .I1 (g8104), .I2 (g7822));
OR2X1 gate8883(.O (g10791), .I1 (g6186), .I2 (g10762));
OR2X1 gate8884(.O (g2499), .I1 (I5570), .I2 (I5571));
OR3X1 gate8885(.O (I14607), .I1 (g8995), .I2 (g9205), .I3 (g9192));
OR2X1 gate8886(.O (g6049), .I1 (g5254), .I2 (g3718));
OR2X1 gate8887(.O (g9920), .I1 (g9860), .I2 (g9701));
OR2X1 gate8888(.O (g10556), .I1 (g4115), .I2 (g10506));
OR2X1 gate8889(.O (g8643), .I1 (g8364), .I2 (g8508));
OR2X1 gate8890(.O (g5810), .I1 (g5588), .I2 (g4823));
OR2X1 gate8891(.O (g11336), .I1 (g11281), .I2 (g11176));
OR2X1 gate8892(.O (g8742), .I1 (g8135), .I2 (g8598));
OR2X1 gate8893(.O (g8926), .I1 (g8848), .I2 (g8764));
OR2X1 gate8894(.O (g7218), .I1 (g6655), .I2 (g6070));
OR4X1 gate8895(.O (I15224), .I1 (g8174), .I2 (g9908), .I3 (g9937), .I4 (g9834));
OR2X1 gate8896(.O (g7293), .I1 (g7063), .I2 (g6319));
OR2X1 gate8897(.O (g11288), .I1 (g11204), .I2 (g11070));
OR2X1 gate8898(.O (g10800), .I1 (g6245), .I2 (g10772));
OR2X1 gate8899(.O (g11308), .I1 (g11218), .I2 (g11098));
OR2X1 gate8900(.O (g8269), .I1 (g7892), .I2 (g3429));
OR2X1 gate8901(.O (g10417), .I1 (g10301), .I2 (g9527));
OR2X1 gate8902(.O (g10936), .I1 (g5170), .I2 (g10808));
OR2X1 gate8903(.O (g9388), .I1 (g9240), .I2 (g9223));
OR2X1 gate8904(.O (g6185), .I1 (g5470), .I2 (g4715));
OR2X1 gate8905(.O (g6470), .I1 (g5699), .I2 (g4960));
OR2X1 gate8906(.O (g6897), .I1 (g6771), .I2 (g6240));
OR2X1 gate8907(.O (g8885), .I1 (g8841), .I2 (g8754));
OR2X1 gate8908(.O (g11260), .I1 (g11237), .I2 (g11022));
OR2X1 gate8909(.O (g11488), .I1 (g6671), .I2 (g11465));
OR2X1 gate8910(.O (g6105), .I1 (g5279), .I2 (g4559));
OR2X1 gate8911(.O (g10807), .I1 (g10701), .I2 (g10761));
OR2X1 gate8912(.O (g10639), .I1 (g10623), .I2 (g7734));
OR2X1 gate8913(.O (g4556), .I1 (g3536), .I2 (g2916));
OR2X1 gate8914(.O (g8288), .I1 (g8119), .I2 (g7825));
OR2X1 gate8915(.O (g6755), .I1 (g6106), .I2 (g5479));
OR3X1 gate8916(.O (I14862), .I1 (g9587), .I2 (g9600), .I3 (g9611));
OR4X1 gate8917(.O (I16160), .I1 (g10394), .I2 (g10392), .I3 (g10482), .I4 (g10481));
OR4X1 gate8918(.O (I15042), .I1 (g7853), .I2 (g9686), .I3 (g9624), .I4 (g9785));
OR2X1 gate8919(.O (g11610), .I1 (g11589), .I2 (g11560));
OR4X1 gate8920(.O (g9711), .I1 (g9660), .I2 (g9390), .I3 (g9359), .I4 (g9589));
OR2X1 gate8921(.O (g6045), .I1 (g5541), .I2 (g3989));
OR2X1 gate8922(.O (g11270), .I1 (g11198), .I2 (g11032));
OR2X1 gate8923(.O (g7258), .I1 (g6549), .I2 (g5913));
OR2X1 gate8924(.O (g6059), .I1 (g5211), .I2 (g4489));
OR2X1 gate8925(.O (g10007), .I1 (I15209), .I2 (I15210));
OR2X1 gate8926(.O (g11267), .I1 (g11192), .I2 (g11029));
OR2X1 gate8927(.O (g11294), .I1 (g6576), .I2 (g11210));
OR3X1 gate8928(.O (g9509), .I1 (g9151), .I2 (g9125), .I3 (g9111));
OR2X1 gate8929(.O (g7211), .I1 (g6647), .I2 (g6067));
OR2X1 gate8930(.O (g5404), .I1 (g4487), .I2 (g3696));
OR2X1 gate8931(.O (g4089), .I1 (g1959), .I2 (g3318));
OR4X1 gate8932(.O (I15219), .I1 (g8172), .I2 (g9907), .I3 (g9936), .I4 (g9833));
OR2X1 gate8933(.O (g11219), .I1 (g11145), .I2 (g11006));
OR2X1 gate8934(.O (g6015), .I1 (g5497), .I2 (g3942));
OR2X1 gate8935(.O (g10720), .I1 (g10304), .I2 (g10667));
OR2X1 gate8936(.O (g8265), .I1 (g7881), .I2 (g3396));
OR2X1 gate8937(.O (g5224), .I1 (g4360), .I2 (g3512));
OR3X1 gate8938(.O (g9700), .I1 (g9358), .I2 (g9667), .I3 (I14827));
OR2X1 gate8939(.O (g7106), .I1 (g6554), .I2 (g5917));
OR2X1 gate8940(.O (g8770), .I1 (g5476), .I2 (g8651));
OR2X1 gate8941(.O (g11201), .I1 (g11152), .I2 (g11011));
OR3X1 gate8942(.O (g9950), .I1 (g9901), .I2 (g9898), .I3 (g9779));
OR4X1 gate8943(.O (g9723), .I1 (g9620), .I2 (g9652), .I3 (g9391), .I4 (I14858));
OR2X1 gate8944(.O (g2309), .I1 (I5357), .I2 (I5358));
OR2X1 gate8945(.O (g11266), .I1 (g11190), .I2 (g11028));
OR2X1 gate8946(.O (g10727), .I1 (g4969), .I2 (g10638));
OR2X1 gate8947(.O (g10863), .I1 (g5531), .I2 (g10750));
OR2X1 gate8948(.O (g8429), .I1 (g8385), .I2 (g8069));
OR2X1 gate8949(.O (g9751), .I1 (g9515), .I2 (g9510));
OR2X1 gate8950(.O (g8281), .I1 (g8097), .I2 (g7818));
OR2X1 gate8951(.O (g6910), .I1 (g6341), .I2 (g5680));
OR2X1 gate8952(.O (g8639), .I1 (g8118), .I2 (g8462));
OR3X1 gate8953(.O (g9673), .I1 (g9454), .I2 (g9292), .I3 (g9274));
OR2X1 gate8954(.O (g11285), .I1 (g11255), .I2 (g11161));
OR2X1 gate8955(.O (g11305), .I1 (g11215), .I2 (g11093));
OR4X1 gate8956(.O (I15177), .I1 (g9844), .I2 (g9960), .I3 (g9863), .I4 (g9876));
OR3X1 gate8957(.O (g9734), .I1 (g9415), .I2 (g9428), .I3 (g9421));
OR3X1 gate8958(.O (I14827), .I1 (g9603), .I2 (g9614), .I3 (g9584));
OR2X1 gate8959(.O (g5824), .I1 (g5602), .I2 (g4839));
OR2X1 gate8960(.O (g8715), .I1 (g8416), .I2 (g8687));
OR2X1 gate8961(.O (g5762), .I1 (g5178), .I2 (g5186));
OR2X1 gate8962(.O (g6538), .I1 (g5782), .I2 (g5006));
OR2X1 gate8963(.O (g5590), .I1 (g4718), .I2 (g4723));
OR2X1 gate8964(.O (g10726), .I1 (g10316), .I2 (g10673));
OR2X1 gate8965(.O (g3120), .I1 (I6350), .I2 (I6351));
OR2X1 gate8966(.O (g9573), .I1 (g9052), .I2 (g9030));
OR3X1 gate8967(.O (g4640), .I1 (g3348), .I2 (g3563), .I3 (g1527));
OR2X1 gate8968(.O (g6093), .I1 (g5264), .I2 (g4534));
OR2X1 gate8969(.O (g8162), .I1 (g7898), .I2 (g6889));
OR2X1 gate8970(.O (g8268), .I1 (g7962), .I2 (g7613));
OR2X1 gate8971(.O (g9569), .I1 (g9052), .I2 (g9030));
OR2X1 gate8972(.O (g11485), .I1 (g6646), .I2 (g11462));
OR2X1 gate8973(.O (g10797), .I1 (g6206), .I2 (g10766));
OR3X1 gate8974(.O (I14779), .I1 (g8995), .I2 (g9205), .I3 (g9192));
OR2X1 gate8975(.O (g10408), .I1 (g10298), .I2 (g9553));
OR2X1 gate8976(.O (g10635), .I1 (g10622), .I2 (g7732));
OR2X1 gate8977(.O (g2305), .I1 (I5351), .I2 (I5352));
OR4X1 gate8978(.O (I15176), .I1 (g8176), .I2 (g9910), .I3 (g9897), .I4 (g9836));
OR2X1 gate8979(.O (g3435), .I1 (g2945), .I2 (g2950));
OR2X1 gate8980(.O (g9924), .I1 (g9866), .I2 (g9709));
OR2X1 gate8981(.O (g10711), .I1 (g5547), .I2 (g10690));
OR2X1 gate8982(.O (g5814), .I1 (g5591), .I2 (g4827));
OR2X1 gate8983(.O (g5038), .I1 (g4878), .I2 (g4884));
OR4X1 gate8984(.O (I15215), .I1 (g9840), .I2 (g9965), .I3 (g9854), .I4 (g9879));
OR2X1 gate8985(.O (g8226), .I1 (g7504), .I2 (g8002));
OR2X1 gate8986(.O (g7367), .I1 (g7224), .I2 (g6744));
OR2X1 gate8987(.O (g7457), .I1 (g6873), .I2 (g6404));
OR2X1 gate8988(.O (g5229), .I1 (g4364), .I2 (g3516));
OR2X1 gate8989(.O (g5993), .I1 (g5090), .I2 (g4400));
OR2X1 gate8990(.O (g8283), .I1 (g8098), .I2 (g7820));
OR2X1 gate8991(.O (g7971), .I1 (g5110), .I2 (g7549));
OR2X1 gate8992(.O (g8602), .I1 (g8401), .I2 (g8550));
OR2X1 gate8993(.O (g8920), .I1 (g8845), .I2 (g8759));
OR2X1 gate8994(.O (g10663), .I1 (g10237), .I2 (g10581));
OR2X1 gate8995(.O (g6074), .I1 (g5349), .I2 (g1));
OR2X1 gate8996(.O (g8261), .I1 (g7876), .I2 (g3383));
OR2X1 gate8997(.O (g10862), .I1 (g5524), .I2 (g10746));
OR2X1 gate8998(.O (g5837), .I1 (g5640), .I2 (g4224));
OR2X1 gate8999(.O (g11333), .I1 (g11274), .I2 (g11173));
OR2X1 gate9000(.O (g6080), .I1 (g5249), .I2 (g4512));
OR2X1 gate9001(.O (g6480), .I1 (g5721), .I2 (g4971));
OR2X1 gate9002(.O (g7740), .I1 (g7209), .I2 (g6741));
OR2X1 gate9003(.O (g10702), .I1 (g10562), .I2 (g3877));
OR3X1 gate9004(.O (g9697), .I1 (g9665), .I2 (g9606), .I3 (I14822));
OR2X1 gate9005(.O (g8203), .I1 (g7453), .I2 (g7999));
OR2X1 gate9006(.O (g9914), .I1 (g9851), .I2 (g9692));
OR2X1 gate9007(.O (g10564), .I1 (g10560), .I2 (g7368));
OR2X1 gate9008(.O (g11484), .I1 (g6639), .I2 (g11461));
OR2X1 gate9009(.O (g5842), .I1 (g5618), .I2 (g4870));
OR4X1 gate9010(.O (I15200), .I1 (g9837), .I2 (g9962), .I3 (g9848), .I4 (g9880));
OR2X1 gate9011(.O (g11609), .I1 (g11588), .I2 (g11559));
OR3X1 gate9012(.O (I14582), .I1 (g8995), .I2 (g9205), .I3 (g9192));
OR2X1 gate9013(.O (g8940), .I1 (g8793), .I2 (g8703));
OR2X1 gate9014(.O (g11312), .I1 (g11222), .I2 (g11101));
OR2X1 gate9015(.O (g11608), .I1 (g11587), .I2 (g11558));
OR2X1 gate9016(.O (g6000), .I1 (g5480), .I2 (g3912));
OR2X1 gate9017(.O (g8428), .I1 (g8382), .I2 (g8068));
OR2X1 gate9018(.O (g8430), .I1 (g8386), .I2 (g8070));
OR2X1 gate9019(.O (g9922), .I1 (g9864), .I2 (g9705));
OR2X1 gate9020(.O (g8247), .I1 (g8010), .I2 (g7704));
OR2X1 gate9021(.O (g3438), .I1 (g2939), .I2 (g2944));
OR4X1 gate9022(.O (I5576), .I1 (g431), .I2 (g435), .I3 (g440), .I4 (g444));
OR2X1 gate9023(.O (g6924), .I1 (g6362), .I2 (g4261));
OR2X1 gate9024(.O (g5405), .I1 (g4476), .I2 (g3440));
OR2X1 gate9025(.O (g8638), .I1 (g8108), .I2 (g8461));
OR2X1 gate9026(.O (g8609), .I1 (g8408), .I2 (g8555));
OR2X1 gate9027(.O (g9995), .I1 (I15199), .I2 (I15200));
OR2X1 gate9028(.O (g8883), .I1 (g8838), .I2 (g8753));
OR4X1 gate9029(.O (I15214), .I1 (g8170), .I2 (g9906), .I3 (g9935), .I4 (g9831));
OR3X1 gate9030(.O (g2538), .I1 (g1466), .I2 (g1458), .I3 (I5649));
OR2X1 gate9031(.O (g11329), .I1 (g11302), .I2 (g11169));
OR2X1 gate9032(.O (g4255), .I1 (g4009), .I2 (g4047));
OR2X1 gate9033(.O (g11328), .I1 (g11299), .I2 (g11168));
OR3X1 gate9034(.O (g9704), .I1 (g9385), .I2 (g9605), .I3 (I14835));
OR4X1 gate9035(.O (I5352), .I1 (g1129), .I2 (g1125), .I3 (g1121), .I4 (g1117));
OR2X1 gate9036(.O (g8774), .I1 (g5499), .I2 (g8654));
OR3X1 gate9037(.O (g9954), .I1 (g9946), .I2 (g9940), .I3 (g9781));
OR2X1 gate9038(.O (g10405), .I1 (g10297), .I2 (g9530));
OR2X1 gate9039(.O (g9363), .I1 (g9205), .I2 (g9192));
OR2X1 gate9040(.O (g5849), .I1 (g4949), .I2 (g4260));
OR4X1 gate9041(.O (I5599), .I1 (g516), .I2 (g511), .I3 (g506), .I4 (g501));
OR2X1 gate9042(.O (g7204), .I1 (g6645), .I2 (g6062));
OR2X1 gate9043(.O (g7300), .I1 (g7139), .I2 (g6326));
OR2X1 gate9044(.O (g4293), .I1 (g4064), .I2 (g4068));
OR2X1 gate9045(.O (g9912), .I1 (g9847), .I2 (g9690));
OR2X1 gate9046(.O (g6533), .I1 (g5771), .I2 (g5002));
OR2X1 gate9047(.O (g8816), .I1 (g7951), .I2 (g8731));
OR2X1 gate9048(.O (g9929), .I1 (g9871), .I2 (g9718));
OR2X1 gate9049(.O (g5819), .I1 (g5625), .I2 (g4876));
OR3X1 gate9050(.O (I14831), .I1 (g9613), .I2 (g9622), .I3 (g9586));
OR2X1 gate9051(.O (g5852), .I1 (g5632), .I2 (g4883));
OR2X1 gate9052(.O (g8263), .I1 (g8032), .I2 (g7720));
OR2X1 gate9053(.O (g3431), .I1 (g2951), .I2 (g2957));
OR3X1 gate9054(.O (g9683), .I1 (g9454), .I2 (g9292), .I3 (g9274));
OR2X1 gate9055(.O (g8631), .I1 (g8474), .I2 (g7449));
OR2X1 gate9056(.O (g6922), .I1 (g6352), .I2 (g5694));
OR2X1 gate9057(.O (g8817), .I1 (g7954), .I2 (g8732));
OR4X1 gate9058(.O (g9735), .I1 (g9649), .I2 (g9651), .I3 (g9384), .I4 (g9361));
OR2X1 gate9059(.O (g8605), .I1 (g8404), .I2 (g8553));
OR2X1 gate9060(.O (g11263), .I1 (g11187), .I2 (g11025));
OR2X1 gate9061(.O (g6739), .I1 (g5769), .I2 (g5780));
OR2X1 gate9062(.O (g11332), .I1 (g11273), .I2 (g11172));
OR2X1 gate9063(.O (g7143), .I1 (g6619), .I2 (g6039));
OR2X1 gate9064(.O (g6479), .I1 (g5707), .I2 (g4968));
OR4X1 gate9065(.O (I15048), .I1 (g7853), .I2 (g9683), .I3 (g9624), .I4 (g9785));
OR2X1 gate9066(.O (g6501), .I1 (g5726), .I2 (g4987));
OR3X1 gate9067(.O (g9702), .I1 (g9365), .I2 (g9647), .I3 (I14831));
OR2X1 gate9068(.O (g11221), .I1 (g11146), .I2 (g11007));
OR3X1 gate9069(.O (g9952), .I1 (g9944), .I2 (g9938), .I3 (g9817));
OR2X1 gate9070(.O (g11613), .I1 (g11600), .I2 (g11591));
OR2X1 gate9071(.O (g7621), .I1 (g5108), .I2 (g6994));
OR2X1 gate9072(.O (g3399), .I1 (g2918), .I2 (g2940));
OR2X1 gate9073(.O (g11605), .I1 (g11584), .I2 (g11555));
OR2X1 gate9074(.O (g4274), .I1 (g4054), .I2 (g4058));
OR3X1 gate9075(.O (I14602), .I1 (g8995), .I2 (g9205), .I3 (g9192));
OR4X1 gate9076(.O (I15033), .I1 (g7853), .I2 (g9804), .I3 (g9624), .I4 (g9785));
OR2X1 gate9077(.O (g10717), .I1 (g6235), .I2 (g10705));
OR3X1 gate9078(.O (I5629), .I1 (g845), .I2 (g841), .I3 (g837));
OR2X1 gate9079(.O (g9925), .I1 (g9867), .I2 (g9712));
OR2X1 gate9080(.O (g3819), .I1 (g3275), .I2 (g9));
OR2X1 gate9081(.O (g6912), .I1 (g6350), .I2 (g4235));
OR2X1 gate9082(.O (g10723), .I1 (g4952), .I2 (g10633));
OR2X1 gate9083(.O (g6929), .I1 (g6360), .I2 (g5704));
OR2X1 gate9084(.O (g10646), .I1 (g10625), .I2 (g7739));
OR2X1 gate9085(.O (g9516), .I1 (g9151), .I2 (g9125));
OR2X1 gate9086(.O (g6626), .I1 (g5934), .I2 (g123));
OR4X1 gate9087(.O (I6350), .I1 (g2445), .I2 (g2437), .I3 (g2433), .I4 (g2419));
OR2X1 gate9088(.O (g11325), .I1 (g11295), .I2 (g11165));
OR4X1 gate9089(.O (I5366), .I1 (g1280), .I2 (g1284), .I3 (g1292), .I4 (g1296));
OR3X1 gate9090(.O (I5649), .I1 (g1499), .I2 (g1486), .I3 (g1482));
OR2X1 gate9091(.O (g6894), .I1 (g6763), .I2 (g4868));
OR3X1 gate9092(.O (g9738), .I1 (g9417), .I2 (g9447), .I3 (g9506));
OR2X1 gate9093(.O (g8383), .I1 (g8163), .I2 (g5051));
OR2X1 gate9094(.O (g8779), .I1 (g5530), .I2 (g8663));
OR2X1 gate9095(.O (g8161), .I1 (g8005), .I2 (g7185));
OR2X1 gate9096(.O (g8451), .I1 (g3440), .I2 (g8366));
OR2X1 gate9097(.O (g9915), .I1 (g9853), .I2 (g9693));
OR4X1 gate9098(.O (g2316), .I1 (g1300), .I2 (g1304), .I3 (g1270), .I4 (I5366));
OR2X1 gate9099(.O (g5576), .I1 (g4675), .I2 (g3664));
OR2X1 gate9100(.O (g10857), .I1 (g6090), .I2 (g10738));
OR2X1 gate9101(.O (g10793), .I1 (g6194), .I2 (g10763));
OR2X1 gate9102(.O (g7511), .I1 (g6890), .I2 (g6438));
OR2X1 gate9103(.O (g8944), .I1 (g8799), .I2 (g8708));
OR2X1 gate9104(.O (g10765), .I1 (g5492), .I2 (g10680));
OR2X1 gate9105(.O (g10549), .I1 (g4951), .I2 (g10451));
OR2X1 gate9106(.O (g7092), .I1 (g6540), .I2 (g5902));
OR2X1 gate9107(.O (g11604), .I1 (g11583), .I2 (g11554));
OR2X1 gate9108(.O (g8434), .I1 (g8400), .I2 (g8074));
OR2X1 gate9109(.O (g6546), .I1 (g5796), .I2 (g5026));
OR2X1 gate9110(.O (g3354), .I1 (g2920), .I2 (g2124));
OR2X1 gate9111(.O (g9928), .I1 (g9870), .I2 (g9717));
OR2X1 gate9112(.O (g11262), .I1 (g11240), .I2 (g11024));
OR4X1 gate9113(.O (g9785), .I1 (g9010), .I2 (g8995), .I3 (g9388), .I4 (g9363));
OR2X1 gate9114(.O (g5867), .I1 (g3440), .I2 (g4921));
OR2X1 gate9115(.O (g8210), .I1 (g7466), .I2 (g7995));
OR2X1 gate9116(.O (g10533), .I1 (g4933), .I2 (g10449));
OR2X1 gate9117(.O (g9563), .I1 (g9052), .I2 (g9030));
OR2X1 gate9118(.O (g6906), .I1 (g6791), .I2 (g5674));
OR2X1 gate9119(.O (g7375), .I1 (g7230), .I2 (g6745));
OR2X1 gate9120(.O (g7651), .I1 (g7135), .I2 (g4084));
OR4X1 gate9121(.O (I5570), .I1 (g416), .I2 (g411), .I3 (g406), .I4 (g401));
OR3X1 gate9122(.O (g9731), .I1 (g9641), .I2 (g9364), .I3 (g9387));
OR2X1 gate9123(.O (g11247), .I1 (g11097), .I2 (g10949));
OR4X1 gate9124(.O (I15045), .I1 (g7853), .I2 (g9676), .I3 (g9624), .I4 (g9785));
OR2X1 gate9125(.O (g10856), .I1 (g6083), .I2 (g10737));
OR2X1 gate9126(.O (g9557), .I1 (g9052), .I2 (g9030));
OR2X1 gate9127(.O (g7184), .I1 (g6625), .I2 (g6047));
OR2X1 gate9128(.O (g11612), .I1 (g11599), .I2 (g11590));
OR2X1 gate9129(.O (g7384), .I1 (g7088), .I2 (g6618));
OR2X1 gate9130(.O (g11324), .I1 (g11271), .I2 (g11164));
OR2X1 gate9131(.O (g8922), .I1 (g8822), .I2 (g8736));
OR4X1 gate9132(.O (I5358), .I1 (g1245), .I2 (g1240), .I3 (g1235), .I4 (g1275));
OR3X1 gate9133(.O (g9955), .I1 (g9947), .I2 (g9941), .I3 (g9808));
OR4X1 gate9134(.O (g2501), .I1 (g448), .I2 (g452), .I3 (g421), .I4 (I5576));
OR2X1 gate9135(.O (g7231), .I1 (g6673), .I2 (g6087));
OR2X1 gate9136(.O (g6078), .I1 (g4503), .I2 (g5256));
OR2X1 gate9137(.O (g6478), .I1 (g5706), .I2 (g4967));
OR2X1 gate9138(.O (g6907), .I1 (g6792), .I2 (g5675));
OR2X1 gate9139(.O (g6035), .I1 (g5518), .I2 (g3974));
OR2X1 gate9140(.O (g8937), .I1 (g8786), .I2 (g8698));
OR2X1 gate9141(.O (g7742), .I1 (g7217), .I2 (g6743));
OR2X1 gate9142(.O (g10722), .I1 (g10308), .I2 (g10671));
OR2X1 gate9143(.O (g9918), .I1 (g9858), .I2 (g9698));
OR2X1 gate9144(.O (g5403), .I1 (g4486), .I2 (g3695));
OR2X1 gate9145(.O (g7926), .I1 (g7435), .I2 (g6892));
OR2X1 gate9146(.O (g6915), .I1 (g6347), .I2 (g5686));
OR2X1 gate9147(.O (g5841), .I1 (g4914), .I2 (g4230));
OR4X1 gate9148(.O (I15220), .I1 (g9841), .I2 (g9966), .I3 (g9857), .I4 (g9877));
OR2X1 gate9149(.O (g10529), .I1 (I16160), .I2 (I16161));
OR2X1 gate9150(.O (g11246), .I1 (g11094), .I2 (g10948));
OR2X1 gate9151(.O (g6002), .I1 (g5489), .I2 (g3939));
OR2X1 gate9152(.O (g7712), .I1 (g7125), .I2 (g3540));
OR2X1 gate9153(.O (g8810), .I1 (g7933), .I2 (g8720));
OR2X1 gate9154(.O (g9921), .I1 (g9862), .I2 (g9703));
OR2X1 gate9155(.O (g8432), .I1 (g8389), .I2 (g8072));
OR4X1 gate9156(.O (I15172), .I1 (g9843), .I2 (g9959), .I3 (g9861), .I4 (g9874));
OR3X1 gate9157(.O (I14822), .I1 (g9597), .I2 (g9604), .I3 (g9582));
OR2X1 gate9158(.O (g6928), .I1 (g6359), .I2 (g5703));
OR2X1 gate9159(.O (g8157), .I1 (g7965), .I2 (g7623));
OR2X1 gate9160(.O (g6930), .I1 (g6364), .I2 (g4269));
OR2X1 gate9161(.O (g7660), .I1 (g7059), .I2 (g6583));
OR2X1 gate9162(.O (g6899), .I1 (g6463), .I2 (g5471));
OR2X1 gate9163(.O (g9392), .I1 (g9328), .I2 (g9324));
OR2X1 gate9164(.O (g11318), .I1 (g11228), .I2 (g11104));
OR3X1 gate9165(.O (I16427), .I1 (g10683), .I2 (g10608), .I3 (g10604));
OR2X1 gate9166(.O (g11227), .I1 (g11151), .I2 (g11010));
OR2X1 gate9167(.O (g11058), .I1 (g10933), .I2 (g5280));
OR4X1 gate9168(.O (I5351), .I1 (g1145), .I2 (g1141), .I3 (g1137), .I4 (g1133));
OR3X1 gate9169(.O (g9708), .I1 (g9653), .I2 (g9389), .I3 (g9646));
OR2X1 gate9170(.O (g6071), .I1 (g5228), .I2 (g4505));
OR2X1 gate9171(.O (g9911), .I1 (g9846), .I2 (g9689));
OR2X1 gate9172(.O (g7102), .I1 (g6550), .I2 (g5915));
OR2X1 gate9173(.O (g7302), .I1 (g7141), .I2 (g6328));
OR2X1 gate9174(.O (g6038), .I1 (g5528), .I2 (g3979));
OR2X1 gate9175(.O (g4239), .I1 (g4000), .I2 (g4008));
OR2X1 gate9176(.O (g8646), .I1 (g8224), .I2 (g8547));
OR2X1 gate9177(.O (g9974), .I1 (I15176), .I2 (I15177));
OR2X1 gate9178(.O (g5823), .I1 (g5631), .I2 (g4882));
OR2X1 gate9179(.O (g6918), .I1 (g6358), .I2 (g4252));
OR2X1 gate9180(.O (g7265), .I1 (g6756), .I2 (g6204));
OR4X1 gate9181(.O (I5804), .I1 (g2111), .I2 (g2109), .I3 (g2106), .I4 (g2104));
OR2X1 gate9182(.O (g5851), .I1 (g4941), .I2 (g4253));
OR2X1 gate9183(.O (g11481), .I1 (g6624), .I2 (g11458));
OR2X1 gate9184(.O (g10336), .I1 (g10230), .I2 (g9572));
OR2X1 gate9185(.O (g7296), .I1 (g7131), .I2 (g6322));
OR2X1 gate9186(.O (g4300), .I1 (g3546), .I2 (g2391));
OR2X1 gate9187(.O (g8647), .I1 (g8130), .I2 (g8470));
ND2X1 gate9188(.O (g8546), .I1 (g3983), .I2 (g8390));
ND2X1 gate9189(.O (g2516), .I1 (I5612), .I2 (I5613));
ND2X1 gate9190(.O (g2987), .I1 (g2481), .I2 (g883));
ND2X1 gate9191(.O (I5593), .I1 (g1703), .I2 (I5591));
ND2X1 gate9192(.O (g8970), .I1 (g5548), .I2 (g8839));
ND2X1 gate9193(.O (I10519), .I1 (g6231), .I2 (g822));
ND2X1 gate9194(.O (I11279), .I1 (g305), .I2 (I11278));
ND4X1 gate9195(.O (g7990), .I1 (g7011), .I2 (g6995), .I3 (g7562), .I4 (g7550));
ND2X1 gate9196(.O (I11278), .I1 (g305), .I2 (g6485));
ND2X1 gate9197(.O (g3978), .I1 (g3207), .I2 (g1822));
ND2X1 gate9198(.O (I5264), .I1 (g456), .I2 (I5263));
ND2X1 gate9199(.O (I8640), .I1 (g4278), .I2 (g516));
ND2X1 gate9200(.O (I6761), .I1 (g2943), .I2 (I6760));
ND2X1 gate9201(.O (I17400), .I1 (g11418), .I2 (g11416));
ND2X1 gate9202(.O (I5450), .I1 (g1235), .I2 (I5449));
ND2X1 gate9203(.O (I16060), .I1 (g10372), .I2 (I16058));
ND2X1 gate9204(.O (I6746), .I1 (g2938), .I2 (g1453));
ND2X1 gate9205(.O (I11975), .I1 (g1462), .I2 (I11973));
ND2X1 gate9206(.O (I12136), .I1 (g7110), .I2 (g131));
ND2X1 gate9207(.O (I11937), .I1 (g1458), .I2 (I11935));
ND2X1 gate9208(.O (g2959), .I1 (I6167), .I2 (I6168));
ND2X1 gate9209(.O (I5878), .I1 (g2120), .I2 (g2115));
ND2X1 gate9210(.O (g2517), .I1 (I5619), .I2 (I5620));
ND2X1 gate9211(.O (g5552), .I1 (g4777), .I2 (g4401));
ND2X1 gate9212(.O (I6468), .I1 (g23), .I2 (I6467));
ND2X1 gate9213(.O (I8796), .I1 (g4672), .I2 (I8795));
ND2X1 gate9214(.O (g10392), .I1 (I15891), .I2 (I15892));
ND2X1 gate9215(.O (I5611), .I1 (g1280), .I2 (g1284));
ND2X1 gate9216(.O (g8738), .I1 (g8688), .I2 (g4921));
ND2X1 gate9217(.O (I6716), .I1 (g201), .I2 (I6714));
ND2X1 gate9218(.O (g2310), .I1 (g591), .I2 (g605));
ND2X1 gate9219(.O (I7685), .I1 (g3460), .I2 (I7683));
ND2X1 gate9220(.O (g3056), .I1 (g2374), .I2 (g599));
ND2X1 gate9221(.O (I12108), .I1 (g135), .I2 (I12106));
ND3X1 gate9222(.O (g3529), .I1 (g2310), .I2 (g3062), .I3 (g2325));
ND2X1 gate9223(.O (I6747), .I1 (g2938), .I2 (I6746));
ND2X1 gate9224(.O (g2236), .I1 (I5230), .I2 (I5231));
ND2X1 gate9225(.O (g7584), .I1 (I12075), .I2 (I12076));
ND2X1 gate9226(.O (I15870), .I1 (g10358), .I2 (g2713));
ND2X1 gate9227(.O (I16067), .I1 (g2765), .I2 (I16065));
ND2X1 gate9228(.O (I7562), .I1 (g3533), .I2 (g654));
ND2X1 gate9229(.O (I13531), .I1 (g8253), .I2 (I13529));
ND2X1 gate9230(.O (I8797), .I1 (g1145), .I2 (I8795));
ND2X1 gate9231(.O (I17584), .I1 (g11354), .I2 (g11515));
ND2X1 gate9232(.O (I11936), .I1 (g7004), .I2 (I11935));
ND2X1 gate9233(.O (I15257), .I1 (g9984), .I2 (I15256));
ND2X1 gate9234(.O (g8402), .I1 (I13505), .I2 (I13506));
ND3X1 gate9235(.O (g8824), .I1 (g8502), .I2 (g8501), .I3 (g8739));
ND2X1 gate9236(.O (I6186), .I1 (g2511), .I2 (g466));
ND2X1 gate9237(.O (g11496), .I1 (I17504), .I2 (I17505));
ND2X1 gate9238(.O (I16001), .I1 (g2683), .I2 (I15999));
ND2X1 gate9239(.O (I6125), .I1 (g2215), .I2 (I6124));
ND2X1 gate9240(.O (I11909), .I1 (g1474), .I2 (I11907));
ND2X1 gate9241(.O (I12040), .I1 (g1466), .I2 (I12038));
ND2X1 gate9242(.O (I13909), .I1 (g1432), .I2 (I13907));
ND2X1 gate9243(.O (g3625), .I1 (I6771), .I2 (I6772));
ND2X1 gate9244(.O (I11908), .I1 (g6967), .I2 (I11907));
ND2X1 gate9245(.O (g10470), .I1 (I16008), .I2 (I16009));
ND2X1 gate9246(.O (I13908), .I1 (g8526), .I2 (I13907));
ND2X1 gate9247(.O (g3813), .I1 (I7034), .I2 (I7035));
ND2X1 gate9248(.O (I8650), .I1 (g4824), .I2 (g778));
ND2X1 gate9249(.O (g6207), .I1 (I9947), .I2 (I9948));
ND2X1 gate9250(.O (I16066), .I1 (g10428), .I2 (I16065));
ND2X1 gate9251(.O (g2948), .I1 (I6144), .I2 (I6145));
ND2X1 gate9252(.O (I11242), .I1 (g6760), .I2 (I11241));
ND2X1 gate9253(.O (g10467), .I1 (I15993), .I2 (I15994));
ND2X1 gate9254(.O (I6187), .I1 (g2511), .I2 (I6186));
ND2X1 gate9255(.O (g6488), .I1 (g6027), .I2 (g6019));
ND2X1 gate9256(.O (I5500), .I1 (g1255), .I2 (g1007));
ND2X1 gate9257(.O (I11974), .I1 (g7001), .I2 (I11973));
ND2X1 gate9258(.O (I12062), .I1 (g1478), .I2 (I12060));
ND2X1 gate9259(.O (g5300), .I1 (I8771), .I2 (I8772));
ND2X1 gate9260(.O (I5184), .I1 (g1415), .I2 (g1515));
ND2X1 gate9261(.O (I13293), .I1 (g1882), .I2 (g8161));
ND2X1 gate9262(.O (I6200), .I1 (g2525), .I2 (I6199));
ND2X1 gate9263(.O (I13265), .I1 (g1909), .I2 (g8154));
ND2X1 gate9264(.O (I5024), .I1 (g995), .I2 (I5023));
ND2X1 gate9265(.O (I7863), .I1 (g4099), .I2 (g774));
ND2X1 gate9266(.O (g8705), .I1 (I13991), .I2 (I13992));
ND2X1 gate9267(.O (g8471), .I1 (I13660), .I2 (I13661));
ND2X1 gate9268(.O (I15256), .I1 (g9984), .I2 (g9980));
ND2X1 gate9269(.O (I6145), .I1 (g646), .I2 (I6143));
ND2X1 gate9270(.O (I13992), .I1 (g8688), .I2 (I13990));
ND2X1 gate9271(.O (I11510), .I1 (g1806), .I2 (I11508));
ND2X1 gate9272(.O (g10853), .I1 (g10731), .I2 (g5034));
ND2X1 gate9273(.O (I5231), .I1 (g148), .I2 (I5229));
ND2X1 gate9274(.O (I12047), .I1 (g1486), .I2 (I12045));
ND2X1 gate9275(.O (I10771), .I1 (g1801), .I2 (I10769));
ND2X1 gate9276(.O (g10477), .I1 (I16045), .I2 (I16046));
ND2X1 gate9277(.O (g7582), .I1 (I12061), .I2 (I12062));
ND2X1 gate9278(.O (I5104), .I1 (g431), .I2 (g435));
ND2X1 gate9279(.O (g8409), .I1 (I13530), .I2 (I13531));
ND2X1 gate9280(.O (I6447), .I1 (g2264), .I2 (g1776));
ND2X1 gate9281(.O (I4956), .I1 (g327), .I2 (I4954));
ND2X1 gate9282(.O (I5613), .I1 (g1284), .I2 (I5611));
ND2X1 gate9283(.O (I8481), .I1 (g3530), .I2 (I8479));
ND2X1 gate9284(.O (g5278), .I1 (I8739), .I2 (I8740));
ND2X1 gate9285(.O (I6880), .I1 (g3301), .I2 (I6879));
ND2X1 gate9286(.O (I15431), .I1 (g10047), .I2 (I15430));
ND2X1 gate9287(.O (g5548), .I1 (g1840), .I2 (g4401));
ND4X1 gate9288(.O (g7671), .I1 (g7011), .I2 (g6995), .I3 (g6984), .I4 (g6974));
ND2X1 gate9289(.O (I12020), .I1 (g7119), .I2 (I12019));
ND2X1 gate9290(.O (g10665), .I1 (I16331), .I2 (I16332));
ND2X1 gate9291(.O (I16469), .I1 (g10518), .I2 (I16467));
ND2X1 gate9292(.O (I5014), .I1 (g1007), .I2 (I5013));
ND2X1 gate9293(.O (I13523), .I1 (g8249), .I2 (I13521));
ND2X1 gate9294(.O (I16039), .I1 (g2707), .I2 (I16037));
ND2X1 gate9295(.O (I16468), .I1 (g10716), .I2 (I16467));
ND2X1 gate9296(.O (I12046), .I1 (g6951), .I2 (I12045));
ND2X1 gate9297(.O (g4476), .I1 (g3807), .I2 (g3071));
ND2X1 gate9298(.O (g10476), .I1 (I16038), .I2 (I16039));
ND2X1 gate9299(.O (I16038), .I1 (g10427), .I2 (I16037));
ND2X1 gate9300(.O (I8676), .I1 (g4374), .I2 (g1027));
ND2X1 gate9301(.O (I12113), .I1 (g7093), .I2 (g162));
ND2X1 gate9302(.O (I8761), .I1 (g4616), .I2 (g1129));
ND2X1 gate9303(.O (g3204), .I1 (g2571), .I2 (g2061));
ND2X1 gate9304(.O (I15993), .I1 (g10422), .I2 (I15992));
ND2X1 gate9305(.O (I5036), .I1 (g1019), .I2 (I5034));
ND2X1 gate9306(.O (I14263), .I1 (g8843), .I2 (g1814));
ND2X1 gate9307(.O (g8298), .I1 (I13249), .I2 (I13250));
ND2X1 gate9308(.O (I5135), .I1 (g521), .I2 (g525));
ND2X1 gate9309(.O (g2405), .I1 (I5485), .I2 (I5486));
ND2X1 gate9310(.O (I7034), .I1 (g3089), .I2 (I7033));
ND2X1 gate9311(.O (I15443), .I1 (g10122), .I2 (I15441));
ND2X1 gate9312(.O (I6166), .I1 (g2236), .I2 (g153));
ND2X1 gate9313(.O (I8624), .I1 (g4267), .I2 (g511));
ND2X1 gate9314(.O (I16015), .I1 (g10425), .I2 (g2695));
ND2X1 gate9315(.O (I8677), .I1 (g4374), .I2 (I8676));
ND2X1 gate9316(.O (I8576), .I1 (g4234), .I2 (I8575));
ND2X1 gate9317(.O (I14613), .I1 (g9204), .I2 (I14612));
ND2X1 gate9318(.O (I8716), .I1 (g4601), .I2 (I8715));
ND2X1 gate9319(.O (g3530), .I1 (I6715), .I2 (I6716));
ND2X1 gate9320(.O (g8405), .I1 (I13514), .I2 (I13515));
ND4X1 gate9321(.O (g4104), .I1 (g3215), .I2 (g3247), .I3 (g2439), .I4 (g3200));
ND2X1 gate9322(.O (I12003), .I1 (g7082), .I2 (I12002));
ND2X1 gate9323(.O (g2177), .I1 (I5127), .I2 (I5128));
ND2X1 gate9324(.O (g3010), .I1 (g2382), .I2 (g2399));
ND2X1 gate9325(.O (g5179), .I1 (I8576), .I2 (I8577));
ND2X1 gate9326(.O (I17395), .I1 (g11414), .I2 (I17393));
ND2X1 gate9327(.O (g7067), .I1 (I11279), .I2 (I11280));
ND4X1 gate9328(.O (g7994), .I1 (g7011), .I2 (g7574), .I3 (g6984), .I4 (g7550));
ND2X1 gate9329(.O (I6167), .I1 (g2236), .I2 (I6166));
ND2X1 gate9330(.O (I5265), .I1 (g461), .I2 (I5263));
ND2X1 gate9331(.O (I6989), .I1 (g2760), .I2 (I6988));
ND2X1 gate9332(.O (I13274), .I1 (g8158), .I2 (I13272));
ND2X1 gate9333(.O (I10507), .I1 (g6221), .I2 (g786));
ND2X1 gate9334(.O (I13530), .I1 (g704), .I2 (I13529));
ND2X1 gate9335(.O (I5164), .I1 (g1508), .I2 (g1499));
ND2X1 gate9336(.O (g9107), .I1 (I14443), .I2 (I14444));
ND2X1 gate9337(.O (I9559), .I1 (g782), .I2 (I9557));
ND2X1 gate9338(.O (I8577), .I1 (g496), .I2 (I8575));
ND2X1 gate9339(.O (g2510), .I1 (I5592), .I2 (I5593));
ND2X1 gate9340(.O (g8177), .I1 (I13077), .I2 (I13078));
ND2X1 gate9341(.O (I8717), .I1 (g4052), .I2 (I8715));
ND2X1 gate9342(.O (I5296), .I1 (g794), .I2 (I5295));
ND2X1 gate9343(.O (g5209), .I1 (I8625), .I2 (I8626));
ND4X1 gate9344(.O (g7950), .I1 (g7395), .I2 (g7390), .I3 (g7380), .I4 (g7273));
ND2X1 gate9345(.O (g2088), .I1 (I4911), .I2 (I4912));
ND2X1 gate9346(.O (I16000), .I1 (g10423), .I2 (I15999));
ND2X1 gate9347(.O (I5371), .I1 (g971), .I2 (g976));
ND2X1 gate9348(.O (g2215), .I1 (I5185), .I2 (I5186));
ND2X1 gate9349(.O (g7101), .I1 (g6617), .I2 (g2364));
ND2X1 gate9350(.O (I5675), .I1 (g1218), .I2 (g1223));
ND2X1 gate9351(.O (I8544), .I1 (g4218), .I2 (I8543));
ND2X1 gate9352(.O (g6577), .I1 (I10520), .I2 (I10521));
ND2X1 gate9353(.O (I5297), .I1 (g798), .I2 (I5295));
ND2X1 gate9354(.O (I13537), .I1 (g658), .I2 (g8157));
ND2X1 gate9355(.O (I13283), .I1 (g1927), .I2 (g8159));
ND2X1 gate9356(.O (g4749), .I1 (g3710), .I2 (g2061));
ND2X1 gate9357(.O (I11982), .I1 (g1482), .I2 (I11980));
ND2X1 gate9358(.O (I8514), .I1 (g4873), .I2 (I8513));
ND2X1 gate9359(.O (I13091), .I1 (g1840), .I2 (I13089));
ND2X1 gate9360(.O (g2943), .I1 (I6125), .I2 (I6126));
ND2X1 gate9361(.O (I15908), .I1 (g10302), .I2 (I15906));
ND2X1 gate9362(.O (I6879), .I1 (g3301), .I2 (g1351));
ND2X1 gate9363(.O (I8763), .I1 (g1129), .I2 (I8761));
ND2X1 gate9364(.O (I5449), .I1 (g1235), .I2 (g991));
ND3X1 gate9365(.O (g8825), .I1 (g8502), .I2 (g8738), .I3 (g8506));
ND2X1 gate9366(.O (I16007), .I1 (g10424), .I2 (g2689));
ND2X1 gate9367(.O (I5865), .I1 (g2107), .I2 (g2105));
ND2X1 gate9368(.O (I5604), .I1 (g1149), .I2 (g1153));
ND2X1 gate9369(.O (g2433), .I1 (I5517), .I2 (I5518));
ND2X1 gate9370(.O (I6111), .I1 (g1494), .I2 (I6109));
ND2X1 gate9371(.O (g2096), .I1 (I4929), .I2 (I4930));
ND2X1 gate9372(.O (I13522), .I1 (g695), .I2 (I13521));
ND2X1 gate9373(.O (I10770), .I1 (g5944), .I2 (I10769));
ND2X1 gate9374(.O (g6027), .I1 (g4566), .I2 (g4921));
ND4X1 gate9375(.O (g7992), .I1 (g7011), .I2 (g7574), .I3 (g6984), .I4 (g6974));
ND2X1 gate9376(.O (I5539), .I1 (g1270), .I2 (I5538));
ND2X1 gate9377(.O (I17394), .I1 (g11415), .I2 (I17393));
ND2X1 gate9378(.O (I13553), .I1 (g668), .I2 (I13552));
ND2X1 gate9379(.O (I8642), .I1 (g516), .I2 (I8640));
ND2X1 gate9380(.O (g7573), .I1 (I12046), .I2 (I12047));
ND2X1 gate9381(.O (g11416), .I1 (I17296), .I2 (I17297));
ND2X1 gate9382(.O (g6003), .I1 (g5552), .I2 (g5548));
ND2X1 gate9383(.O (g8934), .I1 (I14278), .I2 (I14279));
ND2X1 gate9384(.O (I15992), .I1 (g10422), .I2 (g2677));
ND2X1 gate9385(.O (I7683), .I1 (g1023), .I2 (g3460));
ND2X1 gate9386(.O (I4910), .I1 (g386), .I2 (g318));
ND4X1 gate9387(.O (g3209), .I1 (g2550), .I2 (g2061), .I3 (g2564), .I4 (g2571));
ND2X1 gate9388(.O (I6794), .I1 (g143), .I2 (I6792));
ND2X1 gate9389(.O (I10521), .I1 (g822), .I2 (I10519));
ND2X1 gate9390(.O (I5486), .I1 (g1011), .I2 (I5484));
ND2X1 gate9391(.O (I15442), .I1 (g10035), .I2 (I15441));
ND2X1 gate9392(.O (g6858), .I1 (I10931), .I2 (I10932));
ND2X1 gate9393(.O (I5185), .I1 (g1415), .I2 (I5184));
ND2X1 gate9394(.O (g5304), .I1 (I8779), .I2 (I8780));
ND2X1 gate9395(.O (g2354), .I1 (g1515), .I2 (g1520));
ND2X1 gate9396(.O (I15615), .I1 (g10043), .I2 (g10153));
ND2X1 gate9397(.O (I17281), .I1 (g11360), .I2 (g11357));
ND2X1 gate9398(.O (I5470), .I1 (g999), .I2 (I5468));
ND2X1 gate9399(.O (I11509), .I1 (g6580), .I2 (I11508));
ND2X1 gate9400(.O (I5025), .I1 (g1275), .I2 (I5023));
ND2X1 gate9401(.O (I11508), .I1 (g6580), .I2 (g1806));
ND2X1 gate9402(.O (I15430), .I1 (g10047), .I2 (g10044));
ND2X1 gate9403(.O (I14612), .I1 (g9204), .I2 (g611));
ND2X1 gate9404(.O (g4675), .I1 (g4073), .I2 (g3247));
ND2X1 gate9405(.O (I14272), .I1 (g1822), .I2 (I14270));
ND2X1 gate9406(.O (g2979), .I1 (I6208), .I2 (I6209));
ND2X1 gate9407(.O (I17290), .I1 (g11363), .I2 (I17288));
ND2X1 gate9408(.O (g5269), .I1 (I8716), .I2 (I8717));
ND2X1 gate9409(.O (g4297), .I1 (I7563), .I2 (I7564));
ND2X1 gate9410(.O (I12002), .I1 (g7082), .I2 (g153));
ND2X1 gate9411(.O (I5006), .I1 (g421), .I2 (I5005));
ND2X1 gate9412(.O (I12128), .I1 (g170), .I2 (I12126));
ND2X1 gate9413(.O (I5105), .I1 (g431), .I2 (I5104));
ND2X1 gate9414(.O (I6323), .I1 (g2050), .I2 (I6322));
ND2X1 gate9415(.O (g7588), .I1 (I12093), .I2 (I12094));
ND2X1 gate9416(.O (I6666), .I1 (g2776), .I2 (I6664));
ND2X1 gate9417(.O (g3623), .I1 (I6761), .I2 (I6762));
ND2X1 gate9418(.O (I5373), .I1 (g976), .I2 (I5371));
ND2X1 gate9419(.O (I8529), .I1 (g481), .I2 (I8527));
ND2X1 gate9420(.O (I5283), .I1 (g758), .I2 (I5282));
ND2X1 gate9421(.O (I7224), .I1 (g2981), .I2 (I7223));
ND2X1 gate9422(.O (I5007), .I1 (g312), .I2 (I5005));
ND2X1 gate9423(.O (I5459), .I1 (g1240), .I2 (g1003));
ND2X1 gate9424(.O (I17297), .I1 (g11369), .I2 (I17295));
ND3X1 gate9425(.O (g8746), .I1 (g8617), .I2 (g6517), .I3 (g6509));
ND2X1 gate9426(.O (I6143), .I1 (g1976), .I2 (g646));
ND2X1 gate9427(.O (I5015), .I1 (g1011), .I2 (I5013));
ND2X1 gate9428(.O (g8932), .I1 (I14264), .I2 (I14265));
ND2X1 gate9429(.O (I16073), .I1 (g845), .I2 (I16072));
ND2X1 gate9430(.O (I6988), .I1 (g2760), .I2 (g986));
ND2X1 gate9431(.O (g3205), .I1 (g1814), .I2 (g2571));
ND2X1 gate9432(.O (I8652), .I1 (g778), .I2 (I8650));
ND2X1 gate9433(.O (I9558), .I1 (g5598), .I2 (I9557));
ND2X1 gate9434(.O (I5203), .I1 (g369), .I2 (I5202));
ND2X1 gate9435(.O (g7533), .I1 (I11936), .I2 (I11937));
ND2X1 gate9436(.O (g3634), .I1 (I6806), .I2 (I6807));
ND2X1 gate9437(.O (I6792), .I1 (g2959), .I2 (g143));
ND2X1 gate9438(.O (g3304), .I1 (I6468), .I2 (I6469));
ND2X1 gate9439(.O (I12145), .I1 (g158), .I2 (I12143));
ND2X1 gate9440(.O (g7596), .I1 (I12127), .I2 (I12128));
ND2X1 gate9441(.O (I13302), .I1 (g8162), .I2 (I13300));
ND2X1 gate9442(.O (I5502), .I1 (g1007), .I2 (I5500));
ND2X1 gate9443(.O (I9574), .I1 (g5608), .I2 (g818));
ND2X1 gate9444(.O (g3273), .I1 (I6448), .I2 (I6449));
ND2X1 gate9445(.O (I8670), .I1 (g4831), .I2 (I8669));
ND2X1 gate9446(.O (I7035), .I1 (g1868), .I2 (I7033));
ND2X1 gate9447(.O (I15453), .I1 (g10051), .I2 (I15451));
ND2X1 gate9448(.O (I8625), .I1 (g4267), .I2 (I8624));
ND2X1 gate9449(.O (I7876), .I1 (g4109), .I2 (I7875));
ND2X1 gate9450(.O (I14203), .I1 (g8825), .I2 (I14202));
ND2X1 gate9451(.O (I15607), .I1 (g10149), .I2 (g10144));
ND2X1 gate9452(.O (g2274), .I1 (I5324), .I2 (I5325));
ND2X1 gate9453(.O (I8740), .I1 (g1121), .I2 (I8738));
ND2X1 gate9454(.O (I17296), .I1 (g11373), .I2 (I17295));
ND2X1 gate9455(.O (g10507), .I1 (g10434), .I2 (g5859));
ND2X1 gate9456(.O (g2325), .I1 (g611), .I2 (g617));
ND2X1 gate9457(.O (I8606), .I1 (g506), .I2 (I8604));
ND2X1 gate9458(.O (I12087), .I1 (g1470), .I2 (I12085));
ND2X1 gate9459(.O (I13249), .I1 (g1891), .I2 (I13248));
ND2X1 gate9460(.O (I13248), .I1 (g1891), .I2 (g8148));
ND2X1 gate9461(.O (I13552), .I1 (g668), .I2 (g8262));
ND2X1 gate9462(.O (g2106), .I1 (I4979), .I2 (I4980));
ND2X1 gate9463(.O (I12069), .I1 (g139), .I2 (I12067));
ND2X1 gate9464(.O (g9204), .I1 (g6019), .I2 (g8942));
ND2X1 gate9465(.O (I12068), .I1 (g7116), .I2 (I12067));
ND2X1 gate9466(.O (I17503), .I1 (g11475), .I2 (g7603));
ND2X1 gate9467(.O (I7877), .I1 (g810), .I2 (I7875));
ND2X1 gate9468(.O (I5165), .I1 (g1508), .I2 (I5164));
ND2X1 gate9469(.O (g6740), .I1 (g6131), .I2 (g2550));
ND2X1 gate9470(.O (I6289), .I1 (g981), .I2 (I6287));
ND2X1 gate9471(.O (I6777), .I1 (g2892), .I2 (g650));
ND2X1 gate9472(.O (g5171), .I1 (I8562), .I2 (I8563));
ND2X1 gate9473(.O (I15891), .I1 (g853), .I2 (I15890));
ND2X1 gate9474(.O (I13090), .I1 (g8006), .I2 (I13089));
ND2X1 gate9475(.O (g11474), .I1 (I17460), .I2 (I17461));
ND4X1 gate9476(.O (g7942), .I1 (g7395), .I2 (g6847), .I3 (g7380), .I4 (g7369));
ND2X1 gate9477(.O (I5538), .I1 (g1270), .I2 (g1023));
ND2X1 gate9478(.O (I7563), .I1 (g3533), .I2 (I7562));
ND2X1 gate9479(.O (I13513), .I1 (g686), .I2 (g8248));
ND2X1 gate9480(.O (g2107), .I1 (I4986), .I2 (I4987));
ND2X1 gate9481(.O (g2223), .I1 (I5203), .I2 (I5204));
ND2X1 gate9482(.O (I13505), .I1 (g677), .I2 (I13504));
ND2X1 gate9483(.O (I6209), .I1 (g802), .I2 (I6207));
ND2X1 gate9484(.O (I12086), .I1 (g6980), .I2 (I12085));
ND2X1 gate9485(.O (I8545), .I1 (g486), .I2 (I8543));
ND2X1 gate9486(.O (I8180), .I1 (g1786), .I2 (I8178));
ND2X1 gate9487(.O (g2115), .I1 (I5014), .I2 (I5015));
ND2X1 gate9488(.O (I8591), .I1 (g501), .I2 (I8589));
ND2X1 gate9489(.O (I10931), .I1 (g6395), .I2 (I10930));
ND2X1 gate9490(.O (I17402), .I1 (g11416), .I2 (I17400));
ND2X1 gate9491(.O (g8307), .I1 (I13294), .I2 (I13295));
ND2X1 gate9492(.O (I12144), .I1 (g7089), .I2 (I12143));
ND2X1 gate9493(.O (I10520), .I1 (g6231), .I2 (I10519));
ND2X1 gate9494(.O (I5263), .I1 (g456), .I2 (g461));
ND2X1 gate9495(.O (g8757), .I1 (g8599), .I2 (g4401));
ND2X1 gate9496(.O (I6714), .I1 (g2961), .I2 (g201));
ND2X1 gate9497(.O (I14211), .I1 (g599), .I2 (I14209));
ND2X1 gate9498(.O (I8515), .I1 (g3513), .I2 (I8513));
ND2X1 gate9499(.O (g2272), .I1 (I5316), .I2 (I5317));
ND2X1 gate9500(.O (I9946), .I1 (g5233), .I2 (g1796));
ND2X1 gate9501(.O (I8750), .I1 (g4613), .I2 (g1125));
ND2X1 gate9502(.O (I5605), .I1 (g1149), .I2 (I5604));
ND2X1 gate9503(.O (g8880), .I1 (I14203), .I2 (I14204));
ND2X1 gate9504(.O (I16051), .I1 (g837), .I2 (g10371));
ND2X1 gate9505(.O (I16072), .I1 (g845), .I2 (g10373));
ND2X1 gate9506(.O (g10440), .I1 (g10360), .I2 (g6037));
ND2X1 gate9507(.O (g8612), .I1 (I13858), .I2 (I13859));
ND2X1 gate9508(.O (I15872), .I1 (g2713), .I2 (I15870));
ND2X1 gate9509(.O (I8528), .I1 (g4879), .I2 (I8527));
ND2X1 gate9510(.O (g8629), .I1 (I13901), .I2 (I13902));
ND4X1 gate9511(.O (g8542), .I1 (g2571), .I2 (g1828), .I3 (g1814), .I4 (g8390));
ND2X1 gate9512(.O (I9947), .I1 (g5233), .I2 (I9946));
ND2X1 gate9513(.O (I6838), .I1 (g806), .I2 (I6836));
ND2X1 gate9514(.O (g7583), .I1 (I12068), .I2 (I12069));
ND2X1 gate9515(.O (g4803), .I1 (g3664), .I2 (g2356));
ND2X1 gate9516(.O (I17307), .I1 (g11377), .I2 (I17305));
ND2X1 gate9517(.O (g4538), .I1 (g3475), .I2 (g2399));
ND2X1 gate9518(.O (I15452), .I1 (g10058), .I2 (I15451));
ND2X1 gate9519(.O (I13857), .I1 (g8538), .I2 (g1448));
ND2X1 gate9520(.O (I14202), .I1 (g8825), .I2 (g591));
ND2X1 gate9521(.O (I13765), .I1 (g731), .I2 (g8417));
ND2X1 gate9522(.O (g2260), .I1 (I5296), .I2 (I5297));
ND4X1 gate9523(.O (g7986), .I1 (g7011), .I2 (g6995), .I3 (g6984), .I4 (g7550));
ND2X1 gate9524(.O (g5226), .I1 (I8670), .I2 (I8671));
ND2X1 gate9525(.O (g8512), .I1 (g3723), .I2 (g8366));
ND2X1 gate9526(.O (I16046), .I1 (g10370), .I2 (I16044));
ND2X1 gate9527(.O (I13504), .I1 (g677), .I2 (g8247));
ND2X1 gate9528(.O (g10447), .I1 (g10363), .I2 (g5360));
ND2X1 gate9529(.O (g2167), .I1 (I5105), .I2 (I5106));
ND2X1 gate9530(.O (I8804), .I1 (g4677), .I2 (I8803));
ND2X1 gate9531(.O (g10472), .I1 (I16016), .I2 (I16017));
ND2X1 gate9532(.O (I17487), .I1 (g11474), .I2 (I17485));
ND2X1 gate9533(.O (I4995), .I1 (g416), .I2 (g309));
ND2X1 gate9534(.O (I12093), .I1 (g6944), .I2 (I12092));
ND4X1 gate9535(.O (g7987), .I1 (g7011), .I2 (g6995), .I3 (g7562), .I4 (g6974));
ND2X1 gate9536(.O (g5227), .I1 (I8677), .I2 (I8678));
ND2X1 gate9537(.O (I5126), .I1 (g1386), .I2 (g1389));
ND2X1 gate9538(.O (g2321), .I1 (I5372), .I2 (I5373));
ND2X1 gate9539(.O (g7547), .I1 (I11974), .I2 (I11975));
ND2X1 gate9540(.O (I17306), .I1 (g11381), .I2 (I17305));
ND3X1 gate9541(.O (g6548), .I1 (g6132), .I2 (g6124), .I3 (g6122));
ND2X1 gate9542(.O (I11995), .I1 (g7107), .I2 (g127));
ND2X1 gate9543(.O (I7225), .I1 (g1781), .I2 (I7223));
ND2X1 gate9544(.O (I11261), .I1 (g6775), .I2 (g826));
ND3X1 gate9545(.O (g8843), .I1 (g8542), .I2 (g8757), .I3 (g8545));
ND2X1 gate9546(.O (g2938), .I1 (I6110), .I2 (I6111));
ND2X1 gate9547(.O (I4942), .I1 (g396), .I2 (I4941));
ND2X1 gate9548(.O (g10394), .I1 (I15899), .I2 (I15900));
ND2X1 gate9549(.O (g8549), .I1 (g5527), .I2 (g8390));
ND2X1 gate9550(.O (g3070), .I1 (g2016), .I2 (g1206));
ND2X1 gate9551(.O (I4954), .I1 (g401), .I2 (g327));
ND2X1 gate9552(.O (I5023), .I1 (g995), .I2 (g1275));
ND2X1 gate9553(.O (g10446), .I1 (g10443), .I2 (g5350));
ND2X1 gate9554(.O (I16081), .I1 (g10374), .I2 (I16079));
ND2X1 gate9555(.O (I8641), .I1 (g4278), .I2 (I8640));
ND2X1 gate9556(.O (I6178), .I1 (g197), .I2 (I6176));
ND2X1 gate9557(.O (I12075), .I1 (g7098), .I2 (I12074));
ND2X1 gate9558(.O (I5127), .I1 (g1386), .I2 (I5126));
ND2X1 gate9559(.O (I5451), .I1 (g991), .I2 (I5449));
ND2X1 gate9560(.O (g4168), .I1 (I7322), .I2 (I7323));
ND2X1 gate9561(.O (I6288), .I1 (g2091), .I2 (I6287));
ND2X1 gate9562(.O (I8179), .I1 (g3685), .I2 (I8178));
ND2X1 gate9563(.O (I4912), .I1 (g318), .I2 (I4910));
ND2X1 gate9564(.O (I6805), .I1 (g3268), .I2 (g471));
ND3X1 gate9565(.O (g3766), .I1 (g2439), .I2 (g3222), .I3 (g2493));
ND2X1 gate9566(.O (g3087), .I1 (I6288), .I2 (I6289));
ND2X1 gate9567(.O (I17486), .I1 (g11384), .I2 (I17485));
ND2X1 gate9568(.O (I4929), .I1 (g391), .I2 (I4928));
ND2X1 gate9569(.O (I15890), .I1 (g853), .I2 (g10286));
ND2X1 gate9570(.O (I16331), .I1 (g10616), .I2 (I16330));
ND2X1 gate9571(.O (I9575), .I1 (g5608), .I2 (I9574));
ND2X1 gate9572(.O (I13887), .I1 (g8532), .I2 (I13886));
ND2X1 gate9573(.O (g5308), .I1 (I8787), .I2 (I8788));
ND2X1 gate9574(.O (I13529), .I1 (g704), .I2 (g8253));
ND2X1 gate9575(.O (I6208), .I1 (g2534), .I2 (I6207));
ND2X1 gate9576(.O (g5217), .I1 (I8641), .I2 (I8642));
ND2X1 gate9577(.O (I5316), .I1 (g1032), .I2 (I5315));
ND2X1 gate9578(.O (g2111), .I1 (I5006), .I2 (I5007));
ND2X1 gate9579(.O (g10366), .I1 (g10285), .I2 (g5392));
ND2X1 gate9580(.O (I5034), .I1 (g1015), .I2 (g1019));
ND2X1 gate9581(.O (I13869), .I1 (g1403), .I2 (I13867));
ND2X1 gate9582(.O (I13868), .I1 (g8523), .I2 (I13867));
ND2X1 gate9583(.O (I15999), .I1 (g10423), .I2 (g2683));
ND2X1 gate9584(.O (I13259), .I1 (g1900), .I2 (I13258));
ND4X1 gate9585(.O (g3261), .I1 (g2229), .I2 (g2222), .I3 (g2211), .I4 (g2202));
ND2X1 gate9586(.O (g10481), .I1 (I16073), .I2 (I16074));
ND2X1 gate9587(.O (g2180), .I1 (I5136), .I2 (I5137));
ND3X1 gate9588(.O (g4976), .I1 (g2310), .I2 (g4604), .I3 (g3807));
ND2X1 gate9589(.O (g8506), .I1 (g3475), .I2 (g8366));
ND2X1 gate9590(.O (g2380), .I1 (I5460), .I2 (I5461));
ND2X1 gate9591(.O (I13258), .I1 (g1900), .I2 (g8153));
ND2X1 gate9592(.O (I5013), .I1 (g1007), .I2 (g1011));
ND2X1 gate9593(.O (g5196), .I1 (I8605), .I2 (I8606));
ND2X1 gate9594(.O (I10930), .I1 (g6395), .I2 (g5555));
ND2X1 gate9595(.O (I6770), .I1 (g3257), .I2 (g382));
ND2X1 gate9596(.O (g11449), .I1 (I17401), .I2 (I17402));
ND2X1 gate9597(.O (g11448), .I1 (I17394), .I2 (I17395));
ND2X1 gate9598(.O (I15717), .I1 (g10231), .I2 (I15716));
ND2X1 gate9599(.O (I5317), .I1 (g1027), .I2 (I5315));
ND2X1 gate9600(.O (I14210), .I1 (g8824), .I2 (I14209));
ND2X1 gate9601(.O (I17569), .I1 (g1610), .I2 (I17567));
ND2X1 gate9602(.O (I13878), .I1 (g1444), .I2 (I13876));
ND2X1 gate9603(.O (g8545), .I1 (g3710), .I2 (g8390));
ND2X1 gate9604(.O (g2515), .I1 (I5605), .I2 (I5606));
ND2X1 gate9605(.O (I14443), .I1 (g8970), .I2 (I14442));
ND2X1 gate9606(.O (g7557), .I1 (I11996), .I2 (I11997));
ND2X1 gate9607(.O (g8180), .I1 (I13090), .I2 (I13091));
ND2X1 gate9608(.O (I14279), .I1 (g1828), .I2 (I14277));
ND2X1 gate9609(.O (I17568), .I1 (g11496), .I2 (I17567));
ND2X1 gate9610(.O (I13886), .I1 (g8532), .I2 (g1440));
ND2X1 gate9611(.O (I7322), .I1 (g3047), .I2 (I7321));
ND2X1 gate9612(.O (I6990), .I1 (g986), .I2 (I6988));
ND2X1 gate9613(.O (I14278), .I1 (g8847), .I2 (I14277));
ND2X1 gate9614(.O (I7033), .I1 (g3089), .I2 (g1868));
ND2X1 gate9615(.O (I9006), .I1 (g4492), .I2 (g1791));
ND2X1 gate9616(.O (g8507), .I1 (g3738), .I2 (g8366));
ND2X1 gate9617(.O (I5460), .I1 (g1240), .I2 (I5459));
ND2X1 gate9618(.O (g4588), .I1 (g3440), .I2 (g2745));
ND2X1 gate9619(.O (I4986), .I1 (g999), .I2 (I4985));
ND3X1 gate9620(.O (g3247), .I1 (g1828), .I2 (g2564), .I3 (g2571));
ND2X1 gate9621(.O (I8651), .I1 (g4824), .I2 (I8650));
ND2X1 gate9622(.O (I13545), .I1 (g713), .I2 (I13544));
ND2X1 gate9623(.O (g8628), .I1 (I13894), .I2 (I13895));
ND2X1 gate9624(.O (I6138), .I1 (g378), .I2 (I6136));
ND2X1 gate9625(.O (I12074), .I1 (g7098), .I2 (g174));
ND2X1 gate9626(.O (g8630), .I1 (I13908), .I2 (I13909));
ND2X1 gate9627(.O (I13078), .I1 (g7963), .I2 (I13076));
ND2X1 gate9628(.O (I6109), .I1 (g2205), .I2 (g1494));
ND2X1 gate9629(.O (g8300), .I1 (I13259), .I2 (I13260));
ND2X1 gate9630(.O (I5501), .I1 (g1255), .I2 (I5500));
ND2X1 gate9631(.O (I17586), .I1 (g11515), .I2 (I17584));
ND2X1 gate9632(.O (I12092), .I1 (g6944), .I2 (g1490));
ND2X1 gate9633(.O (I13901), .I1 (g8520), .I2 (I13900));
ND2X1 gate9634(.O (I8795), .I1 (g4672), .I2 (g1145));
ND2X1 gate9635(.O (I6201), .I1 (g766), .I2 (I6199));
ND2X1 gate9636(.O (I14217), .I1 (g8826), .I2 (I14216));
ND2X1 gate9637(.O (I9007), .I1 (g4492), .I2 (I9006));
ND2X1 gate9638(.O (I13561), .I1 (g8263), .I2 (I13559));
ND2X1 gate9639(.O (I15716), .I1 (g10231), .I2 (g10229));
ND2X1 gate9640(.O (I6449), .I1 (g1776), .I2 (I6447));
ND2X1 gate9641(.O (I13295), .I1 (g8161), .I2 (I13293));
ND2X1 gate9642(.O (I4987), .I1 (g1003), .I2 (I4985));
ND2X1 gate9643(.O (I6715), .I1 (g2961), .I2 (I6714));
ND2X1 gate9644(.O (I17493), .I1 (g11475), .I2 (I17492));
ND2X1 gate9645(.O (I12215), .I1 (g7061), .I2 (I12214));
ND2X1 gate9646(.O (g2372), .I1 (I5450), .I2 (I5451));
ND2X1 gate9647(.O (g7062), .I1 (I11262), .I2 (I11263));
ND2X1 gate9648(.O (g2988), .I1 (I6225), .I2 (I6226));
ND2X1 gate9649(.O (I13309), .I1 (g617), .I2 (I13307));
ND2X1 gate9650(.O (g8839), .I1 (g8750), .I2 (g4401));
ND2X1 gate9651(.O (g2555), .I1 (I5676), .I2 (I5677));
ND2X1 gate9652(.O (g3662), .I1 (I6826), .I2 (I6827));
ND2X1 gate9653(.O (I13308), .I1 (g8190), .I2 (I13307));
ND2X1 gate9654(.O (g2792), .I1 (I5879), .I2 (I5880));
ND2X1 gate9655(.O (g4117), .I1 (g3041), .I2 (g3061));
ND2X1 gate9656(.O (I8543), .I1 (g4218), .I2 (g486));
ND2X1 gate9657(.O (g11549), .I1 (I17585), .I2 (I17586));
ND2X1 gate9658(.O (I6881), .I1 (g1351), .I2 (I6879));
ND2X1 gate9659(.O (I12138), .I1 (g131), .I2 (I12136));
ND2X1 gate9660(.O (I8729), .I1 (g4605), .I2 (I8728));
ND2X1 gate9661(.O (I14216), .I1 (g8826), .I2 (g605));
ND2X1 gate9662(.O (g10384), .I1 (I15871), .I2 (I15872));
ND2X1 gate9663(.O (I13260), .I1 (g8153), .I2 (I13258));
ND2X1 gate9664(.O (g2776), .I1 (I5866), .I2 (I5867));
ND2X1 gate9665(.O (I8513), .I1 (g4873), .I2 (g3513));
ND2X1 gate9666(.O (I13559), .I1 (g722), .I2 (g8263));
ND2X1 gate9667(.O (I8178), .I1 (g3685), .I2 (g1786));
ND2X1 gate9668(.O (g3631), .I1 (I6793), .I2 (I6794));
ND2X1 gate9669(.O (I6487), .I1 (g2306), .I2 (g1227));
ND2X1 gate9670(.O (I16080), .I1 (g849), .I2 (I16079));
ND2X1 gate9671(.O (I13893), .I1 (g8529), .I2 (g1436));
ND2X1 gate9672(.O (I12115), .I1 (g162), .I2 (I12113));
ND2X1 gate9673(.O (I6748), .I1 (g1453), .I2 (I6746));
ND2X1 gate9674(.O (I13544), .I1 (g713), .I2 (g8259));
ND2X1 gate9675(.O (I5484), .I1 (g1250), .I2 (g1011));
ND2X1 gate9676(.O (I4928), .I1 (g391), .I2 (g321));
ND2X1 gate9677(.O (I6226), .I1 (g1346), .I2 (I6224));
ND2X1 gate9678(.O (I8805), .I1 (g1113), .I2 (I8803));
ND2X1 gate9679(.O (I4930), .I1 (g321), .I2 (I4928));
ND2X1 gate9680(.O (I15880), .I1 (g2719), .I2 (I15878));
ND2X1 gate9681(.O (I14265), .I1 (g1814), .I2 (I14263));
ND2X1 gate9682(.O (I16031), .I1 (g829), .I2 (I16030));
ND2X1 gate9683(.O (g3585), .I1 (I6747), .I2 (I6748));
ND4X1 gate9684(.O (g3041), .I1 (g2364), .I2 (g2399), .I3 (g2374), .I4 (g2382));
ND2X1 gate9685(.O (g8933), .I1 (I14271), .I2 (I14272));
ND2X1 gate9686(.O (I16330), .I1 (g10616), .I2 (g4997));
ND2X1 gate9687(.O (I13267), .I1 (g8154), .I2 (I13265));
ND2X1 gate9688(.O (I13294), .I1 (g1882), .I2 (I13293));
ND2X1 gate9689(.O (g10231), .I1 (I15616), .I2 (I15617));
ND2X1 gate9690(.O (I14442), .I1 (g8970), .I2 (g1834));
ND2X1 gate9691(.O (I6793), .I1 (g2959), .I2 (I6792));
ND2X1 gate9692(.O (I4966), .I1 (g330), .I2 (I4964));
ND2X1 gate9693(.O (I8752), .I1 (g1125), .I2 (I8750));
ND2X1 gate9694(.O (I15432), .I1 (g10044), .I2 (I15430));
ND2X1 gate9695(.O (I12214), .I1 (g7061), .I2 (g2518));
ND2X1 gate9696(.O (g10511), .I1 (g10438), .I2 (g6032));
ND2X1 gate9697(.O (g3011), .I1 (g591), .I2 (g2382));
ND2X1 gate9698(.O (g5103), .I1 (I8480), .I2 (I8481));
ND2X1 gate9699(.O (I16087), .I1 (g861), .I2 (I16086));
ND2X1 gate9700(.O (g3734), .I1 (g3039), .I2 (g599));
ND2X1 gate9701(.O (I6664), .I1 (g2792), .I2 (g2776));
ND2X1 gate9702(.O (g8882), .I1 (I14217), .I2 (I14218));
ND2X1 gate9703(.O (I4955), .I1 (g401), .I2 (I4954));
ND2X1 gate9704(.O (I8786), .I1 (g4639), .I2 (g1141));
ND3X1 gate9705(.O (g3992), .I1 (g2571), .I2 (g2550), .I3 (g2990));
ND2X1 gate9706(.O (g10480), .I1 (I16066), .I2 (I16067));
ND2X1 gate9707(.O (I11915), .I1 (g6935), .I2 (I11914));
ND2X1 gate9708(.O (I8770), .I1 (g4619), .I2 (g1133));
ND2X1 gate9709(.O (I5516), .I1 (g1260), .I2 (g1019));
ND2X1 gate9710(.O (g8541), .I1 (g4001), .I2 (g8390));
ND2X1 gate9711(.O (I6188), .I1 (g466), .I2 (I6186));
ND2X1 gate9712(.O (g5147), .I1 (I8544), .I2 (I8545));
ND3X1 gate9713(.O (g8744), .I1 (g8617), .I2 (g6509), .I3 (g6971));
ND2X1 gate9714(.O (I5892), .I1 (g750), .I2 (I5891));
ND2X1 gate9715(.O (g8558), .I1 (I13766), .I2 (I13767));
ND2X1 gate9716(.O (I15258), .I1 (g9980), .I2 (I15256));
ND2X1 gate9717(.O (I13266), .I1 (g1909), .I2 (I13265));
ND2X1 gate9718(.O (I8787), .I1 (g4639), .I2 (I8786));
ND2X1 gate9719(.O (I6826), .I1 (g3281), .I2 (I6825));
ND2X1 gate9720(.O (I17283), .I1 (g11357), .I2 (I17281));
ND3X1 gate9721(.O (g5013), .I1 (g4749), .I2 (g3247), .I3 (g3205));
ND2X1 gate9722(.O (I17492), .I1 (g11475), .I2 (g3623));
ND2X1 gate9723(.O (g8511), .I1 (g5277), .I2 (g8366));
ND2X1 gate9724(.O (I16079), .I1 (g849), .I2 (g10374));
ND2X1 gate9725(.O (I5035), .I1 (g1015), .I2 (I5034));
ND2X1 gate9726(.O (I5517), .I1 (g1260), .I2 (I5516));
ND2X1 gate9727(.O (I7223), .I1 (g2981), .I2 (g1781));
ND2X1 gate9728(.O (I16086), .I1 (g861), .I2 (g10375));
ND2X1 gate9729(.O (g5317), .I1 (I8796), .I2 (I8797));
ND2X1 gate9730(.O (I15879), .I1 (g10359), .I2 (I15878));
ND2X1 gate9731(.O (I15878), .I1 (g10359), .I2 (g2719));
ND2X1 gate9732(.O (I12114), .I1 (g7093), .I2 (I12113));
ND2X1 gate9733(.O (I12107), .I1 (g7113), .I2 (I12106));
ND2X1 gate9734(.O (g2500), .I1 (g178), .I2 (g182));
ND2X1 gate9735(.O (I15994), .I1 (g2677), .I2 (I15992));
ND4X1 gate9736(.O (g7934), .I1 (g7395), .I2 (g6847), .I3 (g7279), .I4 (g7369));
ND2X1 gate9737(.O (g10469), .I1 (g10430), .I2 (g5999));
ND2X1 gate9738(.O (I14264), .I1 (g8843), .I2 (I14263));
ND2X1 gate9739(.O (I6448), .I1 (g2264), .I2 (I6447));
ND2X1 gate9740(.O (I13285), .I1 (g8159), .I2 (I13283));
ND2X1 gate9741(.O (g10468), .I1 (I16000), .I2 (I16001));
ND2X1 gate9742(.O (I6827), .I1 (g770), .I2 (I6825));
ND2X1 gate9743(.O (g8623), .I1 (I13877), .I2 (I13878));
ND2X1 gate9744(.O (I13900), .I1 (g8520), .I2 (g1428));
ND2X1 gate9745(.O (g2795), .I1 (I5892), .I2 (I5893));
ND2X1 gate9746(.O (I8575), .I1 (g4234), .I2 (g496));
ND2X1 gate9747(.O (I14209), .I1 (g8824), .I2 (g599));
ND2X1 gate9748(.O (I13560), .I1 (g722), .I2 (I13559));
ND2X1 gate9749(.O (I8715), .I1 (g4601), .I2 (g4052));
ND2X1 gate9750(.O (I8604), .I1 (g4259), .I2 (g506));
ND2X1 gate9751(.O (I16017), .I1 (g2695), .I2 (I16015));
ND2X1 gate9752(.O (I4941), .I1 (g396), .I2 (g324));
ND2X1 gate9753(.O (g2205), .I1 (I5165), .I2 (I5166));
ND3X1 gate9754(.O (g3753), .I1 (g2382), .I2 (g2364), .I3 (g2800));
ND2X1 gate9755(.O (I6467), .I1 (g23), .I2 (g2479));
ND2X1 gate9756(.O (I14614), .I1 (g611), .I2 (I14612));
ND2X1 gate9757(.O (g2104), .I1 (I4965), .I2 (I4966));
ND2X1 gate9758(.O (g2099), .I1 (I4942), .I2 (I4943));
ND2X1 gate9759(.O (I16023), .I1 (g10426), .I2 (g2701));
ND2X1 gate9760(.O (g10479), .I1 (I16059), .I2 (I16060));
ND3X1 gate9761(.O (g8737), .I1 (g2317), .I2 (g4921), .I3 (g8688));
ND2X1 gate9762(.O (g5942), .I1 (I9575), .I2 (I9576));
ND2X1 gate9763(.O (g10478), .I1 (I16052), .I2 (I16053));
ND2X1 gate9764(.O (I12004), .I1 (g153), .I2 (I12002));
ND2X1 gate9765(.O (I4911), .I1 (g386), .I2 (I4910));
ND2X1 gate9766(.O (I11914), .I1 (g6935), .I2 (g1494));
ND2X1 gate9767(.O (g7960), .I1 (g7409), .I2 (g5573));
ND2X1 gate9768(.O (I5295), .I1 (g794), .I2 (g798));
ND2X1 gate9769(.O (I12106), .I1 (g7113), .I2 (g135));
ND2X1 gate9770(.O (I8728), .I1 (g4605), .I2 (g1117));
ND2X1 gate9771(.O (g3681), .I1 (I6837), .I2 (I6838));
ND2X1 gate9772(.O (I11907), .I1 (g6967), .I2 (g1474));
ND2X1 gate9773(.O (I13907), .I1 (g8526), .I2 (g1432));
ND2X1 gate9774(.O (I8730), .I1 (g1117), .I2 (I8728));
ND2X1 gate9775(.O (g8551), .I1 (g3967), .I2 (g8390));
ND2X1 gate9776(.O (I4980), .I1 (g333), .I2 (I4978));
ND2X1 gate9777(.O (g2961), .I1 (I6177), .I2 (I6178));
ND2X1 gate9778(.O (g6019), .I1 (g617), .I2 (g4921));
ND2X1 gate9779(.O (I16016), .I1 (g10425), .I2 (I16015));
ND2X1 gate9780(.O (I11935), .I1 (g7004), .I2 (g1458));
ND2X1 gate9781(.O (I8678), .I1 (g1027), .I2 (I8676));
ND2X1 gate9782(.O (I17051), .I1 (g10923), .I2 (g11249));
ND2X1 gate9783(.O (g4482), .I1 (I7864), .I2 (I7865));
ND2X1 gate9784(.O (g7592), .I1 (I12107), .I2 (I12108));
ND2X1 gate9785(.O (g3460), .I1 (I6665), .I2 (I6666));
ND4X1 gate9786(.O (g7932), .I1 (g7395), .I2 (g6847), .I3 (g7279), .I4 (g7273));
ND2X1 gate9787(.O (g7624), .I1 (I12215), .I2 (I12216));
ND4X1 gate9788(.O (g7953), .I1 (g7395), .I2 (g7390), .I3 (g7380), .I4 (g7369));
ND2X1 gate9789(.O (g8414), .I1 (I13553), .I2 (I13554));
ND2X1 gate9790(.O (I6168), .I1 (g153), .I2 (I6166));
ND2X1 gate9791(.O (I5229), .I1 (g182), .I2 (g148));
ND2X1 gate9792(.O (I6772), .I1 (g382), .I2 (I6770));
ND2X1 gate9793(.O (I16030), .I1 (g829), .I2 (g10368));
ND2X1 gate9794(.O (I13284), .I1 (g1927), .I2 (I13283));
ND2X1 gate9795(.O (I16065), .I1 (g10428), .I2 (g2765));
ND2X1 gate9796(.O (g2947), .I1 (I6137), .I2 (I6138));
ND2X1 gate9797(.O (I7321), .I1 (g3047), .I2 (g1231));
ND2X1 gate9798(.O (g2437), .I1 (I5529), .I2 (I5530));
ND2X1 gate9799(.O (g2102), .I1 (I4955), .I2 (I4956));
ND2X1 gate9800(.O (I17282), .I1 (g11360), .I2 (I17281));
ND2X1 gate9801(.O (I5620), .I1 (g1771), .I2 (I5618));
ND2X1 gate9802(.O (I8664), .I1 (g476), .I2 (I8662));
ND2X1 gate9803(.O (g7524), .I1 (I11915), .I2 (I11916));
ND2X1 gate9804(.O (g7717), .I1 (g6863), .I2 (g3206));
ND2X1 gate9805(.O (I16467), .I1 (g10716), .I2 (g10518));
ND2X1 gate9806(.O (I4972), .I1 (g991), .I2 (I4971));
ND2X1 gate9807(.O (I13554), .I1 (g8262), .I2 (I13552));
ND2X1 gate9808(.O (I16037), .I1 (g10427), .I2 (g2707));
ND2X1 gate9809(.O (g8302), .I1 (I13273), .I2 (I13274));
ND2X1 gate9810(.O (I4943), .I1 (g324), .I2 (I4941));
ND2X1 gate9811(.O (I5485), .I1 (g1250), .I2 (I5484));
ND2X1 gate9812(.O (g5527), .I1 (g3978), .I2 (g4749));
ND2X1 gate9813(.O (I10509), .I1 (g786), .I2 (I10507));
ND2X1 gate9814(.O (g7599), .I1 (I12144), .I2 (I12145));
ND2X1 gate9815(.O (I10508), .I1 (g6221), .I2 (I10507));
ND2X1 gate9816(.O (I6126), .I1 (g1419), .I2 (I6124));
ND2X1 gate9817(.O (I8671), .I1 (g814), .I2 (I8669));
ND2X1 gate9818(.O (I6760), .I1 (g2943), .I2 (g1448));
ND2X1 gate9819(.O (g3626), .I1 (I6778), .I2 (I6779));
ND2X1 gate9820(.O (I11973), .I1 (g7001), .I2 (g1462));
ND2X1 gate9821(.O (g2389), .I1 (I5469), .I2 (I5470));
ND2X1 gate9822(.O (I15617), .I1 (g10153), .I2 (I15615));
ND2X1 gate9823(.O (g5277), .I1 (g3734), .I2 (g4538));
ND2X1 gate9824(.O (I5005), .I1 (g421), .I2 (g312));
ND2X1 gate9825(.O (I6779), .I1 (g650), .I2 (I6777));
ND2X1 gate9826(.O (I6665), .I1 (g2792), .I2 (I6664));
ND2X1 gate9827(.O (I8589), .I1 (g4251), .I2 (g501));
ND2X1 gate9828(.O (g8412), .I1 (I13545), .I2 (I13546));
ND2X1 gate9829(.O (g2963), .I1 (I6187), .I2 (I6188));
ND2X1 gate9830(.O (I12045), .I1 (g6951), .I2 (g1486));
ND2X1 gate9831(.O (I16053), .I1 (g10371), .I2 (I16051));
ND2X1 gate9832(.O (g2109), .I1 (I4996), .I2 (I4997));
ND2X1 gate9833(.O (g11418), .I1 (I17306), .I2 (I17307));
ND2X1 gate9834(.O (I13539), .I1 (g8157), .I2 (I13537));
ND2X1 gate9835(.O (g10475), .I1 (I16031), .I2 (I16032));
ND2X1 gate9836(.O (I5324), .I1 (g1336), .I2 (I5323));
ND2X1 gate9837(.O (I13538), .I1 (g658), .I2 (I13537));
ND2X1 gate9838(.O (I5469), .I1 (g1245), .I2 (I5468));
ND2X1 gate9839(.O (I5540), .I1 (g1023), .I2 (I5538));
ND2X1 gate9840(.O (I17505), .I1 (g7603), .I2 (I17503));
ND2X1 gate9841(.O (I11241), .I1 (g6760), .I2 (g790));
ND2X1 gate9842(.O (I8803), .I1 (g4677), .I2 (g1113));
ND2X1 gate9843(.O (I12061), .I1 (g6961), .I2 (I12060));
ND2X1 gate9844(.O (I8780), .I1 (g1137), .I2 (I8778));
ND3X1 gate9845(.O (g8745), .I1 (g8617), .I2 (g6517), .I3 (g6964));
ND2X1 gate9846(.O (I4979), .I1 (g411), .I2 (I4978));
ND2X1 gate9847(.O (g8109), .I1 (g5052), .I2 (g7853));
ND2X1 gate9848(.O (g8309), .I1 (I13308), .I2 (I13309));
ND2X1 gate9849(.O (g6758), .I1 (I10770), .I2 (I10771));
ND2X1 gate9850(.O (I16009), .I1 (g2689), .I2 (I16007));
ND2X1 gate9851(.O (I15616), .I1 (g10043), .I2 (I15615));
ND2X1 gate9852(.O (I8662), .I1 (g4286), .I2 (g476));
ND2X1 gate9853(.O (I16008), .I1 (g10424), .I2 (I16007));
ND2X1 gate9854(.O (I13515), .I1 (g8248), .I2 (I13513));
ND2X1 gate9855(.O (I13991), .I1 (g622), .I2 (I13990));
ND2X1 gate9856(.O (g11276), .I1 (I17052), .I2 (I17053));
ND2X1 gate9857(.O (I15900), .I1 (g10287), .I2 (I15898));
ND2X1 gate9858(.O (g2419), .I1 (I5501), .I2 (I5502));
ND2X1 gate9859(.O (I16074), .I1 (g10373), .I2 (I16072));
ND2X1 gate9860(.O (I10769), .I1 (g5944), .I2 (g1801));
ND2X1 gate9861(.O (I7323), .I1 (g1231), .I2 (I7321));
ND2X1 gate9862(.O (g7978), .I1 (g7697), .I2 (g3038));
ND2X1 gate9863(.O (I7875), .I1 (g4109), .I2 (g810));
ND2X1 gate9864(.O (I8562), .I1 (g4227), .I2 (I8561));
ND2X1 gate9865(.O (I15892), .I1 (g10286), .I2 (I15890));
ND2X1 gate9866(.O (g3771), .I1 (I6989), .I2 (I6990));
ND2X1 gate9867(.O (I8605), .I1 (g4259), .I2 (I8604));
ND2X1 gate9868(.O (g10153), .I1 (I15452), .I2 (I15453));
ND2X1 gate9869(.O (g5295), .I1 (I8762), .I2 (I8763));
ND2X1 gate9870(.O (I8751), .I1 (g4613), .I2 (I8750));
ND2X1 gate9871(.O (I15907), .I1 (g6899), .I2 (I15906));
ND2X1 gate9872(.O (I5136), .I1 (g521), .I2 (I5135));
ND2X1 gate9873(.O (I11263), .I1 (g826), .I2 (I11261));
ND2X1 gate9874(.O (I14204), .I1 (g591), .I2 (I14202));
ND2X1 gate9875(.O (g8881), .I1 (I14210), .I2 (I14211));
ND2X1 gate9876(.O (g2105), .I1 (I4972), .I2 (I4973));
ND3X1 gate9877(.O (g5557), .I1 (g4538), .I2 (g3071), .I3 (g3011));
ND2X1 gate9878(.O (I5230), .I1 (g182), .I2 (I5229));
ND2X1 gate9879(.O (I8669), .I1 (g4831), .I2 (g814));
ND2X1 gate9880(.O (g10474), .I1 (I16024), .I2 (I16025));
ND2X1 gate9881(.O (I8772), .I1 (g1133), .I2 (I8770));
ND2X1 gate9882(.O (g2445), .I1 (I5539), .I2 (I5540));
ND2X1 gate9883(.O (g8006), .I1 (g5552), .I2 (g7717));
ND2X1 gate9884(.O (I10932), .I1 (g5555), .I2 (I10930));
ND2X1 gate9885(.O (I17504), .I1 (g11475), .I2 (I17503));
ND2X1 gate9886(.O (I5137), .I1 (g525), .I2 (I5135));
ND2X1 gate9887(.O (g8305), .I1 (I13284), .I2 (I13285));
ND2X1 gate9888(.O (I5891), .I1 (g750), .I2 (g2057));
ND2X1 gate9889(.O (I13273), .I1 (g1918), .I2 (I13272));
ND2X1 gate9890(.O (I8480), .I1 (g4455), .I2 (I8479));
ND2X1 gate9891(.O (g4144), .I1 (g2160), .I2 (g3044));
ND2X1 gate9892(.O (I15906), .I1 (g6899), .I2 (g10302));
ND2X1 gate9893(.O (I5342), .I1 (g315), .I2 (I5341));
ND2X1 gate9894(.O (I13514), .I1 (g686), .I2 (I13513));
ND2X1 gate9895(.O (g8407), .I1 (I13522), .I2 (I13523));
ND2X1 gate9896(.O (g4088), .I1 (I7224), .I2 (I7225));
ND2X1 gate9897(.O (g4488), .I1 (I7876), .I2 (I7877));
ND2X1 gate9898(.O (g7598), .I1 (I12137), .I2 (I12138));
ND3X1 gate9899(.O (g3222), .I1 (g2557), .I2 (g1814), .I3 (g1834));
ND2X1 gate9900(.O (I16052), .I1 (g837), .I2 (I16051));
ND2X1 gate9901(.O (I12127), .I1 (g7103), .I2 (I12126));
ND2X1 gate9902(.O (g10483), .I1 (I16087), .I2 (I16088));
ND2X1 gate9903(.O (g8415), .I1 (I13560), .I2 (I13561));
ND2X1 gate9904(.O (g11415), .I1 (I17289), .I2 (I17290));
ND2X1 gate9905(.O (g6573), .I1 (I10508), .I2 (I10509));
ND2X1 gate9906(.O (I5676), .I1 (g1218), .I2 (I5675));
ND2X1 gate9907(.O (I6778), .I1 (g2892), .I2 (I6777));
ND2X1 gate9908(.O (g9413), .I1 (I14613), .I2 (I14614));
ND2X1 gate9909(.O (I8779), .I1 (g4630), .I2 (I8778));
ND2X1 gate9910(.O (I5592), .I1 (g1696), .I2 (I5591));
ND4X1 gate9911(.O (g8502), .I1 (g2382), .I2 (g605), .I3 (g591), .I4 (g8366));
ND2X1 gate9912(.O (I15609), .I1 (g10144), .I2 (I15607));
ND2X1 gate9913(.O (I15608), .I1 (g10149), .I2 (I15607));
ND3X1 gate9914(.O (g3071), .I1 (g605), .I2 (g2374), .I3 (g2382));
ND2X1 gate9915(.O (g10509), .I1 (g10436), .I2 (g6023));
ND2X1 gate9916(.O (I17461), .I1 (g11448), .I2 (I17459));
ND2X1 gate9917(.O (I13506), .I1 (g8247), .I2 (I13504));
ND2X1 gate9918(.O (I5468), .I1 (g1245), .I2 (g999));
ND2X1 gate9919(.O (g5219), .I1 (I8651), .I2 (I8652));
ND2X1 gate9920(.O (I5677), .I1 (g1223), .I2 (I5675));
ND3X1 gate9921(.O (g8826), .I1 (g8739), .I2 (g8737), .I3 (g8648));
ND2X1 gate9922(.O (I17393), .I1 (g11415), .I2 (g11414));
ND2X1 gate9923(.O (I5866), .I1 (g2107), .I2 (I5865));
ND2X1 gate9924(.O (I12126), .I1 (g7103), .I2 (g170));
ND2X1 gate9925(.O (I4978), .I1 (g411), .I2 (g333));
ND2X1 gate9926(.O (g7587), .I1 (I12086), .I2 (I12087));
ND2X1 gate9927(.O (g5286), .I1 (I8751), .I2 (I8752));
ND2X1 gate9928(.O (g8308), .I1 (I13301), .I2 (I13302));
ND2X1 gate9929(.O (I7864), .I1 (g4099), .I2 (I7863));
ND2X1 gate9930(.O (I11981), .I1 (g6957), .I2 (I11980));
ND2X1 gate9931(.O (I12060), .I1 (g6961), .I2 (g1478));
ND2X1 gate9932(.O (g5225), .I1 (I8663), .I2 (I8664));
ND2X1 gate9933(.O (g11538), .I1 (I17568), .I2 (I17569));
ND2X1 gate9934(.O (I13767), .I1 (g8417), .I2 (I13765));
ND2X1 gate9935(.O (g10396), .I1 (I15907), .I2 (I15908));
ND2X1 gate9936(.O (I11262), .I1 (g6775), .I2 (I11261));
ND2X1 gate9937(.O (I13990), .I1 (g622), .I2 (g8688));
ND2X1 gate9938(.O (I6224), .I1 (g2544), .I2 (g1346));
ND2X1 gate9939(.O (I5867), .I1 (g2105), .I2 (I5865));
ND2X1 gate9940(.O (g2493), .I1 (g1834), .I2 (g1840));
ND2X1 gate9941(.O (I5893), .I1 (g2057), .I2 (I5891));
ND3X1 gate9942(.O (g3062), .I1 (g2369), .I2 (g591), .I3 (g611));
ND2X1 gate9943(.O (I13521), .I1 (g695), .I2 (g8249));
ND2X1 gate9944(.O (I5186), .I1 (g1515), .I2 (I5184));
ND2X1 gate9945(.O (I6771), .I1 (g3257), .I2 (I6770));
ND2X1 gate9946(.O (I5325), .I1 (g1341), .I2 (I5323));
ND2X1 gate9947(.O (I17459), .I1 (g11449), .I2 (g11448));
ND2X1 gate9948(.O (I9557), .I1 (g5598), .I2 (g782));
ND2X1 gate9949(.O (g11414), .I1 (I17282), .I2 (I17283));
ND2X1 gate9950(.O (I12067), .I1 (g7116), .I2 (g139));
ND2X1 gate9951(.O (I12094), .I1 (g1490), .I2 (I12092));
ND2X1 gate9952(.O (I4964), .I1 (g406), .I2 (g330));
ND2X1 gate9953(.O (I13272), .I1 (g1918), .I2 (g8158));
ND2X1 gate9954(.O (I9948), .I1 (g1796), .I2 (I9946));
ND2X1 gate9955(.O (g10302), .I1 (I15717), .I2 (I15718));
ND2X1 gate9956(.O (I16332), .I1 (g4997), .I2 (I16330));
ND2X1 gate9957(.O (I5106), .I1 (g435), .I2 (I5104));
ND2X1 gate9958(.O (g8847), .I1 (g8760), .I2 (g8683));
ND2X1 gate9959(.O (g2257), .I1 (I5283), .I2 (I5284));
ND2X1 gate9960(.O (I12019), .I1 (g7119), .I2 (g166));
ND2X1 gate9961(.O (I15441), .I1 (g10035), .I2 (g10122));
ND2X1 gate9962(.O (I11997), .I1 (g127), .I2 (I11995));
ND2X1 gate9963(.O (I8739), .I1 (g4607), .I2 (I8738));
ND2X1 gate9964(.O (I5461), .I1 (g1003), .I2 (I5459));
ND2X1 gate9965(.O (I13766), .I1 (g731), .I2 (I13765));
ND2X1 gate9966(.O (I8479), .I1 (g4455), .I2 (g3530));
ND2X1 gate9967(.O (I17295), .I1 (g11373), .I2 (g11369));
ND2X1 gate9968(.O (I14271), .I1 (g8840), .I2 (I14270));
ND2X1 gate9969(.O (I4971), .I1 (g991), .I2 (g995));
ND2X1 gate9970(.O (g8301), .I1 (I13266), .I2 (I13267));
ND2X1 gate9971(.O (I6110), .I1 (g2205), .I2 (I6109));
ND2X1 gate9972(.O (g10482), .I1 (I16080), .I2 (I16081));
ND2X1 gate9973(.O (g10779), .I1 (I16468), .I2 (I16469));
ND2X1 gate9974(.O (I6762), .I1 (g1448), .I2 (I6760));
ND2X1 gate9975(.O (I17289), .I1 (g11366), .I2 (I17288));
ND2X1 gate9976(.O (I5315), .I1 (g1032), .I2 (g1027));
ND2X1 gate9977(.O (I17288), .I1 (g11366), .I2 (g11363));
ND2X1 gate9978(.O (I13859), .I1 (g1448), .I2 (I13857));
ND2X1 gate9979(.O (g7548), .I1 (I11981), .I2 (I11982));
ND2X1 gate9980(.O (I13858), .I1 (g8538), .I2 (I13857));
ND2X1 gate9981(.O (I11996), .I1 (g7107), .I2 (I11995));
ND3X1 gate9982(.O (g8743), .I1 (g8617), .I2 (g6971), .I3 (g6964));
ND2X1 gate9983(.O (I5880), .I1 (g2115), .I2 (I5878));
ND2X1 gate9984(.O (g10513), .I1 (g10441), .I2 (g5345));
ND2X1 gate9985(.O (g8411), .I1 (I13538), .I2 (I13539));
ND2X1 gate9986(.O (I8626), .I1 (g511), .I2 (I8624));
ND2X1 gate9987(.O (g10505), .I1 (g10432), .I2 (g5938));
ND2X1 gate9988(.O (I5612), .I1 (g1280), .I2 (I5611));
ND2X1 gate9989(.O (g4821), .I1 (I8179), .I2 (I8180));
ND2X1 gate9990(.O (I12076), .I1 (g174), .I2 (I12074));
ND2X1 gate9991(.O (I12085), .I1 (g6980), .I2 (g1470));
ND2X1 gate9992(.O (g7567), .I1 (I12020), .I2 (I12021));
ND2X1 gate9993(.O (I5128), .I1 (g1389), .I2 (I5126));
ND2X1 gate9994(.O (I6489), .I1 (g1227), .I2 (I6487));
ND2X1 gate9995(.O (g7593), .I1 (I12114), .I2 (I12115));
ND2X1 gate9996(.O (I8778), .I1 (g4630), .I2 (g1137));
ND2X1 gate9997(.O (g10149), .I1 (I15442), .I2 (I15443));
ND2X1 gate9998(.O (I13902), .I1 (g1428), .I2 (I13900));
ND2X1 gate9999(.O (I13301), .I1 (g1936), .I2 (I13300));
ND2X1 gate10000(.O (g3215), .I1 (g2564), .I2 (g1822));
ND4X1 gate10001(.O (g7996), .I1 (g7011), .I2 (g7574), .I3 (g7562), .I4 (g6974));
ND2X1 gate10002(.O (I4985), .I1 (g999), .I2 (g1003));
ND2X1 gate10003(.O (I14444), .I1 (g1834), .I2 (I14442));
ND4X1 gate10004(.O (g8000), .I1 (g7011), .I2 (g7574), .I3 (g7562), .I4 (g7550));
ND2X1 gate10005(.O (I5166), .I1 (g1499), .I2 (I5164));
ND2X1 gate10006(.O (I17460), .I1 (g11449), .I2 (I17459));
ND2X1 gate10007(.O (g3008), .I1 (g2444), .I2 (g878));
ND2X1 gate10008(.O (I6836), .I1 (g3287), .I2 (g806));
ND2X1 gate10009(.O (I5529), .I1 (g1265), .I2 (I5528));
ND2X1 gate10010(.O (g10229), .I1 (I15608), .I2 (I15609));
ND2X1 gate10011(.O (I13661), .I1 (g8322), .I2 (I13659));
ND2X1 gate10012(.O (I13895), .I1 (g1436), .I2 (I13893));
ND2X1 gate10013(.O (g2303), .I1 (I5342), .I2 (I5343));
ND2X1 gate10014(.O (I12039), .I1 (g6990), .I2 (I12038));
ND2X1 gate10015(.O (g5592), .I1 (I9007), .I2 (I9008));
ND2X1 gate10016(.O (I12038), .I1 (g6990), .I2 (g1466));
ND2X1 gate10017(.O (g3322), .I1 (I6488), .I2 (I6489));
ND2X1 gate10018(.O (I8561), .I1 (g4227), .I2 (g491));
ND2X1 gate10019(.O (I8527), .I1 (g4879), .I2 (g481));
ND2X1 gate10020(.O (I12143), .I1 (g7089), .I2 (g158));
ND2X1 gate10021(.O (I5619), .I1 (g1766), .I2 (I5618));
ND2X1 gate10022(.O (g10386), .I1 (I15879), .I2 (I15880));
ND2X1 gate10023(.O (I11980), .I1 (g6957), .I2 (g1482));
ND2X1 gate10024(.O (I6837), .I1 (g3287), .I2 (I6836));
ND2X1 gate10025(.O (I4973), .I1 (g995), .I2 (I4971));
ND2X1 gate10026(.O (I13888), .I1 (g1440), .I2 (I13886));
ND2X1 gate10027(.O (g7558), .I1 (I12003), .I2 (I12004));
ND2X1 gate10028(.O (I17494), .I1 (g3623), .I2 (I17492));
ND2X1 gate10029(.O (g11491), .I1 (I17493), .I2 (I17494));
ND2X1 gate10030(.O (I16045), .I1 (g833), .I2 (I16044));
ND2X1 gate10031(.O (I7684), .I1 (g1023), .I2 (I7683));
ND2X1 gate10032(.O (g4130), .I1 (g3044), .I2 (g2518));
ND2X1 gate10033(.O (I8771), .I1 (g4619), .I2 (I8770));
ND2X1 gate10034(.O (I13546), .I1 (g8259), .I2 (I13544));
ND2X1 gate10035(.O (I13089), .I1 (g8006), .I2 (g1840));
ND2X1 gate10036(.O (g2117), .I1 (I5024), .I2 (I5025));
ND2X1 gate10037(.O (g5119), .I1 (I8514), .I2 (I8515));
ND2X1 gate10038(.O (g5319), .I1 (I8804), .I2 (I8805));
ND2X1 gate10039(.O (I15899), .I1 (g857), .I2 (I15898));
ND2X1 gate10040(.O (I5606), .I1 (g1153), .I2 (I5604));
ND2X1 gate10041(.O (I15898), .I1 (g857), .I2 (g10287));
ND2X1 gate10042(.O (I16032), .I1 (g10368), .I2 (I16030));
ND2X1 gate10043(.O (I17401), .I1 (g11418), .I2 (I17400));
ND2X1 gate10044(.O (I13659), .I1 (g1945), .I2 (g8322));
ND2X1 gate10045(.O (I8738), .I1 (g4607), .I2 (g1121));
ND2X1 gate10046(.O (I13250), .I1 (g8148), .I2 (I13248));
ND2X1 gate10047(.O (I15718), .I1 (g10229), .I2 (I15716));
ND2X1 gate10048(.O (I9008), .I1 (g1791), .I2 (I9006));
ND2X1 gate10049(.O (I6176), .I1 (g2177), .I2 (g197));
ND2X1 gate10050(.O (I7865), .I1 (g774), .I2 (I7863));
ND2X1 gate10051(.O (g5274), .I1 (I8729), .I2 (I8730));
ND2X1 gate10052(.O (I5341), .I1 (g315), .I2 (g426));
ND2X1 gate10053(.O (I17305), .I1 (g11381), .I2 (g11377));
ND2X1 gate10054(.O (I17053), .I1 (g11249), .I2 (I17051));
ND2X1 gate10055(.O (g5125), .I1 (I8528), .I2 (I8529));
ND2X1 gate10056(.O (I12216), .I1 (g2518), .I2 (I12214));
ND2X1 gate10057(.O (I6225), .I1 (g2544), .I2 (I6224));
ND2X1 gate10058(.O (I5879), .I1 (g2120), .I2 (I5878));
ND2X1 gate10059(.O (g3221), .I1 (g1834), .I2 (g2564));
ND2X1 gate10060(.O (I14270), .I1 (g8840), .I2 (g1822));
ND2X1 gate10061(.O (I6124), .I1 (g2215), .I2 (g1419));
ND2X1 gate10062(.O (I6324), .I1 (g1864), .I2 (I6322));
ND2X1 gate10063(.O (I13867), .I1 (g8523), .I2 (g1403));
ND2X1 gate10064(.O (I13894), .I1 (g8529), .I2 (I13893));
ND2X1 gate10065(.O (I6469), .I1 (g2479), .I2 (I6467));
ND2X1 gate10066(.O (I8663), .I1 (g4286), .I2 (I8662));
ND2X1 gate10067(.O (g7523), .I1 (I11908), .I2 (I11909));
ND2X1 gate10068(.O (I6177), .I1 (g2177), .I2 (I6176));
ND2X1 gate10069(.O (g5187), .I1 (I8590), .I2 (I8591));
ND2X1 gate10070(.O (I6287), .I1 (g2091), .I2 (g981));
ND2X1 gate10071(.O (I8762), .I1 (g4616), .I2 (I8761));
ND2X1 gate10072(.O (I15871), .I1 (g10358), .I2 (I15870));
ND3X1 gate10073(.O (g8840), .I1 (g8542), .I2 (g8541), .I3 (g8760));
ND2X1 gate10074(.O (g2250), .I1 (I5264), .I2 (I5265));
ND2X1 gate10075(.O (I8590), .I1 (g4251), .I2 (I8589));
ND2X1 gate10076(.O (I6199), .I1 (g2525), .I2 (g766));
ND2X1 gate10077(.O (I14218), .I1 (g605), .I2 (I14216));
ND2X1 gate10078(.O (g8190), .I1 (g6027), .I2 (g7978));
ND2X1 gate10079(.O (I5284), .I1 (g762), .I2 (I5282));
ND2X1 gate10080(.O (I17485), .I1 (g11384), .I2 (g11474));
ND2X1 gate10081(.O (I4965), .I1 (g406), .I2 (I4964));
ND2X1 gate10082(.O (I5591), .I1 (g1696), .I2 (g1703));
ND2X1 gate10083(.O (g8501), .I1 (g3760), .I2 (g8366));
ND2X1 gate10084(.O (I15451), .I1 (g10058), .I2 (g10051));
ND2X1 gate10085(.O (g8942), .I1 (g8823), .I2 (g4921));
ND2X1 gate10086(.O (I13877), .I1 (g8535), .I2 (I13876));
ND2X1 gate10087(.O (g7269), .I1 (I11509), .I2 (I11510));
ND2X1 gate10088(.O (I4996), .I1 (g416), .I2 (I4995));
ND2X1 gate10089(.O (I6144), .I1 (g1976), .I2 (I6143));
ND2X1 gate10090(.O (I17567), .I1 (g11496), .I2 (g1610));
ND2X1 gate10091(.O (g7572), .I1 (I12039), .I2 (I12040));
ND2X1 gate10092(.O (I6207), .I1 (g2534), .I2 (g802));
ND2X1 gate10093(.O (I14277), .I1 (g8847), .I2 (g1828));
ND2X1 gate10094(.O (I16059), .I1 (g841), .I2 (I16058));
ND2X1 gate10095(.O (I16025), .I1 (g2701), .I2 (I16023));
ND2X1 gate10096(.O (I8563), .I1 (g491), .I2 (I8561));
ND2X1 gate10097(.O (g3524), .I1 (g3209), .I2 (g3221));
ND2X1 gate10098(.O (I16058), .I1 (g841), .I2 (g10372));
ND2X1 gate10099(.O (I5204), .I1 (g374), .I2 (I5202));
ND2X1 gate10100(.O (I6488), .I1 (g2306), .I2 (I6487));
ND4X1 gate10101(.O (g3818), .I1 (g3056), .I2 (g3071), .I3 (g2310), .I4 (g3003));
ND2X1 gate10102(.O (I16044), .I1 (g833), .I2 (g10370));
ND2X1 gate10103(.O (g3717), .I1 (I6880), .I2 (I6881));
ND2X1 gate10104(.O (I13077), .I1 (g1872), .I2 (I13076));
ND2X1 gate10105(.O (g10043), .I1 (I15257), .I2 (I15258));
ND2X1 gate10106(.O (I11280), .I1 (g6485), .I2 (I11278));
ND2X1 gate10107(.O (I6825), .I1 (g3281), .I2 (g770));
ND2X1 gate10108(.O (I4997), .I1 (g309), .I2 (I4995));
ND2X1 gate10109(.O (I13300), .I1 (g1936), .I2 (g8162));
ND2X1 gate10110(.O (I5323), .I1 (g1336), .I2 (g1341));
ND2X1 gate10111(.O (I6136), .I1 (g2496), .I2 (g378));
ND2X1 gate10112(.O (g5935), .I1 (I9558), .I2 (I9559));
ND2X1 gate10113(.O (I5528), .I1 (g1265), .I2 (g1015));
ND2X1 gate10114(.O (I6806), .I1 (g3268), .I2 (I6805));
ND2X1 gate10115(.O (I5530), .I1 (g1015), .I2 (I5528));
ND2X1 gate10116(.O (g10886), .I1 (g10807), .I2 (g10805));
ND2X1 gate10117(.O (g3106), .I1 (I6323), .I2 (I6324));
ND2X1 gate10118(.O (I13876), .I1 (g8535), .I2 (g1444));
ND2X1 gate10119(.O (I6322), .I1 (g2050), .I2 (g1864));
ND2X1 gate10120(.O (g3061), .I1 (g611), .I2 (g2374));
ND2X1 gate10121(.O (g2439), .I1 (g1814), .I2 (g1828));
ND4X1 gate10122(.O (g7947), .I1 (g7395), .I2 (g7390), .I3 (g7279), .I4 (g7369));
ND2X1 gate10123(.O (I9576), .I1 (g818), .I2 (I9574));
ND2X1 gate10124(.O (I13660), .I1 (g1945), .I2 (I13659));
ND2X1 gate10125(.O (g3200), .I1 (g1822), .I2 (g2061));
ND2X1 gate10126(.O (g4374), .I1 (I7684), .I2 (I7685));
ND2X1 gate10127(.O (I11916), .I1 (g1494), .I2 (I11914));
ND2X1 gate10128(.O (I5372), .I1 (g971), .I2 (I5371));
ND2X1 gate10129(.O (g3003), .I1 (g599), .I2 (g2399));
ND2X1 gate10130(.O (g8627), .I1 (I13887), .I2 (I13888));
ND2X1 gate10131(.O (I5618), .I1 (g1766), .I2 (g1771));
ND2X1 gate10132(.O (I6137), .I1 (g2496), .I2 (I6136));
ND2X1 gate10133(.O (I5343), .I1 (g426), .I2 (I5341));
ND2X1 gate10134(.O (I5282), .I1 (g758), .I2 (g762));
ND2X1 gate10135(.O (I13307), .I1 (g8190), .I2 (g617));
ND2X1 gate10136(.O (I13076), .I1 (g1872), .I2 (g7963));
ND2X1 gate10137(.O (I6807), .I1 (g471), .I2 (I6805));
ND2X1 gate10138(.O (I11243), .I1 (g790), .I2 (I11241));
ND2X1 gate10139(.O (I17585), .I1 (g11354), .I2 (I17584));
ND2X1 gate10140(.O (I12137), .I1 (g7110), .I2 (I12136));
ND2X1 gate10141(.O (I7564), .I1 (g654), .I2 (I7562));
ND2X1 gate10142(.O (g2970), .I1 (I6200), .I2 (I6201));
ND2X1 gate10143(.O (g10144), .I1 (I15431), .I2 (I15432));
ND2X1 gate10144(.O (I8788), .I1 (g1141), .I2 (I8786));
ND2X1 gate10145(.O (g7054), .I1 (I11242), .I2 (I11243));
ND2X1 gate10146(.O (I17052), .I1 (g10923), .I2 (I17051));
ND2X1 gate10147(.O (g2120), .I1 (I5035), .I2 (I5036));
ND2X1 gate10148(.O (g8616), .I1 (I13868), .I2 (I13869));
ND2X1 gate10149(.O (I5202), .I1 (g369), .I2 (g374));
ND2X1 gate10150(.O (I16088), .I1 (g10375), .I2 (I16086));
ND2X1 gate10151(.O (I16024), .I1 (g10426), .I2 (I16023));
ND2X1 gate10152(.O (g11490), .I1 (I17486), .I2 (I17487));
ND2X1 gate10153(.O (I5518), .I1 (g1019), .I2 (I5516));
ND3X1 gate10154(.O (g5118), .I1 (g2439), .I2 (g4806), .I3 (g4073));
ND2X1 gate10155(.O (I12021), .I1 (g166), .I2 (I12019));
NR2X1 gate10156(.O (g6392), .I1 (g5859), .I2 (g5938));
NR2X1 gate10157(.O (g5938), .I1 (g2764), .I2 (g4988));
NR2X1 gate10158(.O (g2478), .I1 (g1610), .I2 (g1737));
NR2X1 gate10159(.O (g10374), .I1 (g10347), .I2 (g3463));
NR4X1 gate10160(.O (g4278), .I1 (g3800), .I2 (g2593), .I3 (g2586), .I4 (g3776));
NR2X1 gate10161(.O (g10424), .I1 (g10292), .I2 (g4620));
NR2X1 gate10162(.O (g10383), .I1 (g10318), .I2 (g2998));
NR2X1 gate10163(.O (g3118), .I1 (g2521), .I2 (g2514));
NR2X1 gate10164(.O (g9815), .I1 (g9392), .I2 (g9367));
NR2X1 gate10165(.O (g11077), .I1 (g10970), .I2 (g10971));
NR3X1 gate10166(.O (g9746), .I1 (g9454), .I2 (g9274), .I3 (g9292));
NR3X1 gate10167(.O (g3879), .I1 (g3141), .I2 (g2354), .I3 (g2353));
NR2X1 gate10168(.O (g10285), .I1 (g10276), .I2 (g3566));
NR2X1 gate10169(.O (g11480), .I1 (g11456), .I2 (g4567));
NR2X1 gate10170(.O (g4076), .I1 (g1707), .I2 (g2864));
NR2X1 gate10171(.O (g10570), .I1 (g10542), .I2 (g10324));
NR2X1 gate10172(.O (g10239), .I1 (g9317), .I2 (g10179));
NR2X1 gate10173(.O (g10594), .I1 (g10480), .I2 (g10521));
NR2X1 gate10174(.O (g9426), .I1 (g9052), .I2 (g9030));
NR2X1 gate10175(.O (g10382), .I1 (g10314), .I2 (g2998));
NR4X1 gate10176(.O (g4672), .I1 (g3501), .I2 (g2669), .I3 (g2662), .I4 (g3479));
NR2X1 gate10177(.O (g5360), .I1 (g2071), .I2 (g4225));
NR4X1 gate10178(.O (g9387), .I1 (g9010), .I2 (g9240), .I3 (g9223), .I4 (I14596));
NR2X1 gate10179(.O (g10438), .I1 (g10356), .I2 (g3566));
NR4X1 gate10180(.O (g4613), .I1 (g3077), .I2 (g3491), .I3 (g2662), .I4 (g2655));
NR4X1 gate10181(.O (g9391), .I1 (g9010), .I2 (g9240), .I3 (g9223), .I4 (I14602));
NR3X1 gate10182(.O (g4572), .I1 (g3419), .I2 (g3408), .I3 (g3628));
NR3X1 gate10183(.O (g9757), .I1 (g9454), .I2 (g9274), .I3 (g9292));
NR2X1 gate10184(.O (g9416), .I1 (g9052), .I2 (g9030));
NR4X1 gate10185(.O (g9874), .I1 (g9519), .I2 (g9536), .I3 (g9579), .I4 (I15033));
NR2X1 gate10186(.O (g9654), .I1 (g9125), .I2 (g9173));
NR4X1 gate10187(.O (g9880), .I1 (g9751), .I2 (g9536), .I3 (g9557), .I4 (I15051));
NR4X1 gate10188(.O (g4873), .I1 (g3292), .I2 (g2593), .I3 (g2586), .I4 (g3776));
NR2X1 gate10189(.O (g2807), .I1 (g22), .I2 (g2320));
NR2X1 gate10190(.O (g10441), .I1 (g10351), .I2 (g3566));
NR4X1 gate10191(.O (g4639), .I1 (g3501), .I2 (g2669), .I3 (g2662), .I4 (g2655));
NR2X1 gate10192(.O (g10435), .I1 (g10332), .I2 (g3507));
NR2X1 gate10193(.O (g10849), .I1 (g10739), .I2 (g3903));
NR4X1 gate10194(.O (g9606), .I1 (g9125), .I2 (g9111), .I3 (g9173), .I4 (g9151));
NR4X1 gate10195(.O (g9879), .I1 (g9747), .I2 (g9536), .I3 (g9566), .I4 (I15048));
NR2X1 gate10196(.O (g9506), .I1 (g9052), .I2 (g9030));
NR2X1 gate10197(.O (g6155), .I1 (g4974), .I2 (g2864));
NR2X1 gate10198(.O (g6355), .I1 (g6032), .I2 (g6023));
NR2X1 gate10199(.O (g9615), .I1 (g9052), .I2 (g9030));
NR2X1 gate10200(.O (g10371), .I1 (g10344), .I2 (g3463));
NR2X1 gate10201(.O (g9591), .I1 (g9125), .I2 (g9151));
NR2X1 gate10202(.O (g10359), .I1 (g10227), .I2 (g4620));
NR2X1 gate10203(.O (g10434), .I1 (g10352), .I2 (g3566));
NR2X1 gate10204(.O (g10358), .I1 (g10226), .I2 (g4620));
NR3X1 gate10205(.O (g9750), .I1 (g9454), .I2 (g9274), .I3 (g9292));
NR2X1 gate10206(.O (g10291), .I1 (g10247), .I2 (g3113));
NR4X1 gate10207(.O (g4227), .I1 (g3292), .I2 (g3793), .I3 (g2586), .I4 (g2579));
NR4X1 gate10208(.O (g9655), .I1 (g9010), .I2 (g9240), .I3 (g9223), .I4 (I14776));
NR4X1 gate10209(.O (g9410), .I1 (g9010), .I2 (g9240), .I3 (g9223), .I4 (I14607));
NR4X1 gate10210(.O (g9667), .I1 (g9125), .I2 (g9111), .I3 (g9173), .I4 (g9151));
NR2X1 gate10211(.O (g10563), .I1 (g10539), .I2 (g10322));
NR2X1 gate10212(.O (g9776), .I1 (g9392), .I2 (g9367));
NR2X1 gate10213(.O (g10324), .I1 (g9317), .I2 (g10244));
NR3X1 gate10214(.O (g4455), .I1 (g3543), .I2 (g3419), .I3 (g3408));
NR4X1 gate10215(.O (g9878), .I1 (g9754), .I2 (g9536), .I3 (g9560), .I4 (I15045));
NR2X1 gate10216(.O (g10360), .I1 (g10277), .I2 (g3566));
NR4X1 gate10217(.O (g9882), .I1 (g9742), .I2 (g9536), .I3 (g9563), .I4 (I15057));
NR2X1 gate10218(.O (g10370), .I1 (g10343), .I2 (g3463));
NR4X1 gate10219(.O (g4605), .I1 (g3077), .I2 (g2669), .I3 (g3485), .I4 (g2655));
NR2X1 gate10220(.O (g10420), .I1 (g10329), .I2 (g3744));
NR2X1 gate10221(.O (g10562), .I1 (g10483), .I2 (g10529));
NR2X1 gate10222(.O (g10427), .I1 (g10296), .I2 (g4620));
NR2X1 gate10223(.O (g5780), .I1 (g2112), .I2 (g4921));
NR2X1 gate10224(.O (g10385), .I1 (g10321), .I2 (g2998));
NR2X1 gate10225(.O (g10376), .I1 (g10323), .I2 (g3113));
NR2X1 gate10226(.O (g10426), .I1 (g10294), .I2 (g4620));
NR4X1 gate10227(.O (g4601), .I1 (g3077), .I2 (g2669), .I3 (g2662), .I4 (g3479));
NR2X1 gate10228(.O (g5573), .I1 (g4117), .I2 (g4432));
NR2X1 gate10229(.O (g9808), .I1 (g9392), .I2 (g9367));
NR2X1 gate10230(.O (g5999), .I1 (g2753), .I2 (g4953));
NR3X1 gate10231(.O (g9759), .I1 (g9454), .I2 (g9274), .I3 (g9292));
NR2X1 gate10232(.O (g6037), .I1 (g3305), .I2 (g5614));
NR2X1 gate10233(.O (g10287), .I1 (g10275), .I2 (g3463));
NR2X1 gate10234(.O (g5034), .I1 (g3524), .I2 (g4593));
NR4X1 gate10235(.O (g9362), .I1 (g9010), .I2 (g9240), .I3 (g9223), .I4 (I14585));
NR4X1 gate10236(.O (g9881), .I1 (g9516), .I2 (g9536), .I3 (g9573), .I4 (I15054));
NR2X1 gate10237(.O (g10443), .I1 (g10353), .I2 (g3566));
NR2X1 gate10238(.O (g10286), .I1 (g10271), .I2 (g3463));
NR3X1 gate10239(.O (g4276), .I1 (g4065), .I2 (g3261), .I3 (g2500));
NR4X1 gate10240(.O (g4616), .I1 (g3077), .I2 (g3491), .I3 (g2662), .I4 (g3479));
NR2X1 gate10241(.O (g10363), .I1 (g10355), .I2 (g3566));
NR2X1 gate10242(.O (g2862), .I1 (g2315), .I2 (g2305));
NR2X1 gate10243(.O (g10373), .I1 (g10346), .I2 (g3463));
NR2X1 gate10244(.O (g10423), .I1 (g10290), .I2 (g4620));
NR3X1 gate10245(.O (g9758), .I1 (g9454), .I2 (g9274), .I3 (g9292));
NR3X1 gate10246(.O (g9589), .I1 (g9125), .I2 (g9173), .I3 (g9151));
NR2X1 gate10247(.O (g9803), .I1 (g9392), .I2 (g9367));
NR2X1 gate10248(.O (g10430), .I1 (g10349), .I2 (g3566));
NR2X1 gate10249(.O (g9421), .I1 (g9052), .I2 (g9030));
NR2X1 gate10250(.O (g10362), .I1 (g10228), .I2 (g3507));
NR2X1 gate10251(.O (g2791), .I1 (g2187), .I2 (g750));
NR2X1 gate10252(.O (g9817), .I1 (g9392), .I2 (g9367));
NR4X1 gate10253(.O (g9605), .I1 (g9125), .I2 (g9111), .I3 (g9173), .I4 (g9151));
NR2X1 gate10254(.O (g10372), .I1 (g10345), .I2 (g3463));
NR2X1 gate10255(.O (g9669), .I1 (g9392), .I2 (g9367));
NR2X1 gate10256(.O (g10422), .I1 (g10289), .I2 (g4620));
NR2X1 gate10257(.O (g10436), .I1 (g10354), .I2 (g3566));
NR4X1 gate10258(.O (g5556), .I1 (g4787), .I2 (g2695), .I3 (g2299), .I4 (g2031));
NR4X1 gate10259(.O (g4286), .I1 (g3800), .I2 (g2593), .I3 (g3784), .I4 (g2579));
NR2X1 gate10260(.O (g4974), .I1 (g4502), .I2 (g3714));
NR2X1 gate10261(.O (g9779), .I1 (g9392), .I2 (g9367));
NR2X1 gate10262(.O (g9423), .I1 (g9052), .I2 (g9030));
NR2X1 gate10263(.O (g5350), .I1 (g4163), .I2 (g4872));
NR4X1 gate10264(.O (g9361), .I1 (g9010), .I2 (g9240), .I3 (g9223), .I4 (I14582));
NR4X1 gate10265(.O (g2459), .I1 (g1645), .I2 (g1642), .I3 (g1651), .I4 (g1648));
NR2X1 gate10266(.O (g10381), .I1 (g10310), .I2 (g2998));
NR4X1 gate10267(.O (g4259), .I1 (g3292), .I2 (g3793), .I3 (g3784), .I4 (g3776));
NR2X1 gate10268(.O (g10522), .I1 (g10486), .I2 (g10239));
NR2X1 gate10269(.O (g5392), .I1 (g3369), .I2 (g4258));
NR3X1 gate10270(.O (g4122), .I1 (g3291), .I2 (g2410), .I3 (g2538));
NR2X1 gate10271(.O (g6023), .I1 (g2763), .I2 (g4975));
NR2X1 gate10272(.O (g3462), .I1 (g2187), .I2 (g2795));
NR4X1 gate10273(.O (g4218), .I1 (g3292), .I2 (g2593), .I3 (g3784), .I4 (g3776));
NR4X1 gate10274(.O (g4267), .I1 (g3800), .I2 (g2593), .I3 (g2586), .I4 (g2579));
NR4X1 gate10275(.O (g4677), .I1 (g3501), .I2 (g2669), .I3 (g3485), .I4 (g2655));
NR2X1 gate10276(.O (g9646), .I1 (g9125), .I2 (g9151));
NR2X1 gate10277(.O (g2863), .I1 (g2316), .I2 (g2309));
NR4X1 gate10278(.O (g9616), .I1 (g9010), .I2 (g9240), .I3 (g9223), .I4 (I14751));
NR2X1 gate10279(.O (g6032), .I1 (g3430), .I2 (g5039));
NR4X1 gate10280(.O (g9647), .I1 (g9125), .I2 (g9111), .I3 (g9173), .I4 (g9151));
NR2X1 gate10281(.O (g5859), .I1 (g3362), .I2 (g4943));
NR2X1 gate10282(.O (g10433), .I1 (g10330), .I2 (g3507));
NR2X1 gate10283(.O (g10368), .I1 (g10342), .I2 (g3463));
NR4X1 gate10284(.O (g4251), .I1 (g3292), .I2 (g3793), .I3 (g3784), .I4 (g2579));
NR4X1 gate10285(.O (g9876), .I1 (g9522), .I2 (g9536), .I3 (g9576), .I4 (I15039));
NR4X1 gate10286(.O (g9656), .I1 (g9010), .I2 (g9240), .I3 (g9223), .I4 (I14779));
NR2X1 gate10287(.O (g8303), .I1 (g8209), .I2 (g4811));
NR2X1 gate10288(.O (g10429), .I1 (g10326), .I2 (g3507));
NR2X1 gate10289(.O (g10428), .I1 (g10335), .I2 (g4620));
NR4X1 gate10290(.O (g4234), .I1 (g3292), .I2 (g3793), .I3 (g2586), .I4 (g3776));
NR4X1 gate10291(.O (g9877), .I1 (g9512), .I2 (g9536), .I3 (g9569), .I4 (I15042));
NR2X1 gate10292(.O (g5186), .I1 (g2047), .I2 (g4401));
NR2X1 gate10293(.O (g9489), .I1 (g9052), .I2 (g9030));
NR4X1 gate10294(.O (g4619), .I1 (g3077), .I2 (g3491), .I3 (g3485), .I4 (g2655));
NR2X1 gate10295(.O (g10432), .I1 (g10350), .I2 (g3566));
NR2X1 gate10296(.O (g5345), .I1 (g2754), .I2 (g4835));
NR2X1 gate10297(.O (g5763), .I1 (g5350), .I2 (g5345));
NR2X1 gate10298(.O (g10375), .I1 (g10288), .I2 (g3463));
NR4X1 gate10299(.O (g4879), .I1 (g3292), .I2 (g2593), .I3 (g3784), .I4 (g2579));
NR4X1 gate10300(.O (g4607), .I1 (g3077), .I2 (g2669), .I3 (g3485), .I4 (g3479));
NR2X1 gate10301(.O (g10425), .I1 (g10293), .I2 (g4620));
NR2X1 gate10302(.O (g3107), .I1 (g2501), .I2 (g2499));
NR2X1 gate10303(.O (g10322), .I1 (g9317), .I2 (g10272));
NR4X1 gate10304(.O (g4630), .I1 (g3077), .I2 (g3491), .I3 (g3485), .I4 (g3479));
NR2X1 gate10305(.O (g10364), .I1 (g10327), .I2 (g3744));
NR2X1 gate10306(.O (g9781), .I1 (g9392), .I2 (g9367));
endmodule